netcdf sampling_error_correction_table.Lanai {
dimensions:
	bins = 200 ;
	ens_sizes = UNLIMITED ; // (40 currently)
variables:
	int count(ens_sizes, bins) ;
		count:description = "number of samples in each bin" ;
	double true_corr_mean(ens_sizes, bins) ;
	double alpha(ens_sizes, bins) ;
		alpha:description = "sampling error correction factors" ;
	int ens_sizes(ens_sizes) ;
		ens_sizes:description = "ensemble size used for calculation" ;

// global attributes:
		:num_samples = 100000000 ;
		:title = "Sampling Error Corrections for fixed ensemble sizes." ;
		:version = "original values as from final_full.nn" ;
		:reference = "Anderson, J., 2012: Localization and Sampling Error Correction in Ensemble Kalman Filter Data Assimilation. Mon. Wea. Rev., 140, 2359-2371, doi: 10.1175/MWR-D-11-00013.1." ;
data:

 count =
  1595111, 1335139, 1202476, 1108193, 1032044, 972567, 923878, 878705, 
    843621, 810724, 780965, 753744, 730593, 706765, 687843, 670227, 652400, 
    637266, 621868, 608162, 595985, 583360, 571664, 561321, 550800, 539950, 
    531544, 524795, 516024, 507443, 501295, 493355, 486254, 480777, 472541, 
    467497, 461633, 456455, 451490, 446090, 441356, 437126, 432731, 428825, 
    424707, 420738, 416533, 411667, 410361, 405248, 402402, 400308, 396944, 
    394242, 392538, 389079, 385135, 384303, 381512, 380006, 377310, 374221, 
    372652, 369642, 368548, 367687, 364874, 363338, 362465, 360560, 359552, 
    357804, 355872, 353660, 353987, 352615, 350843, 350571, 350051, 348216, 
    347249, 346969, 345261, 345698, 344547, 343728, 343819, 343168, 342391, 
    341424, 341107, 340567, 340182, 340382, 339327, 339172, 338873, 339027, 
    338815, 338822, 339042, 338994, 338783, 339155, 339272, 339456, 341262, 
    339713, 340491, 341506, 341276, 342084, 343221, 342982, 343520, 344331, 
    345638, 345837, 347060, 348506, 349012, 349367, 351800, 351309, 352008, 
    354390, 356307, 358118, 357725, 360592, 361144, 362988, 364284, 366403, 
    368082, 369802, 371474, 374354, 375266, 376959, 380985, 381576, 384335, 
    387385, 389636, 392904, 395954, 399230, 401882, 404021, 408702, 410771, 
    415803, 418922, 422247, 425668, 429091, 435115, 438581, 444647, 446836, 
    453191, 459023, 463366, 468984, 474953, 481818, 488505, 495273, 502777, 
    509544, 516885, 525532, 534718, 544033, 553238, 562186, 572772, 585218, 
    598488, 609839, 623066, 638879, 656184, 670997, 688257, 710282, 730055, 
    754217, 782803, 812167, 844026, 882253, 923157, 972622, 1032701, 1108366, 
    1204064, 1338799, 1595636,
  1165121, 1064500, 997879, 944350, 900836, 865493, 832286, 803534, 779990, 
    758056, 733530, 715958, 698534, 681550, 667325, 652075, 639336, 627456, 
    614658, 603693, 594263, 583977, 572658, 564161, 557758, 547219, 539834, 
    532181, 526005, 519656, 512460, 506545, 501376, 494959, 489079, 485058, 
    480510, 476022, 470391, 466511, 461680, 458067, 453792, 450377, 446209, 
    443508, 439127, 436269, 433596, 429587, 426403, 425054, 422239, 419529, 
    416862, 414537, 412049, 408874, 407719, 404078, 403280, 401721, 399644, 
    397300, 396555, 393032, 392472, 389586, 388504, 388229, 386802, 385568, 
    383476, 382144, 381397, 380141, 378233, 377286, 376895, 376005, 375385, 
    373951, 374300, 373324, 372640, 372544, 371138, 369894, 369496, 368415, 
    369605, 369359, 368383, 368110, 368755, 368327, 367629, 367946, 367724, 
    368101, 367087, 367633, 367830, 368615, 367665, 368478, 368610, 369234, 
    369573, 369162, 370129, 370572, 371575, 371683, 372038, 374328, 373733, 
    374521, 374956, 376490, 377550, 377953, 378276, 380302, 379745, 381311, 
    383073, 385766, 386019, 387502, 389999, 390463, 391939, 393176, 395527, 
    396070, 398998, 400807, 402487, 404789, 406252, 408836, 411736, 412771, 
    414741, 418263, 421274, 422696, 425026, 428748, 431149, 434267, 437538, 
    442017, 445543, 448432, 452969, 454613, 459336, 463494, 468118, 473456, 
    478105, 482830, 486219, 490531, 497315, 501963, 508311, 515976, 519582, 
    527289, 534407, 542993, 549254, 557704, 565914, 576366, 584722, 593546, 
    604590, 614920, 626150, 640277, 653971, 667935, 682893, 699060, 717399, 
    735795, 756646, 781235, 804251, 834564, 868346, 903953, 945960, 1000868, 
    1065825, 1165760,
  967014, 917065, 877665, 845191, 818791, 791981, 770308, 750047, 730591, 
    714452, 697711, 683259, 670193, 657172, 644870, 633929, 624438, 612575, 
    604082, 593554, 586349, 578345, 570571, 561967, 555349, 548805, 541878, 
    534849, 529584, 524044, 520667, 514080, 507523, 502924, 498134, 493901, 
    489516, 486087, 481142, 477754, 473111, 470511, 467128, 463552, 460300, 
    456981, 453319, 451048, 447826, 445301, 442176, 440112, 437585, 435611, 
    432751, 431081, 427119, 427021, 423956, 422644, 420404, 418062, 416897, 
    415137, 414495, 410986, 409776, 408886, 408644, 406188, 404230, 404256, 
    402293, 401315, 399988, 400124, 398079, 397038, 395721, 395850, 394145, 
    395028, 393735, 392730, 392009, 391991, 390244, 390231, 389574, 389007, 
    389310, 388651, 388645, 388016, 388310, 388187, 387888, 387521, 387682, 
    387816, 387624, 387659, 387370, 387866, 388882, 387947, 388197, 389115, 
    388856, 389887, 390271, 390614, 391449, 391892, 392955, 392759, 393283, 
    393107, 394412, 395412, 396357, 397238, 398244, 398906, 401345, 401280, 
    401586, 403385, 405078, 405476, 407606, 408065, 409572, 411248, 412588, 
    414210, 416490, 417900, 419637, 420962, 422571, 424537, 428407, 429242, 
    430906, 434613, 435515, 439353, 440551, 444376, 445881, 449345, 452446, 
    454563, 457603, 462134, 464864, 467473, 472707, 475264, 479290, 481916, 
    487602, 490601, 495405, 499839, 503643, 509077, 514179, 521289, 527665, 
    531199, 537933, 543790, 549834, 556639, 563194, 572554, 578921, 588005, 
    594665, 605295, 614504, 624129, 636274, 647847, 658542, 671664, 684151, 
    699180, 714783, 732298, 752442, 772038, 794430, 817802, 846809, 880567, 
    917780, 966564,
  857367, 827066, 800879, 781709, 759474, 742200, 724617, 709940, 696597, 
    682666, 669966, 657279, 646751, 637793, 626552, 618283, 608931, 600999, 
    593109, 586733, 578534, 572279, 564430, 558415, 552659, 547977, 540727, 
    535564, 529451, 526423, 520370, 515862, 511504, 507615, 503761, 499770, 
    495232, 491747, 487928, 484507, 482236, 477305, 474920, 471715, 468342, 
    465855, 462356, 460920, 458762, 455392, 453482, 450558, 447679, 446218, 
    442850, 441701, 439608, 438489, 437141, 433285, 433702, 431716, 429593, 
    428204, 427311, 424217, 423284, 421778, 421222, 419330, 418236, 416863, 
    416816, 414143, 414646, 412986, 412675, 411567, 410986, 410183, 408381, 
    408181, 408435, 406517, 406112, 406365, 405328, 404148, 404948, 405721, 
    401761, 403298, 402111, 403206, 402557, 401706, 402845, 403529, 401976, 
    402105, 402887, 401614, 402728, 402671, 402960, 402506, 402860, 403374, 
    403844, 404185, 404168, 404896, 405694, 406903, 405867, 407101, 407803, 
    408959, 409774, 409157, 410446, 410233, 412783, 412228, 413347, 415123, 
    415769, 416626, 417624, 419480, 420373, 421293, 423059, 424451, 425222, 
    426932, 429343, 430250, 433311, 433317, 435472, 438264, 438871, 440443, 
    442452, 444545, 447443, 448895, 451852, 454235, 456772, 459089, 462264, 
    465124, 466220, 469606, 473218, 475806, 478785, 481952, 486444, 488552, 
    493216, 496742, 500729, 505310, 509313, 512903, 518279, 521817, 525809, 
    532600, 537551, 543312, 548769, 554499, 560110, 566247, 572248, 579499, 
    588290, 594781, 602518, 611657, 619551, 629159, 638253, 649592, 659631, 
    671198, 683293, 695974, 711025, 724906, 744197, 760295, 779765, 803944, 
    826691, 857693,
  789427, 767816, 749642, 735932, 718890, 705776, 692203, 680746, 669979, 
    657605, 647836, 638263, 628711, 621393, 612211, 605480, 598198, 591624, 
    586031, 577085, 572018, 567892, 559630, 553773, 550067, 545968, 539578, 
    535207, 531362, 526393, 520233, 515907, 513308, 510456, 505525, 502062, 
    498636, 497009, 493743, 488730, 486186, 481699, 480188, 477362, 474735, 
    471653, 469679, 467135, 465069, 462402, 460068, 457203, 455879, 454143, 
    451963, 450106, 448026, 446481, 445008, 443798, 441848, 440923, 437722, 
    435345, 436074, 436403, 433190, 431462, 429666, 430694, 429874, 428849, 
    427320, 424851, 423739, 422815, 422140, 422647, 421123, 420940, 418957, 
    418822, 418516, 418102, 416849, 417429, 416646, 415892, 415802, 416426, 
    415157, 414820, 414431, 414336, 414062, 414531, 411851, 413410, 413770, 
    413738, 413931, 413377, 414013, 413751, 413406, 413283, 414805, 414734, 
    414720, 413260, 414384, 416110, 416742, 418108, 417218, 417641, 418120, 
    418604, 419603, 420045, 421521, 422893, 421742, 423909, 424851, 425816, 
    426447, 426130, 429023, 429202, 430066, 431445, 432547, 432949, 436848, 
    435957, 437686, 440253, 441008, 442827, 444184, 446410, 448610, 449541, 
    450472, 453191, 456358, 458345, 459333, 461171, 462271, 466060, 468426, 
    471522, 473396, 477352, 478046, 480654, 483295, 487204, 489748, 491997, 
    498603, 500444, 503526, 506020, 513136, 514275, 519330, 523816, 526369, 
    530345, 536396, 541070, 545680, 550226, 556165, 561971, 565464, 573938, 
    578570, 586233, 592994, 600201, 606987, 613509, 622487, 630341, 638559, 
    648003, 660090, 668864, 679352, 693222, 705792, 718738, 734827, 749170, 
    767715, 788710,
  741603, 727507, 711825, 701965, 690974, 676531, 664683, 657416, 649189, 
    640837, 632684, 623280, 617164, 608208, 602324, 595617, 589128, 582149, 
    575855, 571673, 567430, 561628, 554128, 550383, 545267, 540449, 535266, 
    532972, 529037, 523452, 520109, 517933, 515710, 511366, 507881, 504540, 
    501370, 499690, 496120, 493272, 489074, 486736, 483160, 481673, 478723, 
    477202, 474058, 471360, 470343, 468094, 466121, 463604, 462940, 460705, 
    458896, 456856, 454991, 454152, 451069, 450068, 447214, 446528, 445166, 
    444530, 443328, 442445, 440656, 439661, 440241, 438284, 436093, 435363, 
    434395, 434859, 432387, 432068, 431206, 428948, 429314, 428594, 428530, 
    426523, 426649, 427514, 426406, 425197, 424839, 424595, 423854, 424070, 
    423918, 424467, 423380, 422900, 423373, 423251, 422955, 421950, 423032, 
    423504, 421300, 421044, 421885, 422566, 422040, 423922, 423019, 424610, 
    425209, 423466, 423933, 424335, 426017, 426497, 427073, 426146, 425580, 
    427439, 429117, 427707, 429486, 430767, 431071, 431430, 433342, 433747, 
    434312, 434118, 435859, 437237, 439065, 438893, 440683, 441400, 443187, 
    444176, 444367, 446865, 449528, 450910, 450670, 453311, 454517, 456401, 
    457621, 458704, 460050, 461949, 464740, 465537, 469964, 471389, 472382, 
    476669, 478935, 479797, 482624, 486395, 487142, 489294, 492598, 496099, 
    498385, 502554, 504580, 509513, 510745, 517036, 518964, 523174, 525262, 
    530806, 533238, 539135, 543226, 547784, 550414, 556820, 561637, 565451, 
    571725, 577605, 583369, 589480, 596511, 602200, 608152, 615931, 623997, 
    632261, 639224, 647672, 659298, 667715, 677147, 689017, 698954, 713322, 
    725681, 741251,
  682532, 672433, 662470, 656685, 647358, 640528, 631088, 626600, 617530, 
    612023, 604592, 601066, 594977, 591459, 583295, 579810, 574472, 569790, 
    565700, 559090, 555745, 553137, 549995, 545176, 540486, 537348, 531798, 
    530159, 526702, 524017, 521549, 518883, 515242, 510873, 508194, 503748, 
    502678, 499076, 497956, 496104, 492744, 490018, 490422, 486348, 486945, 
    481479, 480878, 480137, 478683, 475268, 473705, 472387, 470366, 468465, 
    464770, 464078, 464797, 461905, 461094, 460210, 457998, 458962, 456902, 
    454025, 453905, 452620, 451973, 450731, 449204, 447587, 448086, 448216, 
    446610, 447488, 446299, 444292, 443093, 444402, 442384, 442573, 440642, 
    440786, 440053, 439045, 438629, 437575, 437206, 437868, 439678, 437263, 
    438255, 436423, 435203, 436226, 436476, 435612, 436511, 435042, 435738, 
    434694, 435021, 435582, 436830, 436427, 435850, 437452, 436788, 436177, 
    437952, 437527, 435554, 436023, 438957, 439876, 438585, 439813, 438202, 
    440910, 438961, 440403, 442633, 442750, 441406, 443890, 443824, 445496, 
    444788, 448378, 448518, 448615, 448990, 449575, 451601, 452326, 452478, 
    455205, 455825, 457083, 458825, 460192, 461902, 461801, 464330, 465817, 
    467397, 467362, 470451, 471450, 472846, 473952, 475572, 477500, 480538, 
    481967, 481811, 485919, 488652, 490937, 492341, 494339, 496538, 500423, 
    501265, 503208, 505547, 509788, 514619, 514763, 517025, 521180, 524706, 
    525579, 530752, 532334, 535802, 539349, 543182, 545745, 552733, 556839, 
    560711, 565600, 571475, 574715, 579059, 583438, 588217, 592688, 599776, 
    607083, 613344, 619859, 625804, 632052, 639854, 647415, 654260, 662723, 
    672584, 682455,
  646519, 639574, 632616, 627078, 620831, 615044, 609412, 603480, 599396, 
    593981, 589074, 583958, 579848, 576234, 572433, 566914, 563609, 559763, 
    556289, 551076, 549963, 545851, 542087, 538756, 535387, 532294, 529479, 
    526365, 523369, 521640, 519248, 516568, 513188, 510842, 509865, 505954, 
    503920, 501795, 499584, 498490, 495673, 494258, 492500, 490355, 488432, 
    486177, 485334, 483196, 482013, 480216, 478818, 478600, 475893, 473288, 
    472887, 472138, 471123, 468646, 468163, 466962, 465069, 463812, 463372, 
    462983, 461551, 460457, 459066, 457690, 457833, 457113, 456899, 456299, 
    454608, 454569, 452861, 453655, 451773, 451613, 451628, 449255, 450316, 
    449222, 448539, 448075, 448234, 447251, 447601, 446756, 446619, 445877, 
    445946, 446413, 445022, 445440, 445609, 444691, 445288, 443968, 445815, 
    445402, 445078, 444369, 444806, 445899, 445364, 445888, 445842, 446011, 
    447417, 445193, 446909, 446790, 447150, 447549, 448492, 447892, 448822, 
    448459, 448588, 450291, 449983, 450863, 451693, 452993, 452832, 453536, 
    454763, 454486, 455308, 457235, 456826, 458918, 459145, 460122, 460174, 
    462171, 463088, 464267, 464579, 466214, 467274, 468007, 468842, 470290, 
    471772, 473585, 475531, 476485, 476939, 478942, 481367, 482796, 483754, 
    485700, 487513, 488305, 490757, 493020, 494158, 496473, 498647, 500693, 
    502484, 504698, 507376, 509853, 511980, 513872, 516456, 518464, 521786, 
    524830, 526602, 529937, 532462, 536061, 539388, 542154, 545192, 549096, 
    553042, 555458, 559156, 563810, 566977, 571693, 575609, 579406, 583494, 
    588849, 592599, 598995, 603185, 609178, 613932, 619316, 626626, 633207, 
    639391, 645894,
  633279, 626601, 621914, 617245, 610211, 605809, 602022, 594893, 588452, 
    584474, 581750, 580940, 574665, 569555, 566736, 563740, 561038, 555457, 
    553516, 549438, 546208, 542511, 539557, 535220, 532382, 530633, 526872, 
    523836, 522571, 519474, 518041, 516846, 515061, 510025, 506459, 508952, 
    506369, 503716, 500697, 498636, 497448, 496275, 492110, 492082, 489775, 
    489053, 485571, 484468, 482427, 483381, 480389, 480281, 476584, 475805, 
    474766, 472568, 472899, 472180, 470420, 468796, 469049, 468967, 466651, 
    464701, 463250, 462588, 462930, 462124, 462132, 458349, 458334, 458160, 
    457944, 457012, 456444, 456091, 455655, 453256, 452719, 453851, 453106, 
    452930, 452280, 452709, 452127, 452663, 449917, 449531, 451404, 450459, 
    448819, 449319, 448438, 450840, 448847, 449031, 450275, 449194, 449135, 
    448376, 450218, 448445, 447012, 448423, 450962, 448119, 448742, 449411, 
    450268, 450283, 450750, 449420, 450015, 451507, 453200, 453631, 452446, 
    450527, 451359, 452012, 454400, 454560, 455319, 455376, 455904, 457360, 
    457615, 458568, 458139, 459801, 461742, 461337, 463252, 463271, 463931, 
    464975, 464565, 467350, 466516, 469060, 468216, 472898, 473185, 473587, 
    472851, 474924, 476153, 477232, 478484, 481855, 482845, 482488, 485687, 
    487289, 488227, 491333, 490746, 494938, 496891, 496868, 498943, 501047, 
    502779, 506168, 508282, 509233, 509802, 511857, 516257, 518681, 520661, 
    523262, 524958, 527908, 532323, 535027, 538022, 540108, 542479, 544598, 
    549694, 551159, 555768, 557479, 561847, 565663, 569444, 573779, 578274, 
    581414, 584617, 592645, 594029, 600381, 604614, 610526, 615133, 622177, 
    626918, 632869,
  622097, 617087, 611697, 607939, 601621, 598028, 591913, 589281, 584555, 
    580569, 575840, 573433, 569579, 565083, 561726, 558638, 555436, 551359, 
    549074, 546146, 542198, 540256, 538386, 534492, 532225, 528989, 527488, 
    525411, 520989, 519428, 518118, 514136, 513588, 510344, 508514, 506681, 
    503939, 502296, 500691, 498441, 498012, 495177, 494269, 493813, 490134, 
    488867, 487694, 486627, 484681, 483262, 483004, 480326, 480452, 477714, 
    477591, 476133, 474098, 473841, 472356, 471927, 469815, 470196, 468468, 
    467790, 466558, 467510, 464531, 464154, 464041, 462945, 462573, 461975, 
    460711, 460670, 459371, 458470, 457839, 458955, 457323, 457206, 456083, 
    455935, 455356, 455157, 454745, 453830, 452765, 453214, 453057, 452925, 
    452753, 452686, 451721, 451282, 453599, 453313, 451998, 452454, 451591, 
    451120, 451630, 453096, 451585, 451876, 451248, 452843, 452285, 451735, 
    453321, 453953, 453584, 453456, 454834, 453050, 453981, 454796, 454839, 
    455082, 456610, 456691, 457528, 457205, 458111, 458185, 459417, 459667, 
    460531, 461546, 461321, 462659, 463688, 463864, 465686, 465314, 466194, 
    467259, 468722, 468504, 469366, 470848, 472321, 473231, 473924, 475408, 
    477028, 478121, 478968, 479397, 481483, 482129, 484449, 484742, 486983, 
    487703, 489920, 490763, 492584, 494992, 496504, 497433, 499084, 500936, 
    503577, 505213, 505635, 509662, 511546, 513233, 515551, 517482, 519276, 
    522009, 524192, 527418, 529266, 530682, 534456, 537456, 539261, 543927, 
    545392, 548927, 551457, 555331, 557399, 562899, 564634, 567549, 572419, 
    576791, 579230, 583694, 587645, 593156, 596809, 600911, 606998, 610884, 
    617458, 621987,
  605253, 599782, 597026, 592383, 588186, 584462, 581003, 579423, 575079, 
    570622, 565767, 564844, 559459, 556447, 555235, 551770, 550519, 546309, 
    544931, 540640, 539550, 536573, 531214, 529597, 528020, 526247, 523089, 
    522706, 520345, 518273, 516561, 513955, 512316, 511061, 507440, 507031, 
    504522, 501652, 500991, 500721, 498440, 496234, 495372, 493836, 492237, 
    490010, 489743, 489463, 488033, 487485, 483633, 483567, 483356, 480654, 
    481875, 482160, 478330, 475061, 475143, 476189, 474706, 472837, 471556, 
    471899, 471210, 470407, 468759, 468452, 466256, 465872, 466843, 467680, 
    465485, 464238, 464803, 465130, 464439, 463350, 461754, 461601, 461388, 
    460265, 461160, 460574, 460537, 458964, 457687, 458130, 457598, 457498, 
    459715, 458705, 456718, 457574, 458970, 459227, 457669, 457496, 456776, 
    457089, 455290, 458354, 456377, 458403, 456720, 457603, 457184, 457550, 
    458074, 460548, 459070, 459813, 458639, 458814, 458258, 458344, 459615, 
    460864, 460450, 460261, 463074, 463020, 461431, 462989, 463293, 464369, 
    465364, 466470, 465161, 466304, 467820, 468844, 468793, 469606, 471500, 
    471672, 473179, 474647, 474543, 475587, 474571, 475596, 476864, 478166, 
    479668, 482108, 481708, 482134, 483496, 484890, 486185, 487050, 488759, 
    489947, 489815, 492979, 495159, 495383, 495301, 497584, 499505, 502206, 
    503671, 505507, 506550, 508366, 509784, 511990, 514885, 516101, 517410, 
    519677, 520777, 525734, 525789, 529194, 530412, 534955, 535943, 537386, 
    539478, 542094, 545424, 548821, 552983, 554577, 556011, 560728, 562957, 
    566371, 570619, 573822, 578899, 579598, 581613, 586945, 593274, 596918, 
    599800, 605123,
  591647, 588567, 585647, 582557, 577359, 575513, 570482, 569182, 564382, 
    564253, 558409, 556310, 555330, 550821, 548644, 546960, 546531, 542523, 
    539955, 535928, 533800, 532112, 529289, 526513, 526226, 524401, 522292, 
    520500, 517028, 515456, 513070, 512784, 512750, 510341, 508006, 507874, 
    505403, 502602, 501266, 500131, 500440, 497776, 497055, 495148, 495820, 
    493111, 490716, 490238, 488718, 488638, 486835, 486715, 485535, 483229, 
    479300, 481340, 481268, 479782, 478296, 477730, 475235, 474471, 475764, 
    475072, 472799, 473410, 473787, 472353, 470812, 469710, 468434, 470604, 
    469981, 469005, 468690, 466278, 468084, 466590, 465052, 464691, 465819, 
    465229, 466024, 464251, 461650, 463589, 464259, 462565, 463030, 463068, 
    464510, 463162, 462047, 462072, 462261, 461499, 460524, 463686, 461820, 
    462523, 461479, 461483, 460520, 461328, 460680, 461466, 461373, 462616, 
    463910, 463459, 463054, 461865, 461839, 465333, 464163, 463194, 464569, 
    464467, 463804, 464150, 465644, 466751, 466243, 467470, 468605, 467454, 
    468339, 469587, 469600, 470426, 470039, 471219, 472487, 473552, 473229, 
    474428, 476343, 476520, 477370, 475765, 479064, 479324, 479344, 481016, 
    483217, 483408, 482959, 484950, 486805, 486810, 487976, 489189, 491757, 
    492360, 491747, 492445, 493145, 495316, 497962, 498745, 501722, 503276, 
    504218, 505800, 506982, 506446, 508254, 509589, 513509, 515270, 517691, 
    519056, 520525, 521209, 522840, 526006, 528963, 528419, 530437, 534077, 
    536259, 537901, 541549, 544810, 546642, 547794, 549764, 555077, 557275, 
    558900, 562255, 566509, 567564, 569280, 572298, 576647, 582813, 584712, 
    588145, 591210,
  581830, 579040, 575901, 573020, 570553, 566125, 564375, 562420, 558615, 
    557115, 553268, 551904, 547789, 546755, 544411, 541841, 539842, 537581, 
    535601, 533331, 530820, 530017, 527074, 525126, 523943, 522220, 521065, 
    518680, 516810, 516106, 513163, 512168, 510560, 510117, 508482, 505236, 
    504337, 502839, 502858, 500431, 499333, 497837, 497751, 495877, 494586, 
    493225, 493282, 491135, 490375, 488759, 487678, 486649, 485764, 484746, 
    484629, 483624, 482997, 482439, 481827, 481014, 478971, 478776, 477629, 
    477537, 474575, 476393, 475456, 474570, 474625, 472500, 473878, 473083, 
    471732, 472065, 470230, 470408, 470946, 469373, 468133, 467625, 469223, 
    468461, 468324, 467588, 466650, 467590, 467171, 467048, 465496, 466296, 
    466402, 465347, 465402, 465434, 465119, 464946, 464958, 465348, 465140, 
    464411, 466172, 465162, 466104, 465024, 465061, 465350, 465627, 466011, 
    466489, 465261, 467074, 467031, 466641, 466656, 466611, 468021, 467483, 
    467362, 467540, 469362, 468838, 469119, 469977, 470135, 470910, 471851, 
    471282, 471544, 473241, 473017, 473201, 474293, 474515, 475339, 477090, 
    476122, 478040, 478317, 479687, 479895, 481114, 482543, 481742, 482214, 
    483568, 484178, 486168, 485620, 487757, 488501, 488665, 490558, 490071, 
    492187, 494851, 494918, 495840, 497540, 497521, 499308, 500205, 502997, 
    503188, 505172, 506973, 506952, 508847, 509656, 512170, 513024, 515493, 
    516567, 517659, 520526, 521433, 523948, 525800, 527300, 528927, 531107, 
    532641, 534867, 536207, 539570, 541076, 543650, 546354, 547840, 551518, 
    552851, 555162, 558302, 560602, 564352, 567544, 568424, 572082, 575760, 
    578222, 581957,
  573682, 571452, 568787, 565586, 563847, 559727, 558118, 556672, 552400, 
    552140, 549606, 547845, 544325, 542221, 539420, 538877, 536274, 534573, 
    531322, 530214, 529873, 527745, 524889, 524430, 521179, 520951, 519086, 
    517646, 515528, 513701, 514293, 509401, 510140, 509025, 507341, 506322, 
    505672, 503194, 502265, 501189, 498734, 497240, 496656, 496375, 494563, 
    493635, 494042, 492117, 489977, 490271, 488746, 488629, 487242, 486926, 
    485975, 485280, 485066, 482840, 483128, 481514, 482743, 480442, 479173, 
    479954, 479661, 478236, 477716, 476425, 475119, 476720, 474744, 475220, 
    475034, 473040, 472940, 474390, 474162, 472783, 471945, 471611, 471575, 
    469865, 472369, 470155, 469827, 469897, 469558, 469140, 467597, 469113, 
    468538, 468405, 468237, 468780, 468311, 467670, 467996, 467662, 467817, 
    468410, 468748, 468358, 467065, 468871, 469101, 468739, 469121, 467650, 
    469464, 468035, 469911, 468633, 467917, 469313, 471511, 469755, 470904, 
    471885, 470831, 471728, 471660, 472445, 472797, 472279, 472445, 472991, 
    474090, 475457, 474795, 474989, 474292, 475787, 477331, 479299, 478921, 
    478717, 480213, 479728, 479968, 481630, 482190, 483459, 483006, 484634, 
    486053, 485516, 487114, 488783, 489263, 488717, 490456, 492868, 491339, 
    492237, 493290, 497006, 496391, 498030, 498852, 500426, 499832, 501306, 
    502710, 504264, 506410, 506271, 508714, 510066, 511401, 511488, 514079, 
    515125, 517267, 520064, 519006, 522192, 523068, 525356, 526466, 528031, 
    530361, 533068, 532720, 535965, 538342, 539949, 541898, 544051, 545241, 
    547665, 550347, 553174, 555728, 557657, 560023, 563410, 564280, 568993, 
    569937, 574176,
  561687, 560018, 557293, 554342, 553920, 550606, 549025, 547445, 544718, 
    544612, 540692, 539622, 537821, 535514, 534395, 533785, 530573, 530038, 
    528422, 526296, 524289, 523145, 521126, 521086, 520091, 517202, 515637, 
    514428, 513729, 512135, 511710, 509727, 508748, 507365, 506431, 504932, 
    504777, 503342, 502602, 501121, 499511, 499456, 496468, 497905, 497045, 
    495383, 494054, 494613, 493155, 491105, 491306, 490186, 489303, 489447, 
    488551, 487573, 486554, 485089, 486476, 484953, 483570, 484436, 482972, 
    482548, 480729, 481688, 480290, 480615, 479925, 478969, 479209, 478462, 
    478083, 477833, 478505, 476262, 476720, 476405, 475763, 475563, 474970, 
    475215, 474712, 474353, 475453, 474132, 473078, 472842, 474070, 474019, 
    473176, 473351, 473632, 473411, 472183, 473207, 472473, 471853, 472721, 
    472916, 473286, 472715, 472562, 472486, 472721, 473170, 473366, 473849, 
    473912, 473508, 473699, 473554, 473852, 473815, 474036, 474154, 474500, 
    474849, 474457, 475325, 476269, 476749, 477393, 475577, 477007, 477563, 
    477622, 478526, 478397, 478760, 479664, 480019, 481443, 481898, 481663, 
    482115, 482219, 482930, 483743, 483705, 485546, 486141, 486119, 487289, 
    487177, 489612, 489304, 490649, 489886, 491089, 490939, 492562, 494758, 
    494033, 495479, 496056, 497772, 498482, 500587, 499378, 501060, 502276, 
    504148, 503729, 504074, 506835, 506713, 507942, 509437, 511809, 512474, 
    513455, 514265, 516983, 517278, 517484, 519418, 521610, 522611, 524878, 
    526418, 527546, 528733, 530744, 531612, 533494, 536661, 536441, 538521, 
    540828, 542243, 545043, 546959, 548260, 550758, 551805, 554935, 557169, 
    559007, 561513,
  556665, 555271, 552929, 551444, 549844, 545383, 545071, 543992, 540771, 
    541448, 542104, 538752, 536859, 530015, 529519, 529393, 527618, 526860, 
    527113, 526710, 526137, 520903, 520893, 517705, 516863, 515698, 515231, 
    512995, 512787, 511142, 510195, 510806, 509048, 507589, 506091, 503660, 
    504717, 502972, 506039, 501071, 499937, 499697, 498396, 497610, 496560, 
    498225, 493947, 493948, 494852, 492802, 490488, 492030, 490016, 488487, 
    487503, 487890, 486810, 487913, 485207, 484444, 485156, 485198, 482611, 
    485779, 482580, 482814, 484280, 482331, 481715, 481370, 480542, 481018, 
    479228, 478073, 476738, 477354, 476848, 479036, 477919, 477341, 475690, 
    477830, 476788, 475710, 476404, 475664, 476169, 477675, 475970, 475096, 
    477027, 473097, 474121, 474567, 474229, 474655, 476047, 475953, 472792, 
    471815, 474643, 473663, 474975, 476363, 474764, 475633, 474040, 472849, 
    473023, 474515, 477311, 474772, 474923, 477700, 476166, 476378, 477511, 
    475157, 477094, 478100, 478011, 477023, 476525, 478302, 477996, 478270, 
    478845, 479770, 480923, 483316, 482704, 481639, 484372, 483406, 483935, 
    482004, 481306, 484468, 485204, 484771, 485335, 485548, 488230, 488235, 
    488784, 490253, 491139, 489796, 489779, 491871, 494180, 495029, 493385, 
    494640, 496187, 498402, 496177, 497704, 500432, 500369, 499805, 501997, 
    502184, 503068, 505473, 505980, 505221, 507468, 511020, 511825, 512188, 
    513096, 512410, 513977, 518483, 518232, 518606, 519774, 520886, 523848, 
    524327, 523835, 524111, 527618, 530339, 534042, 534324, 535542, 535451, 
    536088, 539095, 541909, 543028, 544468, 547433, 548052, 550592, 552990, 
    554494, 556580,
  552932, 551533, 549052, 547466, 545362, 543915, 543483, 541010, 539335, 
    537221, 535526, 534225, 532986, 531578, 529576, 528700, 526510, 526456, 
    523684, 523673, 522304, 520098, 519001, 518550, 516828, 515460, 513628, 
    512184, 513743, 510054, 510418, 508818, 508336, 505716, 505959, 505205, 
    504610, 502175, 502189, 501494, 500517, 499159, 498538, 497956, 496411, 
    496580, 495831, 494223, 493445, 494224, 492346, 491007, 490950, 489776, 
    489814, 488863, 487845, 488620, 487000, 487310, 486585, 485701, 485680, 
    485499, 484258, 482906, 483956, 483571, 481798, 482336, 481301, 481614, 
    480732, 480970, 480252, 480353, 478803, 479791, 479281, 478787, 477773, 
    477400, 478114, 478801, 477275, 477145, 477608, 477796, 476803, 476405, 
    476189, 476842, 476036, 476617, 476359, 476139, 475058, 477056, 475947, 
    476016, 476852, 475858, 476897, 475887, 475246, 475800, 476185, 477172, 
    476455, 475711, 477400, 477498, 476928, 476932, 477114, 478577, 477692, 
    478553, 478421, 479053, 479198, 478801, 479739, 479399, 479752, 480086, 
    480879, 481899, 480299, 482308, 481354, 482878, 484777, 483003, 483878, 
    484988, 486621, 484942, 485841, 486013, 487196, 486947, 488782, 489020, 
    489693, 489279, 490501, 491559, 492382, 492461, 494018, 492695, 494473, 
    495624, 495570, 496578, 497893, 498762, 499819, 500354, 501413, 502726, 
    502487, 504307, 504656, 505639, 506755, 507901, 508941, 510420, 510706, 
    510991, 513280, 513645, 514676, 515763, 518967, 518673, 519710, 521387, 
    523071, 523643, 525297, 526850, 528051, 529507, 530149, 531612, 533749, 
    535921, 536528, 538817, 540383, 541496, 544066, 544829, 546925, 548962, 
    551085, 552562,
  546477, 544672, 544684, 541236, 538936, 537702, 537052, 538316, 535506, 
    534471, 529756, 527821, 530939, 527095, 525235, 526353, 524439, 522750, 
    523277, 519553, 518685, 519531, 519098, 516122, 513893, 512677, 512988, 
    512033, 509356, 509598, 508569, 507852, 506363, 505663, 504535, 504481, 
    505714, 502460, 502318, 500438, 502003, 501072, 500712, 498160, 497570, 
    495654, 496158, 496691, 494135, 495164, 492568, 493678, 493917, 491765, 
    489311, 490737, 490824, 488360, 488542, 488053, 486720, 484997, 486293, 
    485919, 486542, 483928, 485072, 484735, 482880, 484403, 485213, 483832, 
    484524, 482664, 482073, 481585, 482023, 480794, 480040, 480861, 482511, 
    481675, 481650, 479013, 480313, 481426, 481858, 480739, 479297, 477495, 
    478581, 478683, 479958, 480758, 478805, 478319, 480647, 478027, 477810, 
    477782, 477862, 477692, 479999, 479706, 480152, 477737, 477769, 479112, 
    478558, 479867, 481340, 480755, 477895, 478220, 479769, 480025, 481208, 
    479773, 481253, 480640, 480391, 483819, 482000, 480298, 482296, 481765, 
    482284, 485130, 483710, 482521, 483585, 484256, 484614, 486200, 486315, 
    486699, 487212, 487632, 488251, 488715, 486022, 489778, 490990, 490720, 
    490875, 492407, 490259, 491312, 491813, 494799, 493592, 495223, 497050, 
    495440, 495656, 496706, 497295, 497942, 500212, 503322, 503438, 501215, 
    499674, 503401, 503437, 504207, 508820, 508022, 508082, 506306, 509643, 
    511600, 512747, 513027, 513541, 512819, 515828, 518077, 520154, 517472, 
    519780, 521042, 520656, 525216, 524748, 527285, 526369, 530246, 531714, 
    530010, 529422, 531044, 535408, 539642, 539532, 540533, 541229, 541879, 
    543461, 546672,
  541031, 540280, 538014, 537660, 536277, 534152, 533257, 531277, 531840, 
    529423, 530180, 525929, 525013, 524723, 524077, 522793, 522235, 520300, 
    518080, 518672, 518448, 517324, 515419, 512587, 512766, 513204, 511245, 
    511744, 511348, 507910, 507308, 508808, 506437, 507286, 503691, 504205, 
    502354, 501800, 502837, 501640, 499775, 498757, 499224, 497940, 498348, 
    497732, 498011, 495025, 494916, 493489, 495172, 494035, 493427, 492953, 
    491048, 490746, 490763, 490760, 489026, 489298, 488457, 489047, 489468, 
    488193, 488187, 486417, 486381, 488192, 487391, 486066, 485661, 484262, 
    484355, 483125, 484212, 483976, 484233, 483675, 484439, 482863, 482040, 
    483287, 481687, 484016, 483871, 482213, 480491, 481267, 480367, 481372, 
    480456, 481165, 482156, 480574, 481069, 481434, 478798, 480213, 482101, 
    480402, 480506, 481073, 481070, 481824, 481710, 481809, 481578, 482697, 
    480923, 480658, 480421, 481161, 481376, 481451, 482038, 480805, 482431, 
    483551, 483860, 482793, 482734, 483277, 482961, 484261, 484453, 485781, 
    484316, 484870, 486308, 485126, 487022, 485005, 484089, 488095, 486961, 
    488305, 487684, 489761, 489216, 487885, 490794, 489660, 491028, 492158, 
    490727, 493548, 492182, 493200, 494041, 494802, 493354, 495244, 495538, 
    496831, 497187, 496755, 499627, 499824, 500648, 500230, 500643, 501692, 
    501087, 505236, 504532, 503557, 506997, 505830, 506202, 507716, 509164, 
    508949, 511310, 510687, 512283, 514624, 512964, 515079, 516432, 516752, 
    518937, 519773, 518962, 520164, 523327, 523882, 524006, 523217, 528926, 
    527155, 528321, 530316, 532005, 533074, 535009, 535283, 535577, 538673, 
    539945, 540890,
  536908, 535994, 534529, 533966, 532673, 531199, 530011, 528933, 527537, 
    526337, 526936, 523376, 523729, 522927, 521577, 521651, 518688, 518502, 
    518735, 516533, 515298, 514652, 513931, 513164, 512457, 511481, 510673, 
    510804, 509617, 507808, 507323, 505952, 505907, 504959, 505284, 503387, 
    502652, 503547, 501062, 500473, 500000, 499895, 499416, 499072, 498611, 
    497791, 496593, 496362, 497162, 496309, 494072, 494403, 492720, 493471, 
    492331, 491932, 491810, 491529, 491089, 490673, 490991, 489681, 488974, 
    488641, 488115, 488056, 488492, 487498, 487160, 487718, 487284, 486634, 
    485629, 486265, 485524, 486296, 485397, 483945, 484632, 484615, 484987, 
    484322, 483202, 483629, 483819, 483366, 484291, 483411, 483696, 482334, 
    483406, 482389, 483608, 483152, 481771, 484530, 482299, 482045, 482271, 
    482678, 483610, 482012, 481305, 483127, 483125, 483455, 482884, 483113, 
    482358, 483273, 483357, 483031, 483933, 483892, 482819, 484511, 483228, 
    483655, 484777, 485315, 484876, 484217, 484909, 485126, 485423, 486076, 
    487180, 486021, 487256, 486514, 486253, 486628, 487733, 489064, 488719, 
    489028, 489583, 490971, 489954, 488681, 490562, 491988, 492021, 491178, 
    492649, 492792, 492676, 494803, 495509, 493737, 496261, 494974, 496483, 
    496929, 497048, 498521, 497244, 499646, 499988, 500892, 501547, 501787, 
    503413, 502548, 503098, 503763, 504681, 505841, 507100, 507832, 507723, 
    508035, 510322, 510630, 511236, 512216, 512456, 514086, 514785, 515129, 
    516698, 517272, 517242, 519908, 520382, 520495, 522364, 523223, 523859, 
    524928, 526248, 527889, 528650, 529982, 529781, 532714, 533050, 534119, 
    536062, 536846,
  533684, 532835, 530770, 532078, 528635, 528803, 526788, 526667, 526021, 
    524242, 523223, 522342, 522477, 520638, 518558, 519790, 518095, 516675, 
    516498, 515249, 514877, 512934, 513313, 511845, 511165, 509225, 510628, 
    508547, 509070, 507841, 507302, 506995, 505290, 504659, 504036, 505240, 
    501958, 501145, 502383, 500960, 500705, 500262, 499756, 497532, 499061, 
    497843, 498296, 496200, 496437, 495624, 494984, 494889, 494373, 492405, 
    493030, 493494, 492705, 492544, 491649, 490821, 490830, 491315, 489739, 
    490807, 488509, 491054, 489094, 488869, 488030, 488279, 488080, 487310, 
    487677, 486946, 487133, 487882, 486348, 485715, 486076, 485708, 484862, 
    486265, 484863, 485735, 484463, 485498, 485053, 484209, 484041, 484615, 
    485837, 484844, 483449, 484093, 485408, 483275, 483762, 483877, 484885, 
    482973, 483989, 483818, 484520, 483755, 484164, 483978, 484102, 485170, 
    484241, 483750, 484892, 485194, 485264, 485496, 484450, 485196, 484849, 
    485248, 485001, 485821, 486920, 486507, 486438, 486903, 487332, 487511, 
    486737, 486623, 488443, 487794, 488326, 488048, 489143, 489150, 489368, 
    489172, 490923, 491455, 490129, 490828, 490343, 492214, 493207, 492180, 
    493953, 494544, 492709, 494803, 494299, 494934, 495008, 496505, 496587, 
    497187, 498271, 498588, 499107, 498119, 500956, 500452, 501479, 502301, 
    503533, 502397, 502636, 502903, 505346, 505821, 506058, 506607, 506557, 
    508436, 509462, 509961, 509444, 511360, 510883, 512769, 512874, 514016, 
    515513, 515688, 517001, 518034, 518280, 518918, 520373, 521513, 521821, 
    522581, 524637, 524823, 525985, 526373, 528559, 529237, 530389, 531180, 
    532493, 533645,
  532584, 531926, 531147, 530561, 528803, 527492, 526675, 526462, 524715, 
    523667, 522844, 522023, 520619, 520635, 519072, 519095, 517252, 516335, 
    517486, 513933, 515475, 513072, 512269, 511864, 510543, 509668, 510306, 
    509166, 508367, 507517, 506981, 506885, 504949, 503809, 504822, 503696, 
    502274, 502837, 502109, 500880, 499592, 500078, 499566, 498499, 499183, 
    496625, 497014, 497655, 495973, 496017, 495962, 494750, 494390, 494266, 
    492964, 493072, 492579, 492939, 492060, 491787, 490639, 490328, 490385, 
    490795, 490062, 489670, 490700, 489563, 488504, 488625, 488643, 487907, 
    487439, 486857, 487029, 486238, 487635, 486123, 485658, 486685, 485425, 
    485797, 485412, 485339, 486101, 485784, 485421, 483984, 484985, 485043, 
    484830, 484670, 484315, 484561, 485227, 484383, 484559, 483781, 484992, 
    483788, 484326, 485195, 484470, 484681, 483975, 483458, 485822, 484543, 
    484232, 484583, 484600, 485334, 485411, 485629, 484457, 487743, 485126, 
    486088, 485304, 485265, 485812, 486131, 486609, 486816, 487209, 487319, 
    488492, 487486, 488249, 488310, 488094, 488000, 489595, 488893, 490084, 
    490015, 489863, 491453, 491198, 491178, 491986, 491789, 492962, 492660, 
    494140, 492772, 494436, 494312, 495337, 495766, 496293, 495890, 497382, 
    496852, 498115, 497788, 498518, 499498, 500537, 500541, 499741, 501563, 
    502294, 503245, 504025, 503717, 504426, 505416, 505976, 506492, 507447, 
    507305, 509340, 509269, 510242, 510422, 511800, 512059, 512829, 514110, 
    515069, 514950, 516660, 516589, 517588, 518807, 521027, 520817, 521190, 
    523318, 522743, 524021, 525663, 526810, 527802, 528232, 529200, 530127, 
    532627, 532751,
  532170, 531459, 529952, 529384, 527983, 528023, 525687, 525933, 524470, 
    522850, 522443, 521605, 520887, 519479, 519005, 518507, 517541, 515857, 
    515548, 514477, 514169, 514564, 511658, 510860, 511082, 510091, 510508, 
    508277, 507836, 506401, 507606, 505532, 506301, 504556, 503970, 502483, 
    502817, 503271, 500981, 501401, 500672, 500089, 499847, 498826, 498132, 
    497845, 496979, 498702, 495913, 495630, 494443, 496152, 494639, 493268, 
    494145, 492589, 493075, 492805, 491728, 492770, 491522, 491449, 490956, 
    490420, 488642, 489178, 490217, 488804, 488356, 489686, 488575, 488087, 
    487746, 487161, 487689, 487906, 486764, 488107, 485780, 486396, 486353, 
    485702, 485812, 485914, 486631, 486009, 485697, 484725, 484605, 484968, 
    485259, 484670, 484910, 484728, 484413, 484469, 484803, 486007, 484287, 
    484884, 484629, 484539, 484987, 485185, 484604, 484534, 484905, 484141, 
    485303, 484690, 484653, 486006, 484970, 485679, 486637, 485710, 485193, 
    486327, 487593, 485947, 485957, 486500, 487276, 486679, 487966, 487660, 
    486753, 487317, 488162, 489189, 489401, 488950, 488581, 490181, 489778, 
    490448, 491279, 491044, 490488, 492884, 491169, 493020, 491984, 493961, 
    493324, 493683, 493740, 494179, 494840, 495273, 495838, 496249, 497377, 
    498579, 497572, 498613, 498982, 499175, 499696, 500089, 500770, 501893, 
    501144, 503572, 502505, 505103, 504391, 504607, 506007, 507645, 506916, 
    506531, 508406, 510086, 509510, 510949, 511484, 511173, 513216, 513140, 
    513786, 515812, 516649, 516300, 517566, 518230, 520219, 519672, 521868, 
    522626, 522863, 523107, 524493, 526326, 527368, 527804, 528773, 529897, 
    530971, 532393,
  530927, 530149, 528940, 528125, 526705, 526654, 525048, 524112, 523479, 
    522850, 521508, 520350, 520086, 519102, 517389, 517942, 516412, 516884, 
    513711, 514938, 513898, 512484, 511648, 511226, 510579, 510431, 509084, 
    508183, 507512, 507338, 505441, 505226, 505357, 504833, 504511, 503133, 
    503379, 502252, 500587, 501694, 500955, 500490, 499137, 498216, 498587, 
    497970, 496736, 497962, 496888, 495149, 496240, 494200, 495451, 495738, 
    494766, 493522, 493181, 492223, 491202, 492535, 491509, 490888, 491716, 
    491809, 489758, 490233, 490230, 491433, 488305, 488826, 488419, 488478, 
    488051, 488291, 487781, 488521, 487193, 486760, 487970, 487034, 487050, 
    486983, 486464, 486354, 485845, 486213, 485835, 484930, 484915, 486426, 
    485377, 485493, 485683, 485554, 486151, 486085, 484353, 485345, 485151, 
    485968, 485884, 484245, 484469, 486609, 485413, 485590, 484770, 485110, 
    485780, 486465, 485786, 486149, 485452, 485207, 487014, 486279, 486422, 
    485996, 486513, 486719, 487728, 486116, 486705, 487990, 488796, 488415, 
    487776, 488865, 488629, 488759, 490249, 489654, 489705, 490744, 490276, 
    489278, 490790, 490714, 491302, 491266, 493541, 493661, 493074, 492425, 
    493596, 494349, 494643, 495526, 494510, 495954, 495668, 497429, 496873, 
    496908, 497842, 499262, 498335, 500060, 499975, 500692, 499947, 500821, 
    502757, 501873, 503740, 504516, 503880, 505558, 505801, 505204, 507217, 
    506522, 508986, 509229, 509042, 509713, 512134, 511233, 512276, 513363, 
    513449, 514759, 515788, 515300, 516753, 519069, 518020, 519340, 519939, 
    522382, 521239, 522717, 523792, 525103, 526175, 526407, 527897, 528535, 
    530128, 530808,
  528708, 527836, 526807, 525620, 525195, 524352, 522851, 522722, 522262, 
    521050, 518208, 520052, 518679, 517712, 517016, 516247, 515216, 515132, 
    513610, 513133, 512284, 511455, 511534, 510630, 509650, 508391, 508589, 
    508266, 507726, 506626, 506399, 505175, 504917, 503904, 503056, 503105, 
    503485, 501663, 502476, 500667, 500416, 499934, 498254, 499761, 498300, 
    498208, 497866, 497114, 497950, 497556, 495414, 495875, 495241, 494684, 
    493765, 493853, 493505, 493084, 493134, 494087, 491058, 492742, 492696, 
    491383, 491557, 491159, 490558, 490309, 489326, 489729, 489563, 489697, 
    488722, 488461, 489023, 488665, 488516, 488275, 488265, 488069, 487755, 
    488514, 487292, 486986, 486643, 487971, 487071, 487083, 487075, 485955, 
    486964, 486784, 485807, 486695, 486198, 486431, 486331, 487448, 486335, 
    484999, 486395, 487091, 485673, 486167, 486983, 486908, 486361, 485511, 
    487423, 487067, 486064, 487011, 486851, 486191, 487288, 485945, 488257, 
    487428, 488050, 488364, 488049, 488153, 487841, 488681, 489183, 489420, 
    488531, 489121, 489576, 489947, 489980, 489985, 490401, 490515, 491758, 
    491421, 491524, 491894, 491867, 492279, 492942, 492763, 493019, 493793, 
    494680, 495046, 494998, 494780, 495260, 496644, 496700, 496449, 497334, 
    497950, 498050, 498230, 500077, 498809, 499422, 501158, 500358, 500810, 
    501593, 502666, 503895, 503693, 504547, 504780, 505087, 505338, 506382, 
    507938, 506575, 509074, 508108, 509417, 508952, 511318, 512152, 512434, 
    512335, 514586, 513054, 515176, 515997, 516411, 516970, 518054, 519430, 
    519357, 520491, 521493, 521788, 522622, 524296, 524832, 525421, 526722, 
    527601, 528471,
  526541, 526025, 524965, 522672, 524214, 523658, 522574, 518304, 518827, 
    521172, 521638, 516682, 515397, 514218, 517592, 517040, 517499, 513130, 
    510992, 510236, 511333, 510467, 511198, 509892, 508654, 508533, 507343, 
    507730, 507109, 505322, 506468, 506923, 502966, 501766, 504481, 503351, 
    505319, 503259, 503796, 501075, 499434, 498418, 497991, 499456, 498299, 
    495773, 499625, 498177, 498570, 495733, 494861, 495495, 496624, 495558, 
    495223, 495978, 495907, 493577, 494673, 494653, 493147, 491106, 489373, 
    491197, 491047, 492078, 491307, 492269, 491158, 489750, 489471, 489214, 
    490168, 488510, 488328, 490030, 489979, 488511, 489018, 488111, 489734, 
    487787, 487733, 488168, 488231, 487272, 487568, 488402, 490473, 489627, 
    489721, 488257, 484930, 487563, 485927, 486129, 488994, 488047, 489093, 
    487318, 489059, 486415, 484462, 485039, 484851, 487327, 486112, 488085, 
    489975, 484831, 485854, 486929, 486671, 488710, 486957, 491690, 490722, 
    489072, 491695, 489167, 489209, 489158, 488208, 488652, 487860, 491241, 
    489390, 490042, 491555, 486301, 491007, 489334, 490745, 491476, 493420, 
    492476, 489534, 491638, 493491, 493322, 494136, 492548, 492390, 495300, 
    497274, 495057, 495429, 496285, 491600, 494878, 496767, 500631, 499372, 
    500395, 497914, 500215, 501357, 497097, 498481, 497208, 498712, 499961, 
    502116, 503740, 506024, 505416, 504687, 504372, 502402, 501439, 503663, 
    505675, 510077, 512678, 510281, 508378, 505815, 506885, 506567, 512988, 
    513647, 514621, 516141, 518850, 513356, 512155, 514790, 516667, 515232, 
    518694, 521517, 522521, 518687, 516215, 524554, 525793, 523761, 523941, 
    525034, 526799,
  525083, 523820, 523183, 522653, 521924, 521310, 519775, 519562, 519245, 
    517927, 516940, 517838, 514529, 516207, 515048, 513387, 513797, 513216, 
    511576, 511302, 511301, 510592, 509239, 509485, 508628, 508102, 506796, 
    507080, 507417, 505879, 505190, 504566, 504233, 504057, 502033, 503430, 
    502771, 502366, 500705, 500745, 501377, 499796, 499702, 498692, 499631, 
    497923, 497677, 497474, 497970, 497317, 496788, 495803, 496430, 495392, 
    496079, 494841, 493689, 493991, 493763, 492989, 493722, 493324, 492772, 
    492557, 492744, 492472, 491979, 492521, 490322, 490829, 490872, 490438, 
    490323, 490952, 490686, 489890, 490306, 488748, 489743, 489953, 488402, 
    488278, 490492, 490085, 489158, 488831, 487298, 488531, 488465, 488069, 
    489007, 488124, 487142, 488753, 486939, 489452, 487426, 488439, 487541, 
    488870, 487521, 488338, 487212, 487416, 488433, 487610, 488331, 488037, 
    489773, 488779, 487755, 488432, 488335, 489303, 489137, 488563, 488686, 
    489978, 488530, 489520, 489470, 490325, 489526, 489495, 489164, 491043, 
    491232, 490489, 490188, 491597, 491222, 491054, 491881, 491006, 492331, 
    493685, 492581, 491364, 492418, 494302, 494241, 494786, 493984, 494097, 
    496480, 494400, 495755, 495785, 496165, 496194, 495898, 498647, 497479, 
    498105, 498639, 498695, 499022, 499742, 499753, 499268, 500614, 502512, 
    501777, 502528, 502722, 502747, 503396, 504804, 504256, 504766, 506424, 
    506329, 505335, 507556, 507622, 508111, 509369, 509506, 510597, 510143, 
    510509, 512109, 513238, 512818, 513458, 514461, 515449, 515192, 516666, 
    517012, 517933, 518558, 519368, 519761, 521021, 521622, 522049, 522964, 
    524016, 524768,
  522588, 521770, 521230, 520457, 520068, 519163, 518453, 517723, 517456, 
    516673, 515479, 515601, 514394, 514019, 514565, 511990, 511869, 511977, 
    511023, 510555, 510196, 510115, 508586, 507756, 507534, 508188, 506314, 
    507669, 505531, 505246, 505305, 503517, 504410, 502812, 502729, 502994, 
    502911, 501135, 501464, 500513, 500508, 498806, 500034, 499847, 500056, 
    499018, 497928, 497411, 497393, 497513, 496276, 496860, 496425, 496363, 
    496074, 495390, 494389, 496287, 493601, 494159, 492601, 494382, 493277, 
    493460, 493525, 492498, 492963, 492151, 490822, 491884, 492352, 491381, 
    491835, 491660, 491786, 491496, 489419, 489417, 492395, 490504, 490361, 
    489875, 490140, 489706, 489198, 489182, 489561, 490014, 489168, 488715, 
    489171, 489548, 489714, 488855, 490014, 489047, 488496, 489106, 488847, 
    488552, 488657, 488602, 489683, 490016, 489348, 488355, 489244, 489845, 
    489217, 488568, 489625, 488591, 489850, 489113, 490732, 490222, 490965, 
    489447, 489836, 489498, 489928, 491618, 490405, 491162, 491135, 490886, 
    491564, 491261, 490887, 491772, 492175, 493259, 492268, 492251, 492435, 
    493837, 493272, 492056, 494794, 494004, 494729, 494887, 494037, 495402, 
    495479, 495428, 496439, 495942, 496536, 497280, 497012, 497818, 497557, 
    497743, 498222, 499411, 499607, 499182, 500042, 500486, 501260, 499809, 
    502575, 502743, 501373, 503584, 502628, 504403, 503093, 504921, 505600, 
    505770, 506048, 506534, 507613, 506664, 508654, 508999, 508609, 509918, 
    509768, 511306, 511333, 512591, 512311, 513146, 514048, 513436, 515671, 
    515255, 516490, 516638, 517571, 518480, 519166, 518857, 520943, 520806, 
    521839, 522530,
  521956, 521236, 519974, 521362, 519646, 516684, 518165, 517571, 517005, 
    516576, 514497, 517009, 513505, 512743, 513733, 512347, 510364, 511832, 
    512094, 509339, 509223, 510531, 509627, 507968, 506132, 507731, 507729, 
    506665, 504876, 504227, 504851, 505215, 504138, 503764, 501781, 501611, 
    502122, 500610, 502028, 502292, 499830, 499188, 500883, 499516, 497956, 
    497991, 499132, 498267, 497759, 497551, 497136, 497217, 497885, 495048, 
    495937, 494967, 492551, 495320, 495472, 495710, 494326, 493436, 493765, 
    493341, 491324, 492784, 492632, 494122, 493431, 491612, 490928, 491666, 
    492582, 490737, 491354, 492630, 491293, 489394, 489798, 491601, 491505, 
    490431, 490852, 489708, 490046, 490520, 488912, 489058, 491031, 489318, 
    490301, 489953, 489020, 487962, 488719, 490654, 488770, 488631, 488966, 
    488945, 488193, 490412, 487359, 490074, 489888, 489413, 490233, 490899, 
    488454, 490286, 489857, 489081, 490213, 488737, 491297, 490256, 491212, 
    492015, 491546, 490220, 490040, 489346, 490058, 491995, 491876, 489164, 
    490823, 490252, 492743, 491733, 492765, 492140, 493586, 493358, 492252, 
    495017, 493826, 493323, 494617, 494590, 494852, 494625, 494541, 494384, 
    496968, 494671, 494201, 497698, 494782, 496554, 498918, 497547, 498250, 
    498902, 497580, 498824, 500283, 498886, 500842, 502581, 501131, 500061, 
    499866, 502388, 502388, 500713, 504037, 502326, 504739, 505533, 506355, 
    506893, 505643, 506412, 504997, 508703, 507528, 507961, 508853, 508858, 
    509864, 509687, 511353, 512297, 513859, 511683, 511089, 516340, 514938, 
    515205, 515569, 515795, 515942, 520260, 517145, 518672, 520385, 520672, 
    520897, 521791,
  519744, 518995, 518495, 517774, 517887, 516514, 515524, 515654, 515432, 
    514675, 512514, 514190, 512841, 512634, 512098, 510156, 511284, 509792, 
    509562, 508952, 509163, 509245, 507441, 506674, 507787, 506546, 505212, 
    505174, 505920, 503940, 504133, 503806, 503242, 503975, 502247, 502589, 
    501621, 501126, 500983, 501253, 500084, 500558, 500226, 499971, 498752, 
    499113, 497827, 499069, 497901, 498031, 496440, 496465, 496727, 496378, 
    496359, 495729, 496687, 495611, 493541, 494572, 494758, 495974, 493855, 
    494317, 494222, 493976, 492764, 494247, 493193, 491735, 493324, 492837, 
    493200, 492722, 491333, 491797, 491886, 491352, 492926, 490698, 491730, 
    491701, 491294, 491008, 491338, 490276, 490612, 491028, 490385, 490368, 
    490220, 490471, 490618, 490089, 492102, 489570, 491298, 489470, 490945, 
    490717, 490556, 490553, 490175, 490459, 489013, 490917, 490575, 490995, 
    490560, 490529, 491463, 490483, 491839, 489740, 491057, 491967, 489891, 
    491451, 490925, 490838, 492185, 491655, 493225, 492055, 491556, 491348, 
    491921, 492982, 492733, 493346, 493293, 491914, 492981, 495222, 494330, 
    493525, 493994, 493899, 495539, 495043, 494693, 495340, 494821, 495385, 
    495277, 497224, 496456, 496563, 496567, 498189, 497629, 497932, 497384, 
    497676, 499115, 499847, 499455, 500197, 499908, 499311, 501578, 501218, 
    500694, 502249, 502570, 502001, 502548, 504651, 503059, 504484, 504094, 
    505293, 505045, 505559, 507095, 507401, 506046, 508055, 507539, 508819, 
    507570, 510717, 509919, 510818, 510285, 511903, 512152, 512894, 512314, 
    513456, 515300, 513752, 516021, 516043, 516047, 517570, 517293, 518271, 
    519327, 519457,
  518589, 518274, 517799, 516951, 516569, 515944, 515361, 514341, 514056, 
    513680, 513861, 512674, 512312, 511509, 510901, 510452, 510521, 509408, 
    509870, 508696, 507993, 508374, 507603, 507225, 506531, 505896, 504890, 
    506112, 503991, 504987, 503873, 504215, 502743, 503490, 502196, 502832, 
    500585, 502544, 500776, 500335, 500675, 500405, 499999, 499736, 498469, 
    498402, 498409, 499134, 498375, 497200, 497780, 497001, 496650, 496196, 
    496989, 496506, 495637, 495556, 495161, 494696, 495473, 495148, 493790, 
    495211, 494297, 494404, 493144, 493582, 493170, 493368, 493549, 493473, 
    492792, 492001, 491905, 492278, 492529, 491855, 492374, 491917, 492160, 
    492414, 491978, 491805, 490832, 490813, 492183, 491207, 491685, 490687, 
    491190, 489913, 491080, 490796, 490946, 491183, 491223, 490272, 490953, 
    490477, 491237, 490391, 491186, 490595, 491367, 491338, 490440, 491631, 
    489908, 492601, 491287, 490960, 491109, 490194, 491859, 491218, 491680, 
    492467, 490928, 492257, 492214, 491887, 492812, 493326, 491607, 493088, 
    492679, 493136, 492995, 492410, 492870, 493072, 493926, 494170, 494565, 
    493868, 494030, 494613, 495221, 495500, 495193, 494761, 496090, 495379, 
    496042, 496010, 496923, 497321, 496872, 497529, 497921, 498461, 498118, 
    498194, 498801, 499034, 499063, 499472, 500301, 500909, 501748, 501274, 
    500654, 501142, 502812, 501651, 502029, 503375, 503865, 504744, 503306, 
    504779, 505479, 505390, 506222, 507025, 506895, 506144, 508737, 507468, 
    508418, 508875, 509900, 509604, 511398, 510830, 511032, 511870, 512371, 
    513618, 513105, 514634, 514559, 515193, 515371, 516402, 517009, 517328, 
    518180, 518535,
  517832, 517356, 517193, 515621, 515477, 515251, 514895, 514236, 512634, 
    514124, 512025, 513303, 511226, 512486, 508972, 510074, 509633, 509634, 
    508543, 508529, 506867, 509135, 506377, 506923, 506401, 505905, 505052, 
    505291, 504076, 504247, 504395, 503683, 502645, 503479, 501848, 502843, 
    501744, 501324, 501005, 501194, 499437, 499848, 499033, 500449, 499086, 
    499645, 498150, 497843, 499123, 497729, 496834, 498472, 496393, 497736, 
    496737, 496170, 495581, 497025, 495367, 494867, 494524, 494227, 494983, 
    495268, 496628, 493342, 493894, 493596, 493557, 493575, 492209, 493560, 
    493546, 493009, 493222, 492621, 492566, 492701, 493995, 491575, 491044, 
    492001, 491688, 492583, 490572, 491921, 493225, 491411, 491377, 492643, 
    490433, 491936, 491962, 490168, 491038, 492780, 491090, 490364, 492041, 
    491267, 490827, 491434, 491081, 490956, 492779, 490201, 491155, 491086, 
    491690, 492216, 491647, 492227, 491309, 491878, 491117, 491924, 491612, 
    492350, 491863, 491817, 491146, 492366, 492840, 493316, 493306, 492897, 
    492994, 493287, 494123, 492569, 494084, 493762, 493941, 493839, 494786, 
    494665, 494509, 494624, 495091, 494400, 495503, 495249, 496570, 497106, 
    495392, 496816, 496973, 496213, 497766, 497494, 498093, 499396, 497783, 
    498566, 497948, 498991, 499182, 499663, 499665, 502390, 500377, 500778, 
    501222, 502323, 501774, 502192, 502605, 502548, 503550, 503847, 503918, 
    503786, 505051, 505734, 505901, 506503, 506900, 505848, 508280, 507026, 
    508470, 508033, 509415, 509161, 510754, 510571, 510372, 512566, 511143, 
    513144, 511784, 513932, 513745, 515010, 514301, 516508, 515719, 516548, 
    517275, 517767,
  517415, 516919, 517252, 515466, 514670, 513346, 514191, 515294, 517234, 
    509894, 512965, 507389, 509922, 516213, 511732, 508548, 510458, 510994, 
    507523, 506666, 506793, 508188, 504431, 505839, 509406, 506334, 505765, 
    504214, 503266, 500131, 503124, 505303, 505005, 504220, 503408, 503637, 
    498873, 498761, 501280, 500271, 502153, 501665, 501552, 500525, 497605, 
    499358, 497852, 495622, 498487, 497416, 502055, 497440, 497586, 494931, 
    495084, 494386, 495845, 498338, 494539, 497778, 497403, 494953, 493764, 
    494212, 492701, 495827, 497354, 494038, 492072, 492270, 493266, 494054, 
    492540, 493543, 493190, 493784, 491799, 493025, 490390, 491951, 494836, 
    492031, 491606, 492029, 494033, 495010, 489997, 490868, 491385, 491571, 
    490690, 490974, 492854, 492229, 490980, 493713, 489044, 491233, 490372, 
    491217, 491105, 491751, 489799, 489520, 492591, 492401, 492026, 492607, 
    492553, 491849, 493448, 491528, 490234, 492774, 491876, 493972, 491397, 
    490808, 491298, 492081, 493793, 490821, 493594, 491200, 492628, 493801, 
    494468, 492366, 494583, 493909, 493310, 494749, 496527, 494996, 496163, 
    493344, 492529, 492124, 495753, 500760, 496509, 490405, 494559, 497784, 
    499413, 497909, 495963, 492917, 495906, 496095, 498359, 499041, 499037, 
    498941, 498803, 496776, 502235, 502468, 500007, 496591, 499692, 500409, 
    499774, 506147, 506077, 502445, 501713, 500905, 500212, 504098, 507080, 
    506909, 503620, 502452, 504305, 505864, 505498, 507748, 509922, 506944, 
    506663, 509695, 508351, 509428, 508603, 510562, 511511, 514539, 509849, 
    510385, 511393, 515267, 515608, 510904, 514943, 515625, 516491, 516743, 
    516256, 517250,
  516355, 515678, 515245, 515193, 514282, 513758, 513106, 513483, 512368, 
    512093, 511902, 510136, 510639, 510535, 510125, 508750, 509399, 508862, 
    508193, 507311, 506649, 507489, 506470, 505197, 506078, 505939, 504323, 
    504995, 504835, 504315, 502979, 503537, 502873, 502103, 501832, 502097, 
    501342, 502121, 500362, 500883, 500459, 499985, 500401, 499924, 499553, 
    497918, 498625, 498431, 498367, 498859, 497167, 497395, 497129, 497102, 
    496362, 496954, 496898, 496686, 495069, 495835, 495462, 496715, 494299, 
    494378, 495532, 494722, 494741, 494872, 494466, 493950, 493993, 493230, 
    494109, 493221, 493571, 493581, 493042, 493436, 492825, 494615, 492591, 
    492271, 492084, 492393, 492395, 493240, 492314, 492992, 491991, 491775, 
    492400, 491873, 491578, 492780, 491912, 491722, 492794, 492045, 491209, 
    492132, 492842, 491896, 490328, 492456, 491311, 492486, 492030, 493077, 
    492752, 491633, 492134, 492345, 492606, 491853, 492236, 492424, 493136, 
    492109, 492915, 494012, 492353, 492509, 493446, 493346, 493276, 493529, 
    493525, 494419, 493984, 493081, 494275, 494695, 494052, 494562, 494895, 
    495743, 495297, 495050, 495412, 495148, 495225, 496114, 496386, 497130, 
    496437, 496052, 497044, 497646, 497090, 497644, 499096, 498349, 497917, 
    497993, 500315, 498716, 500099, 499804, 499270, 500390, 501029, 499603, 
    501905, 502014, 501865, 502432, 502481, 502843, 502632, 503242, 503281, 
    505452, 504070, 504152, 506084, 505140, 506951, 506194, 506710, 506552, 
    508326, 507316, 508393, 508926, 509292, 509591, 510076, 510304, 511451, 
    511283, 511843, 512057, 512723, 513577, 513672, 514273, 515000, 515005, 
    516116, 516046,
  515714, 515119, 514607, 514238, 514057, 513443, 512773, 512392, 511044, 
    512086, 511354, 509595, 511313, 510110, 508949, 508218, 508945, 508502, 
    507616, 507518, 506780, 506258, 506360, 506130, 505193, 505093, 505291, 
    504493, 503740, 503520, 503972, 502380, 503000, 502288, 502013, 503166, 
    501227, 501295, 500853, 500473, 499566, 500375, 499843, 500324, 499648, 
    498603, 499323, 497321, 499020, 497857, 496870, 499113, 497885, 496675, 
    496906, 495987, 497080, 496128, 497575, 495624, 495272, 495474, 496022, 
    494807, 494329, 496104, 494324, 494750, 495222, 495054, 493237, 493416, 
    493716, 494360, 493516, 494804, 492461, 493325, 493710, 493348, 493283, 
    493072, 492465, 493526, 491752, 494455, 491380, 492157, 492795, 493519, 
    492119, 493281, 492494, 491950, 491818, 491689, 492986, 492203, 493207, 
    492169, 491765, 491873, 492978, 492392, 493336, 492198, 491458, 492698, 
    493250, 492113, 491302, 492772, 491670, 494180, 493079, 492449, 492854, 
    492253, 493098, 492416, 493261, 493633, 494371, 493884, 494380, 493113, 
    493547, 494621, 493722, 493873, 494511, 494364, 494308, 495768, 494169, 
    495609, 494009, 495946, 496652, 495498, 496401, 496371, 495360, 496986, 
    496015, 497391, 497357, 496962, 497618, 497307, 499254, 498312, 498618, 
    499713, 498075, 499708, 499875, 498645, 499613, 500874, 500602, 501558, 
    501158, 500650, 502266, 502031, 502421, 502935, 503047, 503291, 502962, 
    504424, 504647, 504153, 505165, 505225, 505761, 506583, 506315, 506307, 
    507936, 507523, 507895, 509412, 507948, 509582, 510289, 509015, 511252, 
    510289, 511142, 512378, 512168, 512859, 513500, 513503, 514311, 514852, 
    514720, 515684,
  513024, 512242, 512854, 512225, 510531, 510858, 511093, 510544, 508845, 
    510448, 509522, 509582, 505024, 508838, 509082, 508722, 505258, 506955, 
    506420, 506867, 505028, 505397, 505707, 507201, 503727, 503937, 503332, 
    504338, 501391, 502322, 504964, 502109, 503180, 500373, 501273, 502069, 
    502559, 499816, 501117, 500373, 500512, 499941, 499996, 499722, 499351, 
    500271, 497839, 498942, 500903, 497102, 496776, 499261, 498118, 496516, 
    499483, 497590, 494691, 498503, 498386, 495492, 494872, 496320, 496482, 
    497027, 495357, 496093, 495110, 495540, 495961, 497338, 493960, 493515, 
    494953, 495665, 496000, 491837, 494318, 495291, 493886, 495075, 494554, 
    495068, 493664, 495444, 493752, 494369, 493018, 494158, 494021, 492306, 
    495188, 492791, 491721, 495627, 494585, 491725, 493061, 494836, 493477, 
    493331, 495142, 493999, 493705, 494272, 490547, 491947, 495517, 495234, 
    492194, 495126, 494913, 493707, 494220, 493788, 495450, 493349, 493299, 
    494807, 494921, 494629, 493322, 493948, 493414, 492966, 494764, 495986, 
    495322, 492711, 494489, 496943, 495529, 496473, 494415, 496812, 495952, 
    494525, 495856, 495931, 497918, 496264, 497959, 495945, 497421, 496110, 
    496361, 497133, 498096, 496584, 501164, 498549, 497932, 499013, 498180, 
    499309, 499366, 497977, 499538, 499055, 498707, 500819, 502805, 498196, 
    501594, 502947, 500425, 501611, 502879, 501232, 502343, 504377, 504053, 
    500209, 506770, 503914, 502713, 506847, 503556, 503667, 503533, 508344, 
    507511, 505692, 505610, 509620, 506394, 505116, 510658, 509227, 507138, 
    508372, 509632, 511223, 508774, 512357, 511199, 509258, 513314, 512705, 
    511825, 512997,
  511262, 510608, 510509, 509793, 509973, 509508, 509131, 509278, 507735, 
    508928, 507342, 507417, 507170, 507275, 506664, 506700, 505749, 505334, 
    505616, 505156, 504707, 505017, 504223, 503826, 504864, 503832, 502695, 
    503993, 502258, 502406, 503100, 502213, 501171, 502189, 501482, 501320, 
    501030, 500620, 500821, 500534, 500991, 499685, 499593, 499651, 499227, 
    500006, 498771, 498788, 499307, 497898, 498437, 498139, 498928, 497887, 
    497503, 498765, 497265, 497143, 498121, 496730, 496323, 497104, 495902, 
    497104, 496388, 496010, 497263, 496408, 495827, 496933, 494890, 495005, 
    496508, 496203, 495038, 495821, 495885, 494692, 495525, 494402, 495377, 
    494738, 495115, 495258, 495532, 494902, 494527, 493909, 495101, 494918, 
    494098, 494838, 495404, 493934, 494189, 494483, 494662, 493955, 494622, 
    494923, 494676, 494400, 494562, 493990, 495271, 494635, 494564, 495164, 
    493415, 494715, 493942, 494262, 495485, 495347, 494793, 495054, 495233, 
    495192, 495075, 494237, 494598, 496419, 494933, 495553, 494695, 496378, 
    494878, 495903, 494887, 495943, 495783, 495947, 497680, 495119, 496720, 
    496740, 497105, 495374, 497971, 496724, 497535, 496781, 497419, 497240, 
    497535, 498177, 497427, 498734, 498892, 498298, 498758, 498422, 498759, 
    499038, 499894, 498493, 499870, 499414, 500162, 501508, 500277, 500948, 
    500160, 500934, 501635, 501600, 501772, 501666, 502360, 502735, 502648, 
    503040, 502997, 503029, 504090, 503739, 504193, 504992, 504423, 504730, 
    505220, 505889, 505340, 506382, 505867, 507002, 507025, 507284, 507563, 
    508401, 507491, 509051, 508565, 509430, 509323, 510124, 509945, 510546, 
    510797, 511068,
  509800, 509364, 509085, 509241, 508335, 508151, 508058, 507489, 507228, 
    507960, 506223, 506390, 506500, 506407, 505439, 505457, 505201, 505309, 
    505004, 504022, 504389, 504544, 504016, 503416, 503401, 503009, 503253, 
    503109, 501560, 502606, 501297, 502656, 501804, 501837, 500781, 501235, 
    500902, 500996, 500783, 500627, 499652, 500813, 499189, 499168, 499951, 
    499800, 498979, 499060, 500105, 498015, 498336, 499410, 497573, 497899, 
    498769, 497913, 496936, 498067, 497471, 498268, 496645, 497784, 497846, 
    496967, 495655, 496681, 497113, 497351, 495884, 496985, 496800, 495799, 
    496948, 495912, 496049, 496559, 495068, 495565, 496369, 495628, 495368, 
    495912, 495180, 496419, 495301, 495345, 495629, 494581, 494523, 495961, 
    495556, 495800, 495084, 495290, 495653, 494659, 495465, 495784, 495388, 
    494523, 494414, 494591, 495727, 495451, 495523, 495050, 494594, 495988, 
    494528, 495850, 494521, 496912, 494121, 496094, 495326, 495088, 495170, 
    495671, 495570, 495728, 495787, 495604, 495743, 496435, 495801, 496578, 
    496632, 495820, 495775, 496712, 496244, 496362, 497095, 496267, 496106, 
    497431, 497583, 498047, 496631, 497457, 497153, 497478, 497768, 497825, 
    497696, 497481, 499299, 497951, 498554, 498573, 499496, 499084, 499313, 
    498376, 499840, 499821, 499683, 500202, 499661, 500694, 499956, 499489, 
    501944, 500892, 501678, 501045, 501193, 502068, 502340, 501844, 502122, 
    502421, 503550, 503138, 502857, 503470, 503775, 503667, 504605, 504000, 
    505550, 504536, 504899, 505048, 505644, 506163, 506597, 506077, 506933, 
    506694, 506933, 507983, 507290, 508205, 508505, 508365, 508861, 509176, 
    509386, 509838,
  508590, 508542, 508124, 506334, 508961, 507093, 508304, 507608, 507483, 
    502900, 501650, 509568, 506444, 508394, 508404, 499594, 505589, 500925, 
    503898, 502405, 508154, 504775, 504620, 503791, 504466, 497223, 502553, 
    501894, 506279, 501325, 503835, 501388, 496827, 497100, 502220, 502147, 
    504604, 502763, 498329, 499773, 498362, 498978, 501806, 498890, 501060, 
    501301, 499142, 499646, 500645, 494710, 498869, 499918, 501023, 497560, 
    496564, 500075, 498611, 499031, 497443, 496126, 496043, 497603, 494772, 
    498281, 498938, 499396, 492910, 498129, 494876, 497262, 498454, 500493, 
    497050, 494058, 496850, 496755, 495070, 498084, 498746, 496068, 491827, 
    496178, 495838, 496358, 497590, 496259, 493596, 494637, 496009, 497981, 
    496311, 494649, 493292, 494636, 497559, 497717, 497036, 497233, 493594, 
    492819, 495840, 497291, 496167, 496311, 496009, 493591, 493743, 497487, 
    496315, 495834, 500956, 492850, 492484, 495009, 494940, 495668, 499073, 
    498347, 495216, 494401, 495816, 496553, 496302, 498912, 498535, 496102, 
    492525, 493776, 497294, 499073, 497561, 495514, 498497, 496815, 495587, 
    500981, 496258, 495671, 496381, 499130, 498390, 497443, 500969, 499730, 
    498873, 497703, 495920, 497354, 497256, 498440, 501687, 499565, 497093, 
    497850, 500701, 501043, 502712, 498801, 498824, 496850, 499071, 502996, 
    507804, 501541, 501090, 496844, 493950, 501583, 505613, 504572, 506089, 
    504656, 497057, 497268, 500402, 508066, 507080, 508008, 500867, 498644, 
    498359, 510864, 506419, 508027, 500998, 504032, 508150, 507445, 501001, 
    507565, 505777, 508870, 506143, 508812, 506116, 506940, 509007, 507406, 
    508471, 508784,
  507861, 507372, 507328, 506936, 506847, 506710, 506010, 506783, 505788, 
    505380, 505349, 505290, 504710, 505218, 504399, 504422, 504174, 504553, 
    503545, 503734, 502692, 503613, 503791, 502445, 503129, 501746, 502640, 
    502532, 501754, 501631, 502029, 501149, 501590, 501601, 501005, 500517, 
    500314, 500952, 500822, 500639, 499516, 500038, 499264, 500929, 499060, 
    499991, 498960, 499231, 498842, 499698, 498733, 498185, 498231, 499160, 
    498595, 498417, 498201, 497991, 497614, 499411, 497592, 497492, 497269, 
    498198, 497409, 497529, 498002, 496332, 497350, 496226, 498458, 496328, 
    496692, 496812, 496751, 497327, 496608, 497087, 496340, 497223, 496045, 
    496328, 496220, 496755, 496483, 496633, 496595, 495526, 495572, 497082, 
    495931, 496165, 496094, 496803, 496139, 495484, 496458, 496169, 495947, 
    496036, 495911, 495834, 496109, 496248, 495924, 496669, 495222, 497388, 
    495256, 495878, 496841, 496445, 496535, 496548, 495692, 496382, 496011, 
    496859, 496112, 496870, 496446, 496864, 497074, 496280, 496732, 496010, 
    497300, 497907, 496321, 497394, 496293, 497919, 497855, 496920, 497672, 
    496987, 498361, 497670, 497575, 497873, 497663, 498233, 498379, 498867, 
    498549, 497836, 498986, 498491, 498678, 498981, 498982, 499188, 499426, 
    499885, 498885, 500914, 498928, 500682, 499423, 500948, 500225, 500270, 
    500601, 501011, 500718, 501208, 501216, 502015, 501573, 502228, 501454, 
    502260, 502740, 501938, 503117, 502844, 503380, 502543, 503543, 503536, 
    503416, 504320, 504360, 504548, 504007, 505733, 504829, 504682, 505592, 
    505553, 505599, 506127, 506303, 506369, 506496, 507108, 507144, 507395, 
    507475, 507855 ;

 true_corr_mean =
  -0.91422406432208, -0.84410960146685, -0.80063819212064, -0.76698005889334, 
    -0.73877502020302, -0.71442223133084, -0.69217397672413, 
    -0.67271718874234, -0.65442533929941, -0.63721243485131, 
    -0.62086169369425, -0.60574841809919, -0.59137253744634, 
    -0.57821354172648, -0.5653489595091, -0.5535613649943, -0.54087094944442, 
    -0.52987118824606, -0.51832709730631, -0.50803831803807, 
    -0.49756484784239, -0.48762812347576, -0.47725847118502, 
    -0.46736213198784, -0.4588815391273, -0.44944707135721, 
    -0.44046070268354, -0.43132672453554, -0.42281362095163, 
    -0.41524400031395, -0.40726473279983, -0.39880731785881, 
    -0.39111719264474, -0.38357000909152, -0.37486955371378, 
    -0.36812993443296, -0.36079132000696, -0.35295365593026, 
    -0.34558021857764, -0.33917040871049, -0.33152629672594, 
    -0.32555170804078, -0.31956582492203, -0.31164604119077, 
    -0.30625254207282, -0.29909569159832, -0.29194388627021, 
    -0.28560778285507, -0.27932679236584, -0.27387716389391, 
    -0.26723065611815, -0.26170147349808, -0.25530808700615, 
    -0.24945464074073, -0.24226389001207, -0.23797376996038, 
    -0.23151547806015, -0.22600359448068, -0.22060978525014, 
    -0.21452629874148, -0.2085085405703, -0.20204647107039, 
    -0.19726903077983, -0.19117292926468, -0.18554804073335, 
    -0.18066063387642, -0.17460029860471, -0.16902019621277, 
    -0.16335579520582, -0.15827183191941, -0.15250098696828, 
    -0.14722250729318, -0.14282052535051, -0.13675862666148, 
    -0.13122010981152, -0.12627055408607, -0.12095221136971, 
    -0.11620059077544, -0.1108632901438, -0.10564929465438, 
    -0.10062377837472, -0.095361403898802, -0.08999809194018, 
    -0.084413529449511, -0.079779707997484, -0.074470007357889, 
    -0.06940465042844, -0.06576614846818, -0.059298422602588, 
    -0.055820403868636, -0.04966853859115, -0.044218064078325, 
    -0.038172438689745, -0.034031712856491, -0.028674237336581, 
    -0.022931936388374, -0.019429565818024, -0.013495761058513, 
    -0.0081913566329826, -0.0052680421500628, 0.0011555086265932, 
    0.0066153805594955, 0.012809315904064, 0.015896665821187, 
    0.02126283574041, 0.026047896920484, 0.031291152703625, 
    0.037012806817124, 0.041642716437319, 0.046912221847253, 
    0.051932958224994, 0.056338244864607, 0.061792718505379, 
    0.067103827976379, 0.072143787772147, 0.077739816805208, 
    0.082839893505012, 0.08757492160699, 0.093714295596221, 
    0.098554384029508, 0.10239864023278, 0.10905836772215, 0.11383615714416, 
    0.11864557746247, 0.12541219604748, 0.13084765984421, 0.13527342587886, 
    0.13945913710316, 0.14565816593223, 0.15169759965083, 0.15618919819038, 
    0.16174913898423, 0.16776857460018, 0.17275370314835, 0.17829757311887, 
    0.18453964638609, 0.1896614046434, 0.195500852599, 0.20197197784348, 
    0.20678574467681, 0.21166835151976, 0.21791287162081, 0.22425666336843, 
    0.23054139955639, 0.2355525837883, 0.24146048002303, 0.24766715897237, 
    0.25345994987784, 0.2605573659572, 0.26516115841829, 0.27227979204318, 
    0.27900224169338, 0.28538330616215, 0.290751991813, 0.29871048505678, 
    0.30451454565107, 0.31076384849976, 0.317491555095, 0.32515562029063, 
    0.33151806143897, 0.338177819845, 0.34623823172978, 0.35265695040672, 
    0.35954398993445, 0.36823697953954, 0.37499560602309, 0.38286992066235, 
    0.39016078972741, 0.39792449272143, 0.40653854096824, 0.41474740128073, 
    0.42306872977236, 0.43127773565842, 0.43991874185273, 0.44827519657868, 
    0.45820558079136, 0.46822066915064, 0.47751414372781, 0.48713988387448, 
    0.49666501391748, 0.50827286062729, 0.51904102334379, 0.5291989169524, 
    0.5411580543238, 0.55309874213919, 0.56549260606744, 0.57833591585293, 
    0.59171667707737, 0.60540368947133, 0.62140576904267, 0.6366896876883, 
    0.65449836299787, 0.6728720498427, 0.69224822123991, 0.71417113642291, 
    0.73851939587299, 0.76669308161827, 0.79999842499369, 0.84368754682866, 
    0.91501750216605,
  -0.95641968254552, -0.90213248852708, -0.86339281356782, -0.83157966981503, 
    -0.80451750467232, -0.78000942000833, -0.75812938206619, 
    -0.73815247232928, -0.71903663508933, -0.70104488569822, 
    -0.68405857832665, -0.66856439757194, -0.65376993434638, 
    -0.63911145555915, -0.62502296005863, -0.61192294968434, 
    -0.59857348984926, -0.58643541134611, -0.574042473681, -0.56274555652524, 
    -0.55183587234437, -0.54078666149598, -0.53011874188502, 
    -0.51935448304138, -0.50960746768947, -0.50030412641051, 
    -0.48948831463901, -0.4808155600442, -0.47125618349479, 
    -0.46237670946911, -0.45327641369364, -0.44407756261734, 
    -0.43599444575156, -0.42711787227281, -0.41909318081087, 
    -0.40991264976859, -0.40332938953121, -0.39450435217786, 
    -0.38652125847884, -0.37966189588118, -0.37112878085899, 
    -0.36328062414909, -0.35557073774414, -0.34849159492327, 
    -0.3410798040156, -0.3340649233422, -0.3267164516, -0.32003572887252, 
    -0.31173870554805, -0.30558365793579, -0.29892766597056, 
    -0.29256494926598, -0.28543671327774, -0.27839206350423, 
    -0.27233091832167, -0.26473517894368, -0.25849489053831, 
    -0.25263240364353, -0.24620899757222, -0.24041543563962, 
    -0.23372753797614, -0.2266487728444, -0.2203460392612, -0.21361975638407, 
    -0.20801519724382, -0.20108217551039, -0.19415441079217, 
    -0.18990466687689, -0.18319996277618, -0.17746942166066, 
    -0.17115354964367, -0.16495253058818, -0.15929557762703, 
    -0.1538485211512, -0.1466338879456, -0.14082223830929, -0.13560962767593, 
    -0.13019512064771, -0.12278441180752, -0.11793710690066, 
    -0.11209519124083, -0.10588890550015, -0.10154307165891, 
    -0.094729575998406, -0.089612521654823, -0.083514963527927, 
    -0.078560149326742, -0.072393640307653, -0.066613411451206, 
    -0.060955235006016, -0.055384834022522, -0.049615029986024, 
    -0.043158759904934, -0.038010652423138, -0.03259331520554, 
    -0.025572776302094, -0.021202088171323, -0.014733264545969, 
    -0.0090593058641659, -0.0028313912409652, 0.00217285446923, 
    0.0073019878384526, 0.011689761702464, 0.018440647787705, 
    0.02375727771307, 0.030483644819787, 0.036459712666433, 
    0.041464932937276, 0.047956939881558, 0.053402123750221, 
    0.059653166744689, 0.064613115999531, 0.069546067791768, 
    0.074748799980465, 0.080697657885074, 0.087025095449924, 
    0.091788048216327, 0.099073597882204, 0.10440321131323, 0.1106132249678, 
    0.1164728610814, 0.12320886399426, 0.12812036791038, 0.13311829218287, 
    0.13949165507955, 0.14601053406596, 0.1524254760966, 0.15886442867667, 
    0.16408777657007, 0.16965234122277, 0.17557551683787, 0.1827384537784, 
    0.18900265449707, 0.1939556664997, 0.19936787980179, 0.2060196133071, 
    0.21169553631673, 0.21899760874322, 0.22454145860269, 0.23124616297703, 
    0.23768458815907, 0.24461868006792, 0.25118416194585, 0.25708791664529, 
    0.26406700385639, 0.27109539818364, 0.27746736494376, 0.28413298004149, 
    0.29100338983333, 0.29747230729931, 0.30482536256005, 0.31295161378063, 
    0.3185572675701, 0.32555387781976, 0.33287099201248, 0.3403723187029, 
    0.34744451863741, 0.35517857960393, 0.36193338740076, 0.36983477409619, 
    0.37834041615366, 0.3849096512336, 0.39314431326819, 0.40091974357716, 
    0.40927270550557, 0.41772699207791, 0.42635624878417, 0.43490024627741, 
    0.44320020322934, 0.45216685156529, 0.46181865623683, 0.47025207248927, 
    0.48067766699341, 0.4895676695836, 0.49946058281455, 0.50941734154092, 
    0.51989209387133, 0.52952212328197, 0.54171064552613, 0.55134314622923, 
    0.56304013357245, 0.57463606662255, 0.58697561355864, 0.59852238761686, 
    0.61107538220144, 0.62502385341136, 0.63864696677968, 0.6525949690723, 
    0.66838068457924, 0.68371423438429, 0.70050665680128, 0.71820847011246, 
    0.73710672328271, 0.75765349870171, 0.78027402809347, 0.80416617943094, 
    0.83149095557645, 0.86311477651041, 0.90183737446643, 0.95619966151913,
  -0.97307639069551, -0.9315440118424, -0.89815046373525, -0.86980411525962, 
    -0.84455517413096, -0.82113118103997, -0.8001901888558, 
    -0.78029414578644, -0.76150489475609, -0.74405980638381, 
    -0.72722102272073, -0.71107028377493, -0.69590479933687, 
    -0.68102788558212, -0.66675703435158, -0.65355129117552, 
    -0.64036619730328, -0.62698343853487, -0.61512544193136, 
    -0.60312107771159, -0.59103613225559, -0.58004509855493, 
    -0.56915342314904, -0.55784527496809, -0.54718029393368, 
    -0.53692318732542, -0.52684658365455, -0.51714922747134, 
    -0.50664979682958, -0.49750649144299, -0.48760533524565, 
    -0.47846049053922, -0.46890241593541, -0.46023930134435, 
    -0.45131353832578, -0.44278812675827, -0.43310711970053, 
    -0.42528714267802, -0.41720164608834, -0.40873415618155, 
    -0.4003435469265, -0.39207377188027, -0.38450155788632, 
    -0.37640495679383, -0.3690236237688, -0.3606518653809, -0.35287466791548, 
    -0.34596265758135, -0.33771517098913, -0.33036902168253, 
    -0.32322410346499, -0.31609127529756, -0.3083570916597, 
    -0.30052191133121, -0.29474047594691, -0.28720765658298, 
    -0.27984099069703, -0.27188502257438, -0.26618299271882, 
    -0.25843313735899, -0.25205241186197, -0.24416070539279, 
    -0.23792007612272, -0.23229036295218, -0.22575701770608, 
    -0.21872840811187, -0.21128934588886, -0.20581366742085, 
    -0.19729897607929, -0.19182646038084, -0.18494271904479, 
    -0.17921777671896, -0.17256348438148, -0.16564687054199, 
    -0.15963935154144, -0.15283163403764, -0.14700763826294, 
    -0.13992200400925, -0.1343583320511, -0.12732605298355, -0.1224059067321, 
    -0.11523925122195, -0.1086414662357, -0.10311881904642, 
    -0.096994948114717, -0.090023373718709, -0.084387594228376, 
    -0.078088580974186, -0.071916264658538, -0.065045381492781, 
    -0.059126041474212, -0.053378883003383, -0.04672952961958, 
    -0.040750276348133, -0.035182285270467, -0.028521227104992, 
    -0.022579753509271, -0.017080276385069, -0.010146538751492, 
    -0.0032755107870317, 0.0021140214808052, 0.0086097517927013, 
    0.014744460345342, 0.021048830289636, 0.026212076681186, 
    0.032650573018009, 0.038420100860528, 0.045260027629368, 
    0.051936589758108, 0.057838820757187, 0.063087820596362, 
    0.070465695016431, 0.075605543350087, 0.082336576260628, 
    0.087862477402271, 0.094321905212631, 0.10125254439357, 0.10758409161152, 
    0.11358049369815, 0.12063416794099, 0.12604378200268, 0.13223266964112, 
    0.13898152884328, 0.14460118329046, 0.15181534047344, 0.15840171333421, 
    0.16460082970012, 0.17065136238654, 0.17684163279183, 0.18309110823908, 
    0.19048465657191, 0.19739563951153, 0.20350054516061, 0.21050238491325, 
    0.21707155785275, 0.22326071422324, 0.23049605258314, 0.23730662028309, 
    0.24410646645246, 0.250179758568, 0.2576296821045, 0.2642025365361, 
    0.27175106336417, 0.27805522527579, 0.28604257681474, 0.29275014013621, 
    0.30043980650294, 0.30754353057931, 0.31475266641356, 0.32244087754742, 
    0.32957001223411, 0.33772380667286, 0.34434134201191, 0.35193512400763, 
    0.35942493575578, 0.36834341147936, 0.37494097986674, 0.3836282174317, 
    0.39118140559156, 0.39934645529189, 0.40767836486987, 0.4152187123123, 
    0.42435714131746, 0.43258836878782, 0.44189719585642, 0.45065781168824, 
    0.45974110803122, 0.46827179003587, 0.47819383188703, 0.48685048221112, 
    0.49611984565897, 0.50634875209864, 0.51634149593265, 0.52612639790543, 
    0.53595657542097, 0.54621605279673, 0.55696016813613, 0.56834004121549, 
    0.57939885327544, 0.59096704198912, 0.60302983887139, 0.61464066235351, 
    0.6274813623486, 0.64047231732954, 0.65354321930849, 0.66689889341169, 
    0.68074354488773, 0.6956145636294, 0.71082860999534, 0.72688818306422, 
    0.74340235017717, 0.76115982556054, 0.77973651932612, 0.79977853673633, 
    0.82098567326844, 0.84412066198856, 0.86950937259416, 0.89834361950787, 
    0.93135983980689, 0.97306033742775,
  -0.98059113239332, -0.94723468857226, -0.91850295778626, -0.89292417063092, 
    -0.86961238119388, -0.84819591632845, -0.82817072972195, 
    -0.80888481316382, -0.79098641929162, -0.77372887917093, 
    -0.75711265114012, -0.74172631579557, -0.72672095376987, 
    -0.71204715173673, -0.69773014770622, -0.68389741121651, 
    -0.67045760347567, -0.65776695470944, -0.6455224239162, -0.6327943243208, 
    -0.62123376857675, -0.60935530577737, -0.59832929359986, 
    -0.58691026284981, -0.57592685188602, -0.56523762068282, 
    -0.55487088902376, -0.54447612711052, -0.53420563483318, 
    -0.52446169361992, -0.51462982340766, -0.50461223668665, 
    -0.49508516207994, -0.48546191109992, -0.47664979344233, 
    -0.46761465277847, -0.45829875567102, -0.45023531128347, 
    -0.44061136060947, -0.43212423272329, -0.42344325383076, 
    -0.41476781857783, -0.40637797914418, -0.39777308380896, 
    -0.38914699305441, -0.38181888732596, -0.37363935320785, 
    -0.36554631885112, -0.35810686109857, -0.35060158750604, 
    -0.34222809653271, -0.33477434218603, -0.32639243581294, 
    -0.31892498368152, -0.31161898690076, -0.30377195912537, 
    -0.29649756265093, -0.28914660337765, -0.28173294363123, 
    -0.27408121714927, -0.26776162908709, -0.26001696585194, 
    -0.25373485996457, -0.24487487321119, -0.23919643088725, 
    -0.23142582194735, -0.22369319679368, -0.21752663997695, 
    -0.21079497385377, -0.20311310212722, -0.19658353215066, 
    -0.18880932261727, -0.18267074746071, -0.1755570565089, 
    -0.16973008322439, -0.16246302879441, -0.15569729945427, 
    -0.14909810668442, -0.14291579821208, -0.13603384937889, 
    -0.12892001846627, -0.12212228849081, -0.11549120954789, 
    -0.10801043666649, -0.10234330974851, -0.095800895273832, 
    -0.089252216087431, -0.081951001943509, -0.075906927325395, 
    -0.069004304686659, -0.062754642214986, -0.056156034374322, 
    -0.049618077545133, -0.043513428794832, -0.036044779748387, 
    -0.030563824841987, -0.023297142093166, -0.017828801720461, 
    -0.010792265441573, -0.0045105641263034, 0.0022339166974139, 
    0.0090043000533902, 0.016097417105558, 0.021345506852452, 
    0.028847629156401, 0.034367678242738, 0.042529953037325, 
    0.048064360576935, 0.05369498335482, 0.061710956528507, 
    0.067623201187854, 0.075403524820758, 0.080489340618992, 
    0.08793688809438, 0.094840613998025, 0.10069772200169, 0.10780160045377, 
    0.11392140883889, 0.12075342822906, 0.12790748270398, 0.13430876011311, 
    0.14014943677746, 0.14743463263292, 0.15401659579795, 0.16129113493249, 
    0.16714483225402, 0.17449289528776, 0.1816495116878, 0.18819746163199, 
    0.19574264906041, 0.20244575853496, 0.20848975948753, 0.21597070971149, 
    0.22366650443111, 0.23046630650948, 0.23674936289909, 0.24361011355456, 
    0.25054332643566, 0.25763382477016, 0.26530257663348, 0.27330650138753, 
    0.28078541150562, 0.28810639474325, 0.29528133341153, 0.30199497117329, 
    0.31048983109975, 0.31733810623573, 0.32535744600359, 0.33301836081866, 
    0.3406399977586, 0.3488048204257, 0.35776605184868, 0.36389449558332, 
    0.3730415106518, 0.38063159796547, 0.38882197533816, 0.39741485425693, 
    0.40551722278381, 0.41351150329907, 0.42276058608016, 0.43068421965796, 
    0.44005775970863, 0.44907426879125, 0.45705363816698, 0.46677282896675, 
    0.47589253600098, 0.48505373055408, 0.4944752838117, 0.50376697685014, 
    0.51388347529003, 0.52343426269299, 0.53361203675042, 0.5443082571551, 
    0.55423971429891, 0.56464053729904, 0.57580539486812, 0.58643236863315, 
    0.5971960609108, 0.6090414575871, 0.62115363287734, 0.63249697110969, 
    0.64511229882535, 0.65755495434443, 0.67089464628405, 0.68409315951926, 
    0.69728577344714, 0.71177563791888, 0.72675009052015, 0.74166192222384, 
    0.7572313470823, 0.7734393576335, 0.79097124722114, 0.808686400587, 
    0.82775937557782, 0.84810782191398, 0.86982409171684, 0.89297662423788, 
    0.91846967106963, 0.94706334628638, 0.98059577211378,
  -0.98453050618317, -0.95638323169049, -0.93109234066881, -0.90785601148585, 
    -0.88645402671436, -0.86637324950131, -0.8475814078245, 
    -0.82945569074979, -0.81192181628762, -0.79538594315209, 
    -0.77923709899345, -0.76396092676975, -0.7484357991487, 
    -0.73415379256996, -0.72050887106444, -0.70677005852504, 
    -0.69329062222143, -0.68038319485063, -0.66755104491097, 
    -0.65589476601296, -0.64380780540071, -0.63185025018048, 
    -0.62015076088275, -0.60922102049782, -0.59831565190844, 
    -0.58706305556871, -0.57546525135468, -0.56596329109146, 
    -0.55515677394516, -0.54456489363835, -0.53506625253723, 
    -0.5243723799786, -0.51525949571617, -0.50552738618262, 
    -0.49613946839686, -0.48686040509558, -0.47764317265312, 
    -0.4681675811243, -0.45854489347261, -0.44995942617536, 
    -0.44036586847507, -0.43214905177966, -0.42492978422482, 
    -0.41593998997063, -0.40641954612616, -0.39790368935406, 
    -0.39024600997675, -0.38221077011633, -0.37353157672184, 
    -0.36613228807195, -0.35768034365596, -0.34901928070251, 
    -0.34087347224075, -0.33303522031993, -0.32617739995972, 
    -0.31815985338484, -0.31041607907298, -0.30218107600689, 
    -0.29377615408174, -0.28718650612497, -0.27962916201865, 
    -0.27192130724483, -0.26429178766757, -0.25660992243032, 
    -0.24874714433289, -0.24149695897593, -0.23419308978068, 
    -0.22751613392986, -0.21989376224293, -0.21336362645559, 
    -0.20655755899067, -0.19861378343604, -0.19115135293511, 
    -0.18467558196155, -0.17750350170794, -0.17025356704977, 
    -0.16342546878724, -0.15649675266523, -0.14869060331676, 
    -0.14227648665168, -0.1347480137304, -0.12776683836531, 
    -0.12119850778602, -0.11401551818533, -0.10662520506537, 
    -0.099809499504984, -0.092941027163904, -0.085728609394218, 
    -0.079313908175688, -0.072140623249209, -0.065510506617258, 
    -0.058653593155606, -0.05197614235913, -0.044626294081047, 
    -0.037960500805048, -0.031020655703719, -0.024743016939464, 
    -0.018372087457179, -0.011198240263612, -0.0047551654108496, 
    0.0019078369712503, 0.009325495623367, 0.016209434246992, 
    0.022957025605432, 0.030451514868021, 0.036488027402453, 
    0.042762566007428, 0.050777544020723, 0.056400702023452, 
    0.06404237194348, 0.070543573854786, 0.07777322169898, 0.08444063500031, 
    0.091879119417744, 0.098445234035757, 0.10603177133903, 0.11291830683745, 
    0.11955415369571, 0.12632353408638, 0.13374338353884, 0.14011427714159, 
    0.1472135171287, 0.15556924715054, 0.16161527429781, 0.1681632362679, 
    0.17537916054092, 0.18239353452059, 0.18974056113759, 0.1967503272486, 
    0.20492719722282, 0.21141541566631, 0.21881182232828, 0.22598808718441, 
    0.23398372123349, 0.24067650593468, 0.24795001031139, 0.25548910457922, 
    0.26381459702194, 0.27046913402915, 0.27835825639136, 0.28457542040843, 
    0.29358125186553, 0.30085942268752, 0.30845178909034, 0.31680647337043, 
    0.32468308988794, 0.3320506513404, 0.34018813340883, 0.34783407967345, 
    0.35641514288117, 0.36383535490388, 0.37240949014267, 0.38105240951058, 
    0.3896383300513, 0.39800403991689, 0.40592248462862, 0.4144667600395, 
    0.42288692711128, 0.4320279663353, 0.44081333662991, 0.449457185052, 
    0.45946120043391, 0.46836557605228, 0.47691027442073, 0.48601771918043, 
    0.49616575717742, 0.5046323051553, 0.514673547583, 0.52521915528185, 
    0.53503625669775, 0.54576732101957, 0.55456677870114, 0.5657495903559, 
    0.576826926609, 0.58735234357191, 0.59802985249729, 0.60856350083766, 
    0.62052220217113, 0.63162556794126, 0.64387156445236, 0.65623994184418, 
    0.66881508123818, 0.6809449041665, 0.69372491476858, 0.7071245990065, 
    0.72101128177699, 0.73502809064036, 0.74919160794201, 0.76394423782525, 
    0.77961056159563, 0.79535452431426, 0.81221736942292, 0.82951945707565, 
    0.84722191255327, 0.86651536403004, 0.88667798495835, 0.90830488535106, 
    0.93126884025385, 0.95636643531402, 0.98458600829509,
  -0.98692108394874, -0.96216541392244, -0.93969203641566, -0.91832515706478, 
    -0.89827488702818, -0.87945882234701, -0.86138369600949, 
    -0.84399239819833, -0.82747427725838, -0.81134541761832, 
    -0.79549129578568, -0.7805186422965, -0.76553984102606, 
    -0.75195471493996, -0.73781689288248, -0.72413242671552, 
    -0.71150166904376, -0.69819705709669, -0.68529949861269, 
    -0.67288756701931, -0.66112016799281, -0.64938834629148, 
    -0.63837421390333, -0.62606130508473, -0.61549140083281, 
    -0.60469443529874, -0.5928780503571, -0.58252693184296, 
    -0.57177434131444, -0.56204175681709, -0.55164862673118, 
    -0.54183633723547, -0.53210992530264, -0.52219046912736, 
    -0.5130063593774, -0.50283117894808, -0.49270179182967, 
    -0.48367775491096, -0.47506737657277, -0.4662186089009, 
    -0.45734692412882, -0.4480799913128, -0.43857642851235, 
    -0.42928332916759, -0.42113861639979, -0.41286900993756, 
    -0.40354898897396, -0.39462103792893, -0.38619602648229, 
    -0.37839826161776, -0.3691923582123, -0.36188596438372, -0.3536442694547, 
    -0.34639301779252, -0.33661138377697, -0.32918536564525, 
    -0.32104043083711, -0.31346638559211, -0.30478229038043, 
    -0.29700692466347, -0.28923110978902, -0.28202170502266, 
    -0.27342150588526, -0.26598618257524, -0.25832607238134, 
    -0.25066200611938, -0.24432622226012, -0.23507353286981, 
    -0.22769139859159, -0.21982700349035, -0.21317680452133, 
    -0.20559447719603, -0.19808290868751, -0.190972013459, -0.18327865261111, 
    -0.17627315190451, -0.16817560524816, -0.161717962225, -0.15483734247665, 
    -0.14690513939189, -0.1402696276837, -0.13321450708159, 
    -0.12546280784869, -0.11746952042558, -0.11035045511053, 
    -0.10308537597911, -0.096347742405082, -0.089515107049557, 
    -0.082663534206482, -0.075002080748604, -0.06806756980612, 
    -0.060384926320598, -0.054034545334954, -0.047199040404411, 
    -0.03944375743121, -0.033196421305925, -0.026569542792041, 
    -0.018095344729595, -0.011007113837686, -0.0050633694643769, 
    0.0019632149297667, 0.0098811542400421, 0.016733562002314, 
    0.023504047426956, 0.031276624480566, 0.038570223044776, 
    0.045398029230586, 0.052708588725383, 0.059843577973917, 
    0.066940262104605, 0.073220737889992, 0.080521023158044, 
    0.087925237706917, 0.095362195661132, 0.10209790596058, 0.11021212607394, 
    0.11627807108129, 0.12414552974295, 0.13112175306859, 0.13915468960149, 
    0.14572435551335, 0.15336054141217, 0.16091229244137, 0.16799627703388, 
    0.17556975546782, 0.18262076044035, 0.18998719412891, 0.19767210542417, 
    0.20375417882061, 0.21205251239681, 0.22019391956267, 0.22705257741921, 
    0.23503651423081, 0.24285802718598, 0.25084058402287, 0.25808863156146, 
    0.26465574477045, 0.27262528045803, 0.28084607133767, 0.28857920589495, 
    0.29485764277368, 0.30383275236414, 0.31167051708781, 0.31943338970183, 
    0.3279054570631, 0.3366012302031, 0.34478945592093, 0.35239541841411, 
    0.36046506032406, 0.36910980415166, 0.3774655017327, 0.38606411154956, 
    0.39402203949903, 0.40328346350267, 0.41117210838464, 0.42048676128139, 
    0.42934510857998, 0.43811630479396, 0.44659130315508, 0.45512658678669, 
    0.4650277317443, 0.47375512323881, 0.48361109824207, 0.49360889056605, 
    0.50300642935449, 0.51236772654521, 0.52208759566858, 0.53257861990053, 
    0.54161128589946, 0.55163036931126, 0.56235043991657, 0.57259433645547, 
    0.58361451846661, 0.5937597515382, 0.60467569423851, 0.61551810496288, 
    0.62687035083191, 0.63804413548201, 0.64980842461016, 0.661594167002, 
    0.67423699913736, 0.68578500037901, 0.69925822402327, 0.71195775191995, 
    0.72491493339854, 0.73846153047604, 0.75227484778836, 0.76673063791039, 
    0.78106878902846, 0.79560669579219, 0.81158491368626, 0.82744249703834, 
    0.84410224450396, 0.86157285756156, 0.87954841309534, 0.89831049764212, 
    0.91858027142574, 0.93967631311412, 0.96239776234364, 0.9869194101149,
  -0.98944428453551, -0.96905741282638, -0.94965647449589, -0.93104975233375, 
    -0.91348385524595, -0.8961773858258, -0.87991674757833, 
    -0.86361733736398, -0.84827185229546, -0.8329145720352, 
    -0.81824624370735, -0.80383124050345, -0.79012226846032, 
    -0.77594287104227, -0.76309052770519, -0.74952153693874, 
    -0.7369050415259, -0.72427569176878, -0.71110059742837, -0.6996994761584, 
    -0.68722396644304, -0.67566003903724, -0.6639035713301, 
    -0.65261022118213, -0.64117630423096, -0.62956510554903, 
    -0.61941301162246, -0.60846741362401, -0.59728276662017, 
    -0.5869868853131, -0.57666933971427, -0.56634897480369, 
    -0.55691611141631, -0.5463415867203, -0.5359937118691, -0.52714161374844, 
    -0.51657138578949, -0.50811952740327, -0.49773725616522, 
    -0.48804822829469, -0.47897961728374, -0.46986264961796, 
    -0.46106956966285, -0.45109868788691, -0.44205281993121, 
    -0.4331446436931, -0.4240918603609, -0.4155189938124, -0.40665995440703, 
    -0.39826548759959, -0.38949962740339, -0.38086490711914, 
    -0.37170356301828, -0.36298338557212, -0.35557827748064, 
    -0.34701455865543, -0.33777577935112, -0.33024062992604, 
    -0.32163607236416, -0.31321158040649, -0.30501141763928, 
    -0.29646787047798, -0.2884452595267, -0.28014977998282, 
    -0.27102558425906, -0.26439375990474, -0.256756734758, -0.24829727031282, 
    -0.2413039362399, -0.23358635520534, -0.22514112800526, 
    -0.21742218686196, -0.20923051478888, -0.20103920131232, 
    -0.19341177912978, -0.18537267955758, -0.17802809701282, 
    -0.17080490193051, -0.16266668913291, -0.15526907718123, 
    -0.14823442701727, -0.14031061183571, -0.13279051498602, 
    -0.12551972789599, -0.11766742301028, -0.10976351472573, 
    -0.1009129708009, -0.094602189535633, -0.086660882728838, 
    -0.079508464633527, -0.072009062205962, -0.065202533771344, 
    -0.056500355481097, -0.049237618360911, -0.042501132886451, 
    -0.03465578662393, -0.026651686828482, -0.019246289984669, 
    -0.012387959087937, -0.0051732234210468, 0.0029374768781016, 
    0.01016517031883, 0.01788185828032, 0.025151999564964, 0.033263899017098, 
    0.042296961593155, 0.049171814361699, 0.055940114971325, 
    0.063206199922759, 0.071079228406567, 0.078091161327251, 
    0.085850383700763, 0.092972906485695, 0.10047737874409, 0.10850956919429, 
    0.11619844952288, 0.12335959495891, 0.13200214950437, 0.13954113285563, 
    0.14687983431723, 0.15449616635082, 0.16220615679311, 0.17019069063563, 
    0.17722795180418, 0.18497859130646, 0.19287208508902, 0.20104718400481, 
    0.20844160831568, 0.21689374137253, 0.22482142045668, 0.23231439475024, 
    0.24044044858538, 0.24774750878926, 0.25561698803929, 0.26448157094122, 
    0.27247653612006, 0.28084253390972, 0.28826481550349, 0.29677490670079, 
    0.30523337826229, 0.31253634240435, 0.32104173635238, 0.32904778347319, 
    0.33752921720534, 0.34558610922747, 0.35538105695234, 0.36317555359664, 
    0.3717305559779, 0.38048213708446, 0.38934852777548, 0.39753840142599, 
    0.40661385048972, 0.41490836173883, 0.42362976239278, 0.433260325515, 
    0.44253742960382, 0.45079960588311, 0.46015046748417, 0.46969748808484, 
    0.47905693754447, 0.48801743058009, 0.49729273399122, 0.50714100757849, 
    0.51780380259748, 0.5275486174629, 0.53647620628692, 0.54724798927621, 
    0.55651973358721, 0.56716932434071, 0.57829001169476, 0.58724637138951, 
    0.5976712899079, 0.60860379240499, 0.61920696723353, 0.63101838360293, 
    0.64184284666969, 0.65304349796741, 0.6648449875331, 0.67614430948483, 
    0.68811711975401, 0.69970119485919, 0.71239467986254, 0.72451198784618, 
    0.737098364346, 0.7496469592149, 0.76304901235758, 0.77648472240222, 
    0.7903529312941, 0.80392156762039, 0.81885033043815, 0.83351042388431, 
    0.84809282344455, 0.86365562125779, 0.8798488763052, 0.89631407134844, 
    0.91329566197101, 0.93121383549418, 0.94978119694713, 0.96905200326114, 
    0.98942106247002,
  -0.99078427609444, -0.97279372592768, -0.95539839133846, -0.93863065452524, 
    -0.92236523141767, -0.90643337442274, -0.89103178765765, 
    -0.87584798454425, -0.86098412989347, -0.84690771776916, 
    -0.83270168380867, -0.81878225854403, -0.80531005403958, 
    -0.79226006558776, -0.77902305964738, -0.76621385317601, 
    -0.75371797274083, -0.74133181245985, -0.72910926879469, 
    -0.71689054237457, -0.70494154622427, -0.69351948113865, 
    -0.68205128279038, -0.67045903596825, -0.65978170253252, 
    -0.64826753595881, -0.63719830178707, -0.62648209477228, 
    -0.61581825331739, -0.60509981037474, -0.59484585492841, 
    -0.58427094248776, -0.57395410621824, -0.56389309766207, 
    -0.55377600987709, -0.54432131333228, -0.53367651204764, 
    -0.52410100962109, -0.51420840926124, -0.50498449153598, 
    -0.49547990348364, -0.48611921140813, -0.47643943678471, 
    -0.46730109068461, -0.45795827926553, -0.44848519020715, 
    -0.43911260468997, -0.43021146334044, -0.42085607950693, 
    -0.41217817789501, -0.4034688049478, -0.39480482639627, 
    -0.38570158132042, -0.37697459686127, -0.36857243715395, 
    -0.35926394040391, -0.35046837870966, -0.34201894011424, 
    -0.33411234385306, -0.32523950546747, -0.31658283327175, 
    -0.3087220912504, -0.29979906653717, -0.29153818045001, 
    -0.28316480483961, -0.27454114540661, -0.26704691164334, 
    -0.25816113134501, -0.24997266278457, -0.24177527027088, 
    -0.2338603069807, -0.22538852766759, -0.21791540638611, 
    -0.20992123066651, -0.20171127727043, -0.1935569685381, 
    -0.18486969818418, -0.17792830743159, -0.16980097302556, 
    -0.16166013604224, -0.15314191465816, -0.14556576065694, 
    -0.13775384605434, -0.12927254345971, -0.12185827942344, 
    -0.11388617898633, -0.10576614735137, -0.097939297789106, 
    -0.090394462599956, -0.082457867943828, -0.074295645482091, 
    -0.066904188634558, -0.059397302255641, -0.050955687423798, 
    -0.04273021630066, -0.035705300610918, -0.027157366765487, 
    -0.01987673531571, -0.011891673005048, -0.0041686182233261, 
    0.0036355100924805, 0.011265913368061, 0.019275813245188, 
    0.026773679607073, 0.034370904278513, 0.042537583172028, 
    0.050111645402315, 0.05859829249087, 0.065454372694967, 
    0.073484796947342, 0.082111670195039, 0.089596837706907, 
    0.097313069157496, 0.1053594372186, 0.11351629036356, 0.12103294314236, 
    0.1292290633716, 0.13695199019644, 0.14471180350179, 0.1532099012082, 
    0.16074978940604, 0.16882633408913, 0.176413823395, 0.18498942627228, 
    0.19316401423854, 0.2008885320532, 0.20925957789834, 0.21676582723791, 
    0.22535362181849, 0.23308698750691, 0.24115988475565, 0.25017381897536, 
    0.25809992544809, 0.26643859147848, 0.27402073871208, 0.28276630820751, 
    0.29141906287627, 0.2995219847401, 0.30807437628252, 0.31707925768995, 
    0.32503064029166, 0.3341402825222, 0.34238847853576, 0.35025855224595, 
    0.35972190599236, 0.36799097928715, 0.37645743507284, 0.38572079185073, 
    0.39489561661207, 0.40344083945407, 0.41232402844188, 0.42129543938378, 
    0.43058633738285, 0.4393132552794, 0.44838520587402, 0.45752176036124, 
    0.46666212993597, 0.47669355393682, 0.48563854314742, 0.49563280389442, 
    0.50512319609582, 0.51484197669237, 0.52422627778447, 0.53414761934511, 
    0.5438978035781, 0.5538617981674, 0.56438354321085, 0.57460758425294, 
    0.58501047141142, 0.59519224756013, 0.6058988089944, 0.61627554773038, 
    0.62726120279485, 0.6375471795049, 0.64866788812769, 0.6601509771698, 
    0.67137904155402, 0.68230933467884, 0.69379737821632, 0.70602507047194, 
    0.71732626450005, 0.72947207171199, 0.74162014587829, 0.75399279304297, 
    0.7669342197676, 0.77933168986692, 0.79267338353592, 0.80595297351295, 
    0.8191813339688, 0.83294119146496, 0.84710352097737, 0.86141174623735, 
    0.87601772304086, 0.89112527103546, 0.90643797993237, 0.92231177070097, 
    0.93861429020346, 0.95536902237491, 0.97279216329416, 0.99077849243671,
  -0.9912591465225, -0.97412719262498, -0.95740343183285, -0.94122073296115, 
    -0.92536272170492, -0.91012519547523, -0.89512516031168, 
    -0.8804838788947, -0.8661848683879, -0.85182267321048, -0.83793159383654, 
    -0.82453646577958, -0.81128535687273, -0.79836885987464, 
    -0.78545278725816, -0.77287923969751, -0.76004700375526, 
    -0.74811725073784, -0.73630155892393, -0.72433679299616, 
    -0.71200423953791, -0.70004742857302, -0.68863813482891, 
    -0.67745247258783, -0.6662718549536, -0.65499581273658, 
    -0.64454348213259, -0.63328135499087, -0.62316903389406, 
    -0.61225695822159, -0.60192078212506, -0.59133880949131, 
    -0.58080893138278, -0.57169668133496, -0.56131193916283, 
    -0.55061297712233, -0.54123577578596, -0.53110609188253, 
    -0.52087980270448, -0.51170765814542, -0.50166846679894, 
    -0.49234883861105, -0.48332285690905, -0.47323372990856, 
    -0.46395472848297, -0.45471074998466, -0.44573326300998, 
    -0.43630223735811, -0.42656761699304, -0.41758926152281, 
    -0.40984624475637, -0.40075856986294, -0.39171745273345, 
    -0.38286095806409, -0.37353384114654, -0.36551580160132, 
    -0.35544055740499, -0.34746632149106, -0.33847988169902, 
    -0.33033073022157, -0.32114926427886, -0.3128053184031, 
    -0.30470853391832, -0.29615770499563, -0.28698600604425, 
    -0.27922877591304, -0.27068287836241, -0.26194630944123, 
    -0.25348650106996, -0.24491340328371, -0.23743419132415, 
    -0.22932900728373, -0.22162183719241, -0.21274909940909, 
    -0.20486272976506, -0.19631051375622, -0.18906752547829, 
    -0.18014549898619, -0.17216446029469, -0.16356623353942, 
    -0.15603705613458, -0.14736742335476, -0.14005432142734, 
    -0.13149534104213, -0.12388632257661, -0.11582680967677, 
    -0.10857331107568, -0.099912678475366, -0.09202954478145, 
    -0.083567571452957, -0.075581947319195, -0.067890817994595, 
    -0.060652637813092, -0.052047158148053, -0.043813755102665, 
    -0.035906381474198, -0.027751713383925, -0.02018095325136, 
    -0.012032029402854, -0.0047661957623276, 0.0037831005296831, 
    0.011956967207018, 0.019637818593956, 0.027219327720406, 
    0.03549652314784, 0.044393091058636, 0.052201792383266, 
    0.059209981609721, 0.06682210166798, 0.074724290718507, 
    0.083089859799063, 0.09140890596322, 0.09887201714518, 0.10690958631324, 
    0.11531075936736, 0.12371904064753, 0.13199589777642, 0.13972709605369, 
    0.14683829767692, 0.15578536117627, 0.16425017481191, 0.17102098478699, 
    0.17977797394585, 0.1877550663755, 0.19562915185794, 0.20402687832613, 
    0.21197491627569, 0.22006814971085, 0.22857326458074, 0.23726320843415, 
    0.24555619107588, 0.25414292375935, 0.26218735434262, 0.27064206676247, 
    0.27927473203522, 0.28739423346111, 0.29592107312211, 0.30358463620508, 
    0.31245499771843, 0.32163441291779, 0.33102800903579, 0.33806799292372, 
    0.3463660236595, 0.35565039085128, 0.36528276875762, 0.37352236255584, 
    0.38250648421476, 0.3914943541704, 0.40012332591946, 0.40878795647342, 
    0.41806629262298, 0.42661008098362, 0.43576187159818, 0.44601144523359, 
    0.45451795254206, 0.46363326796277, 0.47397513099305, 0.48305222604797, 
    0.49253632323355, 0.5019412985523, 0.51229318108257, 0.52186726787725, 
    0.53181225776401, 0.54143184518522, 0.55110038463374, 0.56033240985875, 
    0.57127595405647, 0.58157126093847, 0.5922275619232, 0.60307606875143, 
    0.61271455757289, 0.62281385753537, 0.63365586621479, 0.64498905284624, 
    0.6557728695391, 0.66693852453419, 0.67859645268565, 0.6890674016202, 
    0.70113103704736, 0.71253189735828, 0.72474354085666, 0.7365458212924, 
    0.74843729158662, 0.76045293947891, 0.77330917857683, 0.78571463316836, 
    0.7988208061423, 0.81160517987234, 0.82479786589316, 0.83851769814589, 
    0.85230410519789, 0.86618439211822, 0.88057381549545, 0.89513381462175, 
    0.91008156007037, 0.92545901501396, 0.94113234255802, 0.95732583526316, 
    0.9740734487135, 0.99123758442883,
  -0.99160957570338, -0.97512529565252, -0.95910347532319, -0.94343032357109, 
    -0.92808108829148, -0.91314492767405, -0.89857635517875, 
    -0.88407013671627, -0.87018898621772, -0.8562440360856, 
    -0.84281441779971, -0.82935083661902, -0.81636610957267, 
    -0.80341213668158, -0.79079206532468, -0.77791651067579, 
    -0.76601269424277, -0.75352032147627, -0.7415202058738, 
    -0.72982273050393, -0.71817249564982, -0.70657835402934, 
    -0.6952330164985, -0.6841058225534, -0.67277177066333, -0.66178183510775, 
    -0.65064081960689, -0.63953728722048, -0.62922080657225, 
    -0.6186358749727, -0.60790836060592, -0.59745458240881, 
    -0.58723578773206, -0.57726271777078, -0.56697048469893, 
    -0.55694627340336, -0.54677998964069, -0.53693823302086, 
    -0.5268608858244, -0.51749931357071, -0.50773264445268, -0.4977682314245, 
    -0.48872425994419, -0.47924790282974, -0.46939138284409, 
    -0.46007424090754, -0.45107284304981, -0.4416049075594, 
    -0.43231873214281, -0.42360145014498, -0.41457389897551, 
    -0.40520442143578, -0.39595285709698, -0.38721989237367, 
    -0.37851192348372, -0.36968459506109, -0.36071929994238, 
    -0.35201509603963, -0.34320117720584, -0.33438757627604, 
    -0.32558461109039, -0.3170903075113, -0.30862738440282, 
    -0.30006092176138, -0.29153782237469, -0.28295395566453, 
    -0.27425048362083, -0.26576879161165, -0.25790684401996, 
    -0.24921329437226, -0.24021928487076, -0.23214789844787, 
    -0.22371314851507, -0.21571845309599, -0.2069362422313, 
    -0.19901294164206, -0.19128523940111, -0.18214488889227, 
    -0.17436922092276, -0.16619670992169, -0.1579560633019, 
    -0.14992116220727, -0.14164700673855, -0.13323926330997, 
    -0.12578894462415, -0.11678293136011, -0.1091505064434, 
    -0.10047441046618, -0.093600046930991, -0.08488006436473, 
    -0.076771254716447, -0.068298720982529, -0.060776628528868, 
    -0.052636455094997, -0.04425315457265, -0.037206936112209, 
    -0.028316778766748, -0.019939586771376, -0.012165416326781, 
    -0.0045474201436798, 0.0034994534582872, 0.01151421731344, 
    0.019933616540558, 0.027651160952583, 0.03593706390447, 
    0.044088381763441, 0.051772170434988, 0.060687739939874, 
    0.068791698890493, 0.076019544062937, 0.08446730915383, 
    0.092240197710798, 0.10092145942969, 0.10821518462609, 0.11666935297964, 
    0.12453873660828, 0.13335705814688, 0.14110672870321, 0.14886931587099, 
    0.15784091084833, 0.16559889876196, 0.17410662842225, 0.18226054071254, 
    0.19074553882667, 0.19908535213852, 0.20699984490416, 0.21553517748767, 
    0.22353715236433, 0.2322528019968, 0.24028369958981, 0.24853638395402, 
    0.25738403415685, 0.26569021454479, 0.27397837056005, 0.28273470508392, 
    0.29155957497793, 0.29943278535418, 0.30799452882231, 0.31704271791597, 
    0.32604879891905, 0.33428083732205, 0.34252992365202, 0.35187600599397, 
    0.36048745117736, 0.36976893320887, 0.37848127183183, 0.38731543768118, 
    0.39633106719777, 0.40565817662535, 0.41398610045859, 0.42364369141157, 
    0.43247961559884, 0.44193982257685, 0.45119234798726, 0.46061300875436, 
    0.46998835294444, 0.47951629102618, 0.48893333327275, 0.49874921116396, 
    0.50772890208552, 0.51801789446265, 0.52719775568844, 0.5369729156915, 
    0.54722445788565, 0.55696655556106, 0.56739941523527, 0.57745053210788, 
    0.58748141425718, 0.59779452076921, 0.60850266027022, 0.61922285138432, 
    0.62977153359237, 0.64035171231219, 0.65101535785335, 0.66223378386295, 
    0.673104531025, 0.68427932280472, 0.69571943056445, 0.70707447957934, 
    0.71854648870762, 0.73052149300883, 0.74216475207589, 0.75399137488658, 
    0.76640833942127, 0.77870196944113, 0.79091585591312, 0.80386057758558, 
    0.81664961872544, 0.82970679581869, 0.84310339979277, 0.85646046644909, 
    0.87036514247813, 0.88436233314301, 0.89862386081989, 0.91312712196071, 
    0.92808182875006, 0.94339952050624, 0.95900601011671, 0.97507187480826, 
    0.99159973087893,
  -0.99215854840574, -0.97670357961185, -0.96151388325688, -0.94670940351809, 
    -0.93217249638666, -0.91786485781008, -0.90387095749889, 
    -0.89003392144952, -0.87657670600548, -0.86340552589157, 
    -0.85017927922612, -0.8371936402569, -0.82418403783286, -0.8116716283968, 
    -0.79882710464895, -0.78659914463957, -0.775253775917, -0.76328297710881, 
    -0.75114939867018, -0.73965437862865, -0.72734463600681, 
    -0.71630706751133, -0.704822393902, -0.69365854567392, -0.68243884800439, 
    -0.67164083053832, -0.66089194174719, -0.64998481572728, 
    -0.63954171247384, -0.62848394020647, -0.61838790840236, 
    -0.60785761724231, -0.59801231122506, -0.58713167936608, 
    -0.5770805446205, -0.56644851789092, -0.55663557949282, 
    -0.54667777947224, -0.53717558595192, -0.52705795550772, 
    -0.51709917842265, -0.50792218349691, -0.49828216498647, 
    -0.48834889946522, -0.47881007466263, -0.46965810099996, 
    -0.46069178345217, -0.45030393315441, -0.44114608563709, 
    -0.4327056993955, -0.42278452763561, -0.41418171258613, 
    -0.40532410083788, -0.39579563046188, -0.38651881775653, 
    -0.37720495607383, -0.36845340660963, -0.35917287495774, 
    -0.35076116506919, -0.34187369198686, -0.33314111117715, 
    -0.32413857329849, -0.31528223522324, -0.30634452375124, 
    -0.29807860109232, -0.28904967562662, -0.28039044300494, 
    -0.27175006302276, -0.26299263002578, -0.25411330261377, 
    -0.2458335265964, -0.237362475327, -0.22953977146344, -0.22059290293124, 
    -0.21125820950021, -0.20318779022313, -0.19453084146962, 
    -0.18684586237701, -0.17798315668343, -0.16979508574896, 
    -0.16135392875564, -0.15273629828282, -0.14495641957907, 
    -0.13728488828314, -0.12792032286077, -0.11946496419327, 
    -0.11197344281973, -0.10378762165286, -0.095842828535383, 
    -0.087452003159811, -0.077991510656362, -0.070270811038522, 
    -0.062209368650508, -0.053796466519817, -0.045387944251733, 
    -0.036185395933304, -0.028223384681333, -0.020998298685471, 
    -0.012402796457678, -0.0036224836271044, 0.0037701633827351, 
    0.012181285549845, 0.021096506914874, 0.028702452076979, 
    0.037141143568948, 0.044773446694043, 0.053137253729735, 
    0.062419798793403, 0.070737566500326, 0.078629408300516, 
    0.086491678993176, 0.094297692997206, 0.10299538179262, 0.11127199650257, 
    0.11966780294033, 0.12746579478019, 0.1361990362859, 0.14488297044897, 
    0.15255493803288, 0.16111995162663, 0.16968533422984, 0.17835698923794, 
    0.18720581693188, 0.19510952611, 0.20342066678353, 0.21173853804177, 
    0.22021237078646, 0.22885170864412, 0.23759498379174, 0.24523702515653, 
    0.25456558475685, 0.26339520367861, 0.27235362610612, 0.28074422994168, 
    0.28876088073545, 0.29704970464196, 0.30640559651873, 0.31576971337924, 
    0.32420609946607, 0.33313246379073, 0.34151536548213, 0.35048791613926, 
    0.35971911447338, 0.36876875548576, 0.3774975191886, 0.3865573422544, 
    0.39610414900485, 0.40516009889337, 0.41338159795292, 0.42278363226227, 
    0.43193446677336, 0.44139892191655, 0.45071218663131, 0.45999828701222, 
    0.46994086996965, 0.4804899941114, 0.48859861743491, 0.49859720900232, 
    0.5081162973939, 0.51771708142685, 0.52714097230255, 0.53665250301933, 
    0.54686977462724, 0.55727776651305, 0.56772425809404, 0.57774327359169, 
    0.58755618144125, 0.59729294510205, 0.60787880961306, 0.61896981102219, 
    0.62945209092701, 0.63991243557011, 0.65070736110709, 0.66126470481986, 
    0.67192229278871, 0.68305487967449, 0.69473152304375, 0.70568485145922, 
    0.71719477269271, 0.72772633618378, 0.73984069517212, 0.75174270644503, 
    0.76344807696924, 0.77529230628369, 0.78727621062663, 0.79985005756739, 
    0.81207644128623, 0.82443253324882, 0.83747430549415, 0.85000987916033, 
    0.86337304481259, 0.87660492082209, 0.89009338443266, 0.90406599618947, 
    0.91805062594692, 0.9321571448925, 0.94674644975672, 0.96149667702771, 
    0.97666425320054, 0.99214494777523,
  -0.99257365415625, -0.9778039789183, -0.96335990806578, -0.9490524422007, 
    -0.93534362993725, -0.92118109395495, -0.90759944002621, 
    -0.89459164955089, -0.88172444125201, -0.8682735409381, -0.8556045122485, 
    -0.84289542525566, -0.83047176071319, -0.81825599996147, 
    -0.80542422066108, -0.79366879206023, -0.78187989222648, 
    -0.77039963524662, -0.75862431425874, -0.74685863482228, 
    -0.73533551809664, -0.72417874017814, -0.71268117204367, 
    -0.70162592467223, -0.69032898367585, -0.67963278927346, 
    -0.66867663840195, -0.65852931622492, -0.64770700226765, 
    -0.63670072813698, -0.62658315241175, -0.61605570905556, 
    -0.60559907041131, -0.59485607246133, -0.58555917339489, 
    -0.5751826447313, -0.56481046254902, -0.55457982007333, 
    -0.54526588527111, -0.53502896015911, -0.52484602297243, 
    -0.51579055034903, -0.5059444416664, -0.4959655447607, -0.48668049595576, 
    -0.4771924421653, -0.46761878753563, -0.45747951088917, 
    -0.44782529812891, -0.43862027522241, -0.43003798191113, 
    -0.42100721734066, -0.41106398943743, -0.40227107490138, 
    -0.39265087065804, -0.38417597736721, -0.3747120798106, 
    -0.36526489739369, -0.35640901838674, -0.34737438936549, 
    -0.33821513119673, -0.32971754924285, -0.32002583146416, 
    -0.31195733459964, -0.30333027121879, -0.2948848079043, 
    -0.28554051106341, -0.27633972975823, -0.26840978685816, 
    -0.25964900666989, -0.25127836187718, -0.24161578735199, 
    -0.23247276879076, -0.22470956396804, -0.21621597673102, 
    -0.20752494284037, -0.19904191741355, -0.19042858712986, 
    -0.18143267981416, -0.17301554427583, -0.16450145313967, 
    -0.15625612808527, -0.14794946406022, -0.13957717684361, -0.130294757413, 
    -0.1215931172936, -0.11399548158658, -0.10511462605933, 
    -0.096469507855956, -0.087819412631067, -0.079618349853686, 
    -0.071133140021428, -0.063062406870532, -0.055162285911743, 
    -0.046298159615174, -0.037892755774645, -0.029606969392753, 
    -0.020596782372998, -0.012548593152812, -0.0048127103828112, 
    0.0039059859455712, 0.012833916772137, 0.020455585904505, 
    0.029235253847958, 0.037311506528233, 0.045701498116605, 
    0.054224163082852, 0.063338098254692, 0.071452054208001, 
    0.079762889506684, 0.088572852761751, 0.096050814945958, 
    0.10495709001051, 0.11351688616595, 0.12281167067314, 0.13036056104903, 
    0.13884989562343, 0.14733489141509, 0.15530870643679, 0.16426156036062, 
    0.17244718114416, 0.18107859965013, 0.18988620694325, 0.19900305772366, 
    0.20683725359657, 0.21642528558692, 0.22479465368835, 0.23310971819058, 
    0.24207641032047, 0.25102067519038, 0.25937007168914, 0.26790672334642, 
    0.27643724950731, 0.28536792031031, 0.29448198740116, 0.30311643538381, 
    0.31218499445891, 0.32133411725402, 0.32968535343918, 0.33918041487997, 
    0.34770041688356, 0.35692336754758, 0.36600317808742, 0.37470171244851, 
    0.38441290843844, 0.39346680036885, 0.40316152562775, 0.41149943212898, 
    0.42083916984402, 0.43037635944934, 0.43905351931947, 0.44898569777505, 
    0.45735685034937, 0.46654113371757, 0.47661216348857, 0.48704596681495, 
    0.4967647664989, 0.50659328058205, 0.51619751793585, 0.52593387340949, 
    0.53495480073173, 0.54547656293051, 0.55568337332923, 0.56512315045443, 
    0.5756544017746, 0.58534531617381, 0.59560615961258, 0.60600175427874, 
    0.61613319890112, 0.62678280449228, 0.63750723396241, 0.64809108365081, 
    0.65904200797025, 0.66919414940231, 0.67987852310385, 0.69115252681146, 
    0.70265983155914, 0.71373049769875, 0.72455181075988, 0.73606481076912, 
    0.74731455634831, 0.75871715463969, 0.77034021073852, 0.78236480942198, 
    0.79438936893596, 0.80622895811497, 0.81827296425273, 0.83102081722804, 
    0.84325105311682, 0.85586677936078, 0.86858025069537, 0.88141407636822, 
    0.89468037859728, 0.90799601552262, 0.9215607909428, 0.93521013422458, 
    0.94919341750286, 0.96335154761359, 0.97784443043923, 0.99257056902782,
  -0.99285014376049, -0.97868961313554, -0.9647778996196, -0.95100619779317, 
    -0.93745753492922, -0.92413211770402, -0.9109113177994, 
    -0.89806813086023, -0.88502291111102, -0.87233948743487, 
    -0.85989892623959, -0.84757192265054, -0.83513579581006, 
    -0.8231422368118, -0.81099727808675, -0.79936796023896, 
    -0.78747584894776, -0.77570800966254, -0.7642936788168, 
    -0.75265744330134, -0.74148433277938, -0.73007560499528, 
    -0.71913770071942, -0.70808861889667, -0.69712789720924, 
    -0.68596844329645, -0.67536463548773, -0.66455333563425, 
    -0.65388087209966, -0.64366475566713, -0.63282464295457, 
    -0.62249346097378, -0.61226265764054, -0.60210487333418, 
    -0.59168437096343, -0.58152167132453, -0.57150345830781, 
    -0.56130829011504, -0.55180477944504, -0.54139772933291, 
    -0.53151331619986, -0.52178654269509, -0.5119050754815, 
    -0.50228969495088, -0.49279152571125, -0.48288932841867, 
    -0.47313956868041, -0.46399640959278, -0.45455132769683, 
    -0.4451298493573, -0.43548694981506, -0.42609177795201, 
    -0.41689767933391, -0.40723674328424, -0.39832458453619, 
    -0.38895482856438, -0.37994269501789, -0.37049462377906, 
    -0.36151387074136, -0.35269880307091, -0.34354440464222, 
    -0.33491363630898, -0.32521285285841, -0.31620921005502, 
    -0.30773522154578, -0.29899480113432, -0.28938709312182, 
    -0.28082964014594, -0.27174708628481, -0.2635551679981, 
    -0.25371165630272, -0.24575842318027, -0.23647645651229, 
    -0.22841033921341, -0.21895653570657, -0.21071413400189, 
    -0.20154813697023, -0.19287747770841, -0.18465461492541, 
    -0.17576592138315, -0.16730695159941, -0.15816608197078, 
    -0.14981617072819, -0.14132172248377, -0.13236869604949, -0.124222475957, 
    -0.11512715610394, -0.10688905497777, -0.098171317871739, 
    -0.09001347475743, -0.08068064778491, -0.073090910849317, 
    -0.063896636027597, -0.055412791083094, -0.047233187981829, 
    -0.038337442915541, -0.029985479306002, -0.021502899032519, 
    -0.012930718859328, -0.004224454271081, 0.0045926909256469, 
    0.012758227528275, 0.021899319513356, 0.029608056916988, 
    0.037813794768099, 0.046722340724665, 0.055750442425243, 
    0.063730652870903, 0.072376514463446, 0.081181225447641, 
    0.089940934784746, 0.098373482309791, 0.10657951423697, 0.11574609876302, 
    0.12369489668997, 0.13269558391968, 0.14124813600906, 0.14958503804362, 
    0.15799371579767, 0.16700971722231, 0.17545661609858, 0.18461481364769, 
    0.19320216619097, 0.20153099052182, 0.21043319003816, 0.21935560993933, 
    0.2280813117537, 0.23676547880739, 0.24555291703777, 0.25437708600248, 
    0.26326299705363, 0.27192350248692, 0.28074304688112, 0.29001083488825, 
    0.29863332091163, 0.3074581185102, 0.31628441216017, 0.32518916389011, 
    0.33497652745329, 0.34335112783667, 0.35285688320021, 0.3620463665488, 
    0.3712722575985, 0.37986090556483, 0.38968532715279, 0.39862454931342, 
    0.40798398339596, 0.4169848327501, 0.42647407775685, 0.43551013947718, 
    0.44547928326807, 0.45462708422974, 0.46429432138963, 0.47417398064372, 
    0.48362673076369, 0.49291134335296, 0.5025569176657, 0.51244616935962, 
    0.52188260156425, 0.5319670603699, 0.54165168759799, 0.55204186674614, 
    0.56173102668766, 0.57219447566255, 0.58227137390751, 0.59236622252176, 
    0.60265925055563, 0.61267145985974, 0.62297479928976, 0.63338597681282, 
    0.64383510497963, 0.65460229882432, 0.66486947694406, 0.67607784512356, 
    0.68685712621674, 0.69777833421161, 0.70851545982683, 0.71965297809083, 
    0.73049430025626, 0.74183707023416, 0.75337406635386, 0.7646861117972, 
    0.77620470907049, 0.78792071527968, 0.79954601951793, 0.81129177373901, 
    0.8232987911078, 0.83561409610274, 0.84752649024134, 0.86016205842851, 
    0.87252137520138, 0.8852418218626, 0.8980832269476, 0.91100365104669, 
    0.9242159691796, 0.93755358379692, 0.95104494413873, 0.96473587740162, 
    0.97869986844368, 0.99284967536575,
  -0.99309040310612, -0.97937469128936, -0.96587388969378, -0.95249946619003, 
    -0.93924327420484, -0.92630843475382, -0.91340812198918, 
    -0.90069876467589, -0.88820291730819, -0.87575971664562, 
    -0.86330217403407, -0.85118873663105, -0.83897967581159, 
    -0.82724064532363, -0.81538297539072, -0.80334136135333, 
    -0.79184221448902, -0.78015969170914, -0.76896670193581, 
    -0.75773030224319, -0.74644848520939, -0.73528364905804, 
    -0.7243177821947, -0.71307629391937, -0.70235513743883, 
    -0.69155464876151, -0.68078531026928, -0.6698768098602, 
    -0.65946172395243, -0.64842220349982, -0.63786131680445, 
    -0.62790660058271, -0.61774269149561, -0.60736126114361, 
    -0.5970542564739, -0.58711941723172, -0.57714160084535, -0.566953029848, 
    -0.55700304786554, -0.54656729513298, -0.536901184032, -0.52726237101953, 
    -0.51743850578043, -0.50783072212159, -0.49780072437379, 
    -0.4880741873479, -0.47850220244848, -0.46854933638319, 
    -0.45919300785736, -0.45005521552603, -0.44022468725678, 
    -0.43070981881157, -0.42175463935794, -0.41219030249231, 
    -0.40316611620091, -0.39373656426385, -0.38413402792777, 
    -0.37543904091549, -0.36539511856223, -0.3567206288179, 
    -0.34782698916392, -0.33852077948691, -0.32938166270825, 
    -0.32009593773197, -0.31161911470114, -0.30218928850519, 
    -0.29331510767116, -0.28416793593339, -0.27538106880388, 
    -0.26634776509921, -0.25746021151201, -0.24894471395247, 
    -0.23992433538526, -0.23080522997755, -0.22197560287641, 
    -0.2129895822754, -0.20385561586969, -0.19541226968624, 
    -0.18710615304658, -0.17781990904378, -0.1691706661918, 
    -0.16050962325151, -0.1515098949688, -0.14261961874289, 
    -0.13435470421539, -0.12536798663871, -0.11685731714002, 
    -0.1083842720115, -0.10011955493754, -0.091088073199454, 
    -0.082359026492248, -0.073979320096099, -0.065192180028116, 
    -0.056081854451854, -0.047420792038979, -0.039140355173066, 
    -0.030129436453745, -0.02173560665213, -0.012473054726098, 
    -0.0039178690360861, 0.0045672324997395, 0.012900090173538, 
    0.02153786243278, 0.030385523859355, 0.038930959732244, 
    0.047356161421105, 0.056225348043927, 0.06465251431448, 
    0.073513543708058, 0.082216918791103, 0.090750956676091, 
    0.099127463318193, 0.10756996518594, 0.11709069435445, 0.12552015079918, 
    0.13403408273964, 0.14279578891615, 0.15156137461709, 0.16033295190101, 
    0.16931928429838, 0.17825840820056, 0.18696913946355, 0.19576631363669, 
    0.20432867987057, 0.21342922073364, 0.22226249699308, 0.23091322463481, 
    0.24005752937435, 0.24864119869045, 0.25744681959139, 0.26623457086256, 
    0.27504207204405, 0.28438023120007, 0.29330385917273, 0.30231170205504, 
    0.31146460102546, 0.32030964147406, 0.32985308289998, 0.33847716347148, 
    0.34754529483462, 0.35630077679753, 0.36600430840028, 0.37511675965296, 
    0.38469312941166, 0.39355526289659, 0.40348106136443, 0.41313528260116, 
    0.42165026036623, 0.43135397714191, 0.44071766414746, 0.44964857010502, 
    0.45969771875274, 0.46951388353792, 0.47894010177474, 0.48865348673984, 
    0.49830410207523, 0.50762346849459, 0.5180518840724, 0.52742930291741, 
    0.53770397417751, 0.54735835775067, 0.55702320657369, 0.56683975966024, 
    0.57748861735902, 0.58784590466046, 0.59769835494591, 0.60793164486123, 
    0.61847187459381, 0.62841570799488, 0.63887796034629, 0.64940283210101, 
    0.65980505763901, 0.67070449550353, 0.68104278312366, 0.69191098600327, 
    0.7026960038686, 0.71386057078954, 0.72454990237214, 0.73590343972295, 
    0.7466215254499, 0.75811863636803, 0.76944997441264, 0.7808913933585, 
    0.79242156672996, 0.80364804973049, 0.8156364986653, 0.82749936452362, 
    0.83950283080479, 0.85122677408178, 0.86365592355834, 0.87587621675112, 
    0.88814331082639, 0.90091425605959, 0.91352215868231, 0.92632288664359, 
    0.93937767979685, 0.95251446923167, 0.96584357394754, 0.97937740242547, 
    0.99308333833611,
  -0.99343145087519, -0.98036771478283, -0.96745653235616, -0.95472769897786, 
    -0.94199932994437, -0.9295600322072, -0.91710782930083, 
    -0.90480447566311, -0.89263792583526, -0.88058375830773, 
    -0.86861204788585, -0.85678204147727, -0.84489719997123, 
    -0.83322686041088, -0.82179838842546, -0.8102164792888, 
    -0.79881275634032, -0.78742800380881, -0.7762922721026, 
    -0.76499091620254, -0.75389020123155, -0.742948256762, -0.73207945084601, 
    -0.72110693474147, -0.71027355986621, -0.69962527571924, 
    -0.68873880943783, -0.67828352612092, -0.66792344444865, 
    -0.65721223125237, -0.64681007161156, -0.63635712218256, 
    -0.62606793293416, -0.61584912637779, -0.60576708040287, 
    -0.59510284623158, -0.58536047273012, -0.57531741098521, 
    -0.56512415417121, -0.55540133391975, -0.54530138470253, 
    -0.53564757982995, -0.52536858221825, -0.51572175304355, 
    -0.50591983891254, -0.49628243482924, -0.4863601316208, 
    -0.47682243731073, -0.46705268312506, -0.45772688508165, 
    -0.44795149325434, -0.43833474097015, -0.42930754325978, 
    -0.41964629966455, -0.41032161458276, -0.40050374237371, 
    -0.39120382029386, -0.38207041065493, -0.37292858064857, 
    -0.36325000189348, -0.35420817435735, -0.34478047603172, 
    -0.33564347019782, -0.32590579067721, -0.31746561135188, 
    -0.30792051727886, -0.29903304115627, -0.28969623721568, 
    -0.28072316010133, -0.27167289441814, -0.26247585807441, 
    -0.25364403334043, -0.2443638789392, -0.2356934909102, -0.22647232041783, 
    -0.21720064985639, -0.20831975674204, -0.19968338800892, 
    -0.19044992457224, -0.18221708139609, -0.17286528219449, 
    -0.16391137131918, -0.15465821832105, -0.14585050737497, 
    -0.13728450691301, -0.12786212035015, -0.11895454279165, 
    -0.1107446443415, -0.10161183890339, -0.09270010907311, 
    -0.083770270414693, -0.074760381153161, -0.066092061316995, 
    -0.057019265148772, -0.048817218119538, -0.039828218916875, 
    -0.031218544910523, -0.022287742669593, -0.013326448954305, 
    -0.0046072771996463, 0.0046909900004664, 0.013100349131882, 
    0.022526987110081, 0.030944368216132, 0.03963735775619, 
    0.048388173775299, 0.057135405745491, 0.066207351961981, 
    0.07513895838019, 0.083706640082191, 0.09253478800231, 0.10136146456962, 
    0.1104896398616, 0.11924988975928, 0.12790490854369, 0.13660214463483, 
    0.1460740902215, 0.154585743021, 0.1637670284091, 0.17224025900559, 
    0.18158686227357, 0.19065033192706, 0.19961771597629, 0.20867126793016, 
    0.21736602236978, 0.22650285001134, 0.23546708416974, 0.24461189057416, 
    0.25330968603473, 0.26241392185582, 0.27140856855843, 0.28023554038731, 
    0.2900220477139, 0.29918350736978, 0.30841930959018, 0.31746829368522, 
    0.32609630375743, 0.33584740999841, 0.3448922280826, 0.35404331761415, 
    0.36365769191378, 0.37285120571084, 0.38203654096373, 0.39196000199899, 
    0.40066875121345, 0.4104636628603, 0.41979577830146, 0.42935890773794, 
    0.43888630649282, 0.44844994152367, 0.45783075471919, 0.46758676521883, 
    0.47738602471811, 0.48700623202762, 0.49668259652842, 0.50604571860708, 
    0.51605682027962, 0.5259164048654, 0.53605299367084, 0.54577925563717, 
    0.55566259077662, 0.56586351149801, 0.57557503564277, 0.58592737087442, 
    0.59614383783425, 0.60620262873067, 0.6164285609496, 0.62686260264964, 
    0.63705050717573, 0.64737189029891, 0.65771425892021, 0.66823245109949, 
    0.67890447435562, 0.68929398375688, 0.70015829704236, 0.71110965611897, 
    0.72165461858795, 0.73249125261147, 0.74344794531759, 0.7545085381835, 
    0.76552150922133, 0.77661149492123, 0.78785576690392, 0.79915323692038, 
    0.81050068742048, 0.82209115417866, 0.83356270603341, 0.8452391648201, 
    0.85699814289896, 0.86889955201606, 0.88075587602587, 0.89274459425727, 
    0.90495701016881, 0.9172734729899, 0.92956521994316, 0.94212046870675, 
    0.95468088441398, 0.96749205634089, 0.9803834706314, 0.99343379073794,
  -0.99356383390551, -0.98076327758803, -0.96812203149109, -0.95548683577404, 
    -0.94300239997147, -0.93066836139317, -0.91865705237225, 
    -0.90653912954282, -0.89444208192812, -0.88242584550808, 
    -0.8708176684121, -0.85887131278182, -0.84727063233603, 
    -0.83556600928436, -0.82397190729378, -0.81265576194235, 
    -0.80127505515786, -0.79032529103459, -0.77905849984626, 
    -0.76817840523939, -0.75689748106988, -0.74614046793975, 
    -0.7352225984219, -0.7241539228555, -0.71328130780955, -0.70230388917833, 
    -0.69178612751298, -0.68163977829941, -0.67142359126423, 
    -0.66091859712498, -0.65074798647586, -0.63970503562992, 
    -0.62955508950155, -0.61925955190573, -0.60873580108172, 
    -0.59928176595763, -0.58877228099324, -0.57823097210717, 
    -0.56863633636557, -0.5583099136866, -0.54913524487792, 
    -0.53860859536648, -0.52877264224818, -0.51851133334955, 
    -0.50918392265068, -0.49905796958184, -0.48916569832939, 
    -0.48016795608805, -0.47026834593403, -0.46023930646042, 
    -0.4509426323064, -0.44132249368771, -0.43208307275097, 
    -0.42291787731041, -0.41301875903945, -0.4030188151183, 
    -0.39340694039576, -0.38463546378559, -0.37533955676198, 
    -0.36653313055515, -0.35664315672271, -0.34728809550224, 
    -0.33875579748423, -0.32910978003646, -0.31980425351662, 
    -0.31061938645261, -0.30135150384068, -0.29210634762556, 
    -0.28324345064603, -0.27404111321111, -0.2646379252988, 
    -0.25478778017637, -0.24596470534256, -0.23732324149063, 
    -0.22855846821387, -0.21898712311736, -0.21026203933831, 
    -0.2012734057917, -0.1920040708468, -0.18341732932738, -0.17383104339228, 
    -0.16480848044184, -0.15541879055013, -0.14644959681356, 
    -0.13799691403146, -0.12923709571625, -0.12047877657914, 
    -0.11134142780778, -0.10278306446629, -0.093150135031595, 
    -0.084666677892009, -0.075479326366053, -0.066714392612804, 
    -0.058315677039863, -0.04915531525756, -0.040306926668488, 
    -0.031585865469236, -0.022554426305368, -0.013838684029823, 
    -0.0037944736870812, 0.0043150206099967, 0.013634588688566, 
    0.021495157132242, 0.030261094148125, 0.039490107480695, 
    0.048617332487718, 0.058136899282365, 0.067041986589286, 
    0.075761790438314, 0.084032215431661, 0.093439848086947, 
    0.10294053395531, 0.11070941195818, 0.11990210849808, 0.12980051530081, 
    0.13767930057004, 0.14658502209111, 0.15605915406052, 0.16553928761623, 
    0.17408891850617, 0.18344848251608, 0.19142403130546, 0.20075943539717, 
    0.21059863988655, 0.21886763246713, 0.22879627552835, 0.23766340124126, 
    0.24612835557219, 0.25517668224529, 0.26426494343583, 0.27365982171593, 
    0.28282850446588, 0.29254776513907, 0.3012749571621, 0.31068933815811, 
    0.3197541619212, 0.32860963480642, 0.33893889995858, 0.34768969605491, 
    0.35680627643638, 0.36637393612756, 0.37530833180642, 0.38478452696195, 
    0.3944180126319, 0.40388994763104, 0.41316173236629, 0.42275262123304, 
    0.43231262593907, 0.44152801422237, 0.45135759272941, 0.46027206465753, 
    0.47103867015133, 0.48081120457027, 0.49054307445699, 0.49983494468191, 
    0.50986714927602, 0.51981626028905, 0.52959259249218, 0.53931294721724, 
    0.54843401645975, 0.55884614017345, 0.56905423743047, 0.57926734152125, 
    0.5893121786155, 0.59907082137042, 0.60899556127647, 0.61942121561275, 
    0.63047548370109, 0.64063105328979, 0.65098663895843, 0.66112595314741, 
    0.67174512292863, 0.68236187277808, 0.69280168620016, 0.70296706163397, 
    0.71390645294931, 0.72469241725787, 0.73562576840084, 0.7465393071587, 
    0.75717649479434, 0.76855200491486, 0.77962685278313, 0.79066661513112, 
    0.80202352173663, 0.81300635238487, 0.82452644952804, 0.83608676194653, 
    0.8473604017122, 0.85924586140342, 0.87099037240498, 0.88249696043007, 
    0.89450028172969, 0.9065499135713, 0.91860278881723, 0.93088314934455, 
    0.94317151292919, 0.95559595194204, 0.96807406295879, 0.98076551139889, 
    0.9935667857524,
  -0.99366914105123, -0.98108019169525, -0.96859399488361, -0.95624356771207, 
    -0.94398184381652, -0.93179705535383, -0.91968963450832, 
    -0.90774362076136, -0.89583378352846, -0.88406912651065, 
    -0.87240255666491, -0.86064792234411, -0.84927370394806, 
    -0.83774167992301, -0.82643019027284, -0.81484907085771, 
    -0.80380200279797, -0.79258295703599, -0.78156221859223, 
    -0.77047782856748, -0.75954731881826, -0.74855310971179, 
    -0.73755497765331, -0.72717660624724, -0.71629646530584, 
    -0.70561117864784, -0.694791560896, -0.6843623205326, -0.67403956506401, 
    -0.66342067448634, -0.6531148590657, -0.64274617120881, 
    -0.63223726344032, -0.62212984080063, -0.61196612259328, 
    -0.60170722778572, -0.59161888334446, -0.58131056374738, 
    -0.57162973732992, -0.56151282162987, -0.5513629791442, 
    -0.54183768788931, -0.53192094266543, -0.52169314871516, 
    -0.51197528093828, -0.50233542045542, -0.49240659106037, 
    -0.48278840097584, -0.47296495213985, -0.46348914810011, 
    -0.45383061893518, -0.44441531440314, -0.4344728724651, 
    -0.42535712805848, -0.41571713811398, -0.40602035001241, 
    -0.39648107143741, -0.3874088404207, -0.37772059662755, 
    -0.36798414750615, -0.35894958358253, -0.35015958003607, 
    -0.34035198340436, -0.33115620102601, -0.32182063258019, 
    -0.3124449430212, -0.30339964437222, -0.29358847688861, 
    -0.28468314574215, -0.27574242031809, -0.26629687438451, 
    -0.25747933104385, -0.24791982507155, -0.2391737579313, 
    -0.22969035669472, -0.22075453719972, -0.21146002009868, 
    -0.2023286906839, -0.19314058791739, -0.18419202787862, -0.1757963054725, 
    -0.16656390728252, -0.15725821805484, -0.14804560965134, 
    -0.13921634837604, -0.13005820730729, -0.12130874055874, 
    -0.11210698703903, -0.10304963101019, -0.094731121504546, 
    -0.085237283094065, -0.076051309087717, -0.066882716718367, 
    -0.058436690334734, -0.049465137374333, -0.040345316060418, 
    -0.031672944313127, -0.022335711929155, -0.013372983057397, 
    -0.0045461273848757, 0.0046231360644512, 0.013416843740076, 
    0.022487779335105, 0.031369423844848, 0.040267410485159, 
    0.049135115532125, 0.05808056778538, 0.06674439718505, 0.076242926547719, 
    0.085177465947494, 0.094020446991357, 0.10319179615885, 0.11188509507253, 
    0.12107741064751, 0.13000939781116, 0.13914528007327, 0.14824159853897, 
    0.15681397563457, 0.16618083726377, 0.17484375968677, 0.18410339192939, 
    0.19333873455982, 0.20269729992106, 0.21159070801773, 0.22028200625379, 
    0.23011311439388, 0.239071965636, 0.24810343948504, 0.2573405703824, 
    0.26617566434815, 0.27530090997847, 0.28496803809064, 0.29396024682156, 
    0.3034234258294, 0.31252553120878, 0.32161412472966, 0.33125671514541, 
    0.34053898632202, 0.34989062491116, 0.35906764234899, 0.36861729570498, 
    0.37783456217433, 0.38726030890568, 0.39677922994395, 0.40631447324038, 
    0.41588555326076, 0.42549631310688, 0.43485163741667, 0.44465794877651, 
    0.45433394285272, 0.4638786237059, 0.47325938360306, 0.48308249549214, 
    0.49295847776273, 0.50282088159326, 0.51244137907074, 0.52226332025718, 
    0.53214024151923, 0.54187339757703, 0.55209705702746, 0.5619444924466, 
    0.57176771203575, 0.58227430105485, 0.59208408378074, 0.60236824972735, 
    0.61244508310611, 0.62270828887921, 0.63288734661111, 0.64344936743776, 
    0.65359538554875, 0.6640080471247, 0.67436015063395, 0.68511008471418, 
    0.69539585509858, 0.70620078143614, 0.71676968747448, 0.72745757137354, 
    0.7382415996964, 0.74904774745127, 0.75989584107387, 0.77094049194006, 
    0.78192187884571, 0.79312666895582, 0.80415326557574, 0.81534534109103, 
    0.82670615071618, 0.83804627291271, 0.84945721261926, 0.86097148490463, 
    0.87259624641572, 0.88421403065222, 0.89606217590857, 0.90785476750637, 
    0.91984843052088, 0.93187139351622, 0.94402769528426, 0.95626727992643, 
    0.96862229169415, 0.98109731882669, 0.99367275320645,
  -0.99385040865217, -0.98161546391631, -0.96939128741968, -0.95738516013299, 
    -0.94540522354895, -0.93346583473094, -0.92183586270775, 
    -0.90987492843385, -0.89812555805371, -0.88674383542425, 
    -0.87534000716568, -0.86391476122439, -0.85237432309991, 
    -0.84097956693298, -0.8299053410042, -0.81871690026464, -0.8073626610683, 
    -0.7963930985602, -0.78548430564195, -0.77461594157252, 
    -0.76389888602268, -0.75278359444227, -0.74193668282836, 
    -0.73167185147873, -0.72131383675932, -0.71000495278865, 
    -0.69931862756085, -0.68941163877577, -0.6786849669596, -0.6686562631557, 
    -0.65774308815796, -0.64797053070836, -0.63737959096717, 
    -0.62676132738367, -0.61662191759491, -0.6063596837864, 
    -0.59653369920325, -0.58593027803995, -0.57659557486043, 
    -0.56652061438535, -0.55656793234383, -0.54623887678638, 
    -0.53661894612861, -0.52684827534047, -0.51658227857825, 
    -0.50642654747155, -0.49729110354526, -0.48770570637764, 
    -0.47753245607918, -0.46806745163191, -0.4582485480475, 
    -0.44863144415468, -0.43854421223775, -0.42945612152883, 
    -0.41993681430984, -0.41039285385515, -0.40062475263016, 
    -0.39134282519769, -0.38150275076894, -0.37188538605705, 
    -0.3626242276989, -0.35337446257157, -0.34426765136294, 
    -0.33499229215568, -0.32571642248592, -0.31581166308092, 
    -0.30635326821633, -0.29710589513253, -0.28803042951886, 
    -0.27883166032241, -0.26948451842503, -0.26059280205388, 
    -0.25083475284004, -0.2420151150092, -0.23275122524887, 
    -0.22276596421583, -0.2143183309486, -0.20554385832719, 
    -0.19579602950945, -0.18636979164913, -0.1769333491735, 
    -0.16827199457388, -0.15870872680627, -0.14965478318922, 
    -0.14116300849207, -0.13197138545509, -0.12301364801434, 
    -0.1135119005495, -0.10469920431668, -0.094994729672992, 
    -0.085719194846861, -0.076883697701234, -0.068193177095699, 
    -0.058938950541837, -0.049550842895838, -0.040555716122704, 
    -0.031922274984684, -0.023103163145992, -0.013720064131343, 
    -0.0044493320313421, 0.0046662509674713, 0.01394400602185, 
    0.022224105393607, 0.03171088913255, 0.040769608032948, 
    0.050104374412568, 0.059358929866126, 0.067715516418066, 
    0.077433521397918, 0.085682321610093, 0.094771158748932, 
    0.10438029133127, 0.11318364489269, 0.12208644767944, 0.13096736081258, 
    0.14076995829621, 0.15068879099671, 0.15955274472774, 0.1680363768192, 
    0.17754490938056, 0.18646810251546, 0.19507575263912, 0.20445124094464, 
    0.21382248326065, 0.22348118908405, 0.23309520095819, 0.24206629780127, 
    0.25090296751639, 0.25976174562257, 0.26958562175229, 0.27820365828175, 
    0.28802046973394, 0.29716951082417, 0.30677079324533, 0.31626592996642, 
    0.3254504360813, 0.33489187449618, 0.34363812246894, 0.35322949639153, 
    0.36290851454733, 0.37221036389131, 0.3818778128013, 0.39160195739719, 
    0.40108930970852, 0.41033961702186, 0.41983870754352, 0.42965311314849, 
    0.43910669401449, 0.4486209594459, 0.45912979733468, 0.46850546165462, 
    0.47828948424682, 0.48782632229152, 0.49768624577784, 0.50732027765092, 
    0.51676607713233, 0.52702746385295, 0.53660614048192, 0.54674707597093, 
    0.55694813274555, 0.56680150475402, 0.57696115433654, 0.58713779705715, 
    0.59642218039505, 0.60672716023495, 0.61732010347163, 0.62788850806407, 
    0.6377772019533, 0.64781969366452, 0.65848554032422, 0.66877777772228, 
    0.67921752274492, 0.68949005168825, 0.69992189879771, 0.71081021127791, 
    0.72141512168961, 0.73181363250108, 0.74254149824165, 0.75351227915839, 
    0.76434470227234, 0.77494930121205, 0.78591836959534, 0.79647798531888, 
    0.80807084827741, 0.81915107721088, 0.82997102189787, 0.84148333188971, 
    0.85288252141836, 0.86403307265124, 0.87535868960112, 0.8867786073457, 
    0.89834854631173, 0.91010560194242, 0.92174512897687, 0.93368206410929, 
    0.94544038441102, 0.95740849534932, 0.96954374370737, 0.98158413217396, 
    0.99384486794639,
  -0.99398495592566, -0.9819939540589, -0.9701193832702, -0.95820868305897, 
    -0.94650430751953, -0.93485008216519, -0.92316561240917, 
    -0.91163684926954, -0.90018252822302, -0.88889220667366, 
    -0.8773954205619, -0.86600690575791, -0.85480233179349, 
    -0.84370976381651, -0.83264098221297, -0.82159826048544, 
    -0.81047775543124, -0.79953841332968, -0.78876910928717, 
    -0.77793948243788, -0.76704567954047, -0.75637962967836, 
    -0.74572152559093, -0.7349264419796, -0.72430940768217, 
    -0.71389117090895, -0.70327732986617, -0.69291501494023, 
    -0.68259533173031, -0.67211353555352, -0.66171406201083, 
    -0.65130155643703, -0.64107019584302, -0.63088202564025, 
    -0.62117922175702, -0.61035152801926, -0.60046763468953, 
    -0.58999867459615, -0.58008102953987, -0.5702670015192, 
    -0.56038403682332, -0.5502998546562, -0.54025442366108, -0.5304302344064, 
    -0.52042800836601, -0.5106650150134, -0.50128950486811, 
    -0.49116464832791, -0.48118362547695, -0.47160759540899, 
    -0.46195387296525, -0.45256096372678, -0.44265359509158, 
    -0.43302180861406, -0.42352233249491, -0.41382553719991, 
    -0.40393408165426, -0.39463347368704, -0.38478771893126, 
    -0.37533790245916, -0.36608069502031, -0.35657519903132, 
    -0.34722151019841, -0.337346702521, -0.32812221139485, -0.31839303886494, 
    -0.30961521515454, -0.30006126307075, -0.29070783321792, 
    -0.28132304921321, -0.27209967968581, -0.26276515387149, 
    -0.25298096135689, -0.24379436710483, -0.23488077024436, 
    -0.22511896308444, -0.21618461754117, -0.20703983340345, 
    -0.19800781068997, -0.18810645740461, -0.17869135541607, 
    -0.16974735213598, -0.16083019291443, -0.15124025973726, 
    -0.14162836932395, -0.13262356459465, -0.12376729774127, 
    -0.11511558487273, -0.10524872545302, -0.096312999481282, 
    -0.087154342040601, -0.077953178527688, -0.068663933892985, 
    -0.05984041001269, -0.050566910099655, -0.041286030831279, 
    -0.032008778244722, -0.023037455315202, -0.01366049741305, 
    -0.0044606757507033, 0.0044540520057654, 0.014067056312708, 
    0.023377770437073, 0.031884390611936, 0.040799045809538, 
    0.050430342762398, 0.05943039406286, 0.06760210036102, 0.07769122404257, 
    0.087070284999211, 0.096199180418113, 0.10510031361825, 0.11454373137204, 
    0.12353196082126, 0.13337543639709, 0.14190334426254, 0.15166871424939, 
    0.16079899132132, 0.16961789614214, 0.17891430773511, 0.18854719563441, 
    0.19750954326191, 0.2070109715933, 0.21622613914701, 0.22517905456587, 
    0.23469888511492, 0.24391513910029, 0.25342624276365, 0.26237789600945, 
    0.27192303317202, 0.28093489966329, 0.2903418144933, 0.30007794722168, 
    0.30955292061218, 0.31889228618241, 0.32794458123017, 0.33791337149275, 
    0.34718343058479, 0.35679928212969, 0.36643532813715, 0.37580981191904, 
    0.38483770150301, 0.3947101936597, 0.40413493532073, 0.41424345855112, 
    0.42346556127275, 0.43344574484679, 0.44245261298519, 0.45264226481424, 
    0.46212239867657, 0.47181359134228, 0.48173507873097, 0.49155961342908, 
    0.50112530708457, 0.51103419979586, 0.5209977429653, 0.530887402078, 
    0.54069418161129, 0.55102636982279, 0.56070426458843, 0.57083342132162, 
    0.58058370156583, 0.59049166375098, 0.60107132566901, 0.61101402528813, 
    0.6212299760568, 0.63126057200022, 0.6415998641439, 0.65195613669118, 
    0.66226461314827, 0.6723581884877, 0.68295615179428, 0.69337390432959, 
    0.703749624999, 0.71425201103383, 0.72459253711087, 0.73543604982662, 
    0.74603075636141, 0.75683498726286, 0.76741840271507, 0.77823351646893, 
    0.78895978838181, 0.79997091885944, 0.81084663937104, 0.8219237636377, 
    0.83267672904781, 0.84393590306392, 0.85513071598996, 0.86639345886497, 
    0.87744693639993, 0.88902949704156, 0.90023399035708, 0.91174279961083, 
    0.92327218730205, 0.93488717279198, 0.94653016245455, 0.95831735609605, 
    0.97009759089591, 0.98200612987793, 0.9939906973869,
  -0.99409289916428, -0.98231604044492, -0.97060134619091, -0.9589738528881, 
    -0.94737014687003, -0.93582934655026, -0.92443926469246, 
    -0.91298131256944, -0.90168105239433, -0.89035581754691, 
    -0.87917595090593, -0.86804273067432, -0.85683259535696, 
    -0.84585399452964, -0.8348292352737, -0.82372778445438, 
    -0.81286752577374, -0.80218554709358, -0.79128860848304, 
    -0.78047050824226, -0.76962955795867, -0.75922053248787, 
    -0.74839609126337, -0.73779656872647, -0.72725823832325, 
    -0.71667217436339, -0.70643562406311, -0.69580603091183, 
    -0.68544525972419, -0.67511382058317, -0.6647495467339, 
    -0.65467073584959, -0.64429160586007, -0.63395657502512, 
    -0.62387589069642, -0.61366828125431, -0.60343315636669, 
    -0.59356602203956, -0.58331493977761, -0.57363473074558, 
    -0.56321604221436, -0.55355088435868, -0.54362354780151, 
    -0.53347296656677, -0.52365363142575, -0.51396337090706, 
    -0.50401952474927, -0.49390088418509, -0.48457125597131, 
    -0.47486231550428, -0.46488403286467, -0.45525242810402, -0.445476894443, 
    -0.43564181038317, -0.42608229081081, -0.41624990985609, 
    -0.40656456644621, -0.3972596078141, -0.38778055394292, 
    -0.37806573264227, -0.36838241190368, -0.35897086956925, 
    -0.34970442973042, -0.34005872315934, -0.33084060483561, 
    -0.32104587368696, -0.31166634015716, -0.3021745819495, 
    -0.29223926555371, -0.28300790952792, -0.27403194559488, 
    -0.26467253786921, -0.25539523630274, -0.24596081260583, 
    -0.23659744742554, -0.22731926284219, -0.21735836849384, 
    -0.20825283239033, -0.19898732566721, -0.18969084027969, 
    -0.18041097736942, -0.17105575858193, -0.16231706958522, 
    -0.15252237257976, -0.14318971552913, -0.13398034306752, 
    -0.12466531390889, -0.11563072260722, -0.10637142833837, 
    -0.096878992103397, -0.087693013016126, -0.078890977764896, 
    -0.069222989229477, -0.05988220565574, -0.050910214147262, 
    -0.041403250550455, -0.032289119861203, -0.023168792030359, 
    -0.013732959534616, -0.0047805336596984, 0.0047271949707866, 
    0.013603704919235, 0.022725308768011, 0.032245482864996, 
    0.041467329931901, 0.050790767295076, 0.059812570494623, 
    0.069148104314588, 0.07862799148518, 0.087564276885082, 
    0.096858973857551, 0.1063112691504, 0.11525453245091, 0.12492650618966, 
    0.13423531731093, 0.14326599770538, 0.15245899345825, 0.16184345298825, 
    0.17059281455462, 0.18028342966562, 0.18980531533877, 0.19867754641696, 
    0.20839788057197, 0.21795590698966, 0.2269960598263, 0.23665661601097, 
    0.24616140697251, 0.25475899150138, 0.26476706360917, 0.27423939726555, 
    0.28354060302262, 0.29259967116887, 0.30216418306074, 0.31154945652495, 
    0.32096751052425, 0.33063212488423, 0.34043152889644, 0.34968001712968, 
    0.3587524069736, 0.36854637426911, 0.3785804463909, 0.38790191314318, 
    0.39728821659099, 0.40712434962887, 0.41685390481153, 0.42631495235858, 
    0.43619083937621, 0.4457011021068, 0.45560912706783, 0.46516288131078, 
    0.47514148753344, 0.48456517184673, 0.49445111324673, 0.5041647514953, 
    0.51427128118071, 0.52401319167343, 0.53412698579786, 0.54415952927043, 
    0.55386290856738, 0.5637034514786, 0.57366387536172, 0.58401279181823, 
    0.5939270379302, 0.60391512636943, 0.61427812337566, 0.62416694695246, 
    0.63436740680102, 0.6447781636385, 0.65486754548726, 0.66529765827859, 
    0.67549720531054, 0.6858753521349, 0.69630286990541, 0.70669822476138, 
    0.71722283737735, 0.72755456692483, 0.73828370593115, 0.74877198610281, 
    0.7595073237934, 0.77000108417518, 0.78084659942501, 0.79155400345003, 
    0.80235219683874, 0.81324324389356, 0.8241281338036, 0.83494035766584, 
    0.84602052995629, 0.85704359030432, 0.86817213941786, 0.87929984490311, 
    0.89048485619223, 0.90177584848633, 0.91311482691847, 0.92446520261272, 
    0.9359164691994, 0.94738373953114, 0.95899408608731, 0.9706191719833, 
    0.98231824020209, 0.9940936899903,
  -0.9941769486715, -0.98256346231029, -0.97103421400714, -0.95951094413088, 
    -0.94808772030483, -0.93671918791483, -0.92535660068957, 
    -0.91410380445202, -0.9029233764834, -0.89169234353832, 
    -0.88063790472035, -0.86949413525616, -0.85850009071584, 
    -0.84754704062621, -0.83669688903745, -0.82559020910295, 
    -0.81497094237783, -0.80401769518886, -0.79337240926063, 
    -0.78259087151219, -0.77201029560246, -0.76130177262207, 
    -0.75072072706565, -0.74018489537065, -0.72977057712797, 
    -0.71916295928217, -0.70879714946573, -0.69837317018768, 
    -0.68791482726352, -0.67772511835401, -0.66750154774865, 
    -0.65706602134573, -0.64699085433479, -0.63676825491244, 
    -0.62636162371826, -0.61632944534219, -0.60629409956818, 
    -0.59613079558985, -0.58598132002373, -0.57605298782507, 
    -0.56602693014941, -0.55593854000638, -0.5461194385608, -0.5360845003997, 
    -0.52636212037458, -0.51642968299323, -0.50659150537878, 
    -0.49684011171258, -0.48644822283554, -0.47707298411648, -0.467408019021, 
    -0.45758895100504, -0.44769723778399, -0.43817331699555, 
    -0.42825359586641, -0.41857702093601, -0.40911526472044, 
    -0.39944422080508, -0.38985351595569, -0.38024920755491, 
    -0.37061705659236, -0.36143655393212, -0.35158584771764, 
    -0.34199692509562, -0.33241724234726, -0.32290966281169, 
    -0.31360985533224, -0.30380553456723, -0.29435460664488, 
    -0.28523633214719, -0.27598033195216, -0.26635270319301, 
    -0.25627170632485, -0.24718927307389, -0.23792674033759, 
    -0.22861511108405, -0.2188445552574, -0.2097024931598, -0.20035735744581, 
    -0.19085996610437, -0.18153046327922, -0.17234135552599, 
    -0.16300510779283, -0.15346458852976, -0.14437041781349, 
    -0.13469019917796, -0.12558275861074, -0.11624622506518, 
    -0.10707896134897, -0.097275341075785, -0.088576279163805, 
    -0.078826403509137, -0.069763335827687, -0.060324245822426, 
    -0.051185892938683, -0.042214125381494, -0.032400948835467, 
    -0.022988188423553, -0.014014058101985, -0.0048638597006478, 
    0.0046256558100653, 0.013742295342271, 0.023294962021069, 
    0.032720330508369, 0.042021898355547, 0.05088203165226, 
    0.060203048450087, 0.069665449725571, 0.078988556775417, 
    0.087798140805216, 0.097671755058986, 0.10667703328263, 0.1159970221964, 
    0.1252847715677, 0.13499116749544, 0.14411294242172, 0.15345548141953, 
    0.16272291050166, 0.17249572260741, 0.1815774366376, 0.19118185051471, 
    0.20041889061555, 0.20989863078893, 0.21947000581844, 0.22834182842638, 
    0.23776208475593, 0.24709535648647, 0.25671277891623, 0.26628231654442, 
    0.27551649354677, 0.28513345444899, 0.29462910450006, 0.30415075457051, 
    0.31370572013978, 0.32278857565392, 0.33287908178745, 0.34218193837392, 
    0.35119849525839, 0.36146690851047, 0.37091236545882, 0.38063498665605, 
    0.39014819095934, 0.39985506610166, 0.40950527656874, 0.41907424677904, 
    0.42853660652599, 0.43850165781113, 0.44807992639762, 0.45803625006808, 
    0.46718496844961, 0.47735658657823, 0.48731746646371, 0.49684584755908, 
    0.50685385287558, 0.51667563078686, 0.52680123221257, 0.53639110888382, 
    0.54650623539239, 0.55635076206999, 0.56654500237199, 0.57675661191321, 
    0.58638138213509, 0.59672109122408, 0.60651204692191, 0.61687180024984, 
    0.62686013294244, 0.63707322821057, 0.64720064222124, 0.65751234644682, 
    0.66771881804014, 0.67794553960223, 0.68847865363714, 0.69864480177546, 
    0.70915742861777, 0.71980209437891, 0.73012350515175, 0.74050760398326, 
    0.75108673695676, 0.76160768816524, 0.77216071687588, 0.78285479759176, 
    0.79358959719936, 0.804366346552, 0.81512618650599, 0.82597251657662, 
    0.83683197886684, 0.8477668875145, 0.85863844548318, 0.86968323351245, 
    0.88070553753345, 0.89185776388106, 0.90290062492052, 0.91421363648027, 
    0.92544335774449, 0.93675079014193, 0.94811803168971, 0.95952828783617, 
    0.97103543801252, 0.982571593075, 0.99417752984743,
  -0.99419772297155, -0.98264273237332, -0.97110284057718, -0.95965454382531, 
    -0.94823637216955, -0.93687728655459, -0.92564493882185, 
    -0.91430410317323, -0.90313024896467, -0.89204813949288, 
    -0.88089240366922, -0.86991945610992, -0.85887206337298, 
    -0.84792872970024, -0.83704460727391, -0.82617200623076, 
    -0.81534610065339, -0.80461125571712, -0.79377054994592, 
    -0.78312623269581, -0.77246613946802, -0.7617738663794, 
    -0.75122660246385, -0.74083156081953, -0.73015772292516, 
    -0.71969198502948, -0.70945025650333, -0.69882210404675, 
    -0.68860720646588, -0.67811731669917, -0.66799002224517, 
    -0.65765280701515, -0.64746299286013, -0.63736145867912, 
    -0.62703890558709, -0.61693009461238, -0.60670651651542, 
    -0.59691481883278, -0.58649471930706, -0.57658689326532, 
    -0.56655588628441, -0.55659731237233, -0.54669467557265, 
    -0.53686663680255, -0.52676923039155, -0.51691360444142, 
    -0.50743796873966, -0.49703727255497, -0.48746323896586, 
    -0.47765426096315, -0.46793114050465, -0.4581012163143, 
    -0.44843208685514, -0.43878060793072, -0.4289640321575, 
    -0.41922259042545, -0.40964829855254, -0.4000463073142, -0.3904785097783, 
    -0.38053815613746, -0.37132484067147, -0.36140257692699, 
    -0.35199879186425, -0.34235152777256, -0.33293574651018, 
    -0.3233017443962, -0.31400937461681, -0.30428918766806, 
    -0.29497754127986, -0.28531235617883, -0.27598506987742, 
    -0.26664863964442, -0.25663920272524, -0.24765150084616, 
    -0.23820095560625, -0.22887009416798, -0.21959148508367, 
    -0.20992857449259, -0.20060074971608, -0.19091308323387, 
    -0.18193358384579, -0.17270590552702, -0.16309711445629, 
    -0.15358093136764, -0.14435943553081, -0.13519240180661, 
    -0.12580284135404, -0.11621283258506, -0.10742517784518, 
    -0.097897883789307, -0.088138388191328, -0.079325349642448, 
    -0.069808748919702, -0.060695373987705, -0.051103427464667, 
    -0.041931583748723, -0.032152642793774, -0.023405194306392, 
    -0.014031092201002, -0.0047816348042792, 0.0047160992721866, 
    0.013684713033003, 0.023396353852268, 0.032415221699636, 
    0.042202974802958, 0.051222638734245, 0.060028922123315, 
    0.069754388342293, 0.079238105202745, 0.088157913143401, 
    0.097847552899318, 0.1072675766532, 0.11610455414161, 0.12569655472546, 
    0.13520058232863, 0.14450491162843, 0.15372763174419, 0.16284783397435, 
    0.17250963920993, 0.18159125223692, 0.19148121237384, 0.20050777507121, 
    0.21016049095021, 0.21936470100051, 0.228823395109, 0.23828978445745, 
    0.24744443243891, 0.25709390376227, 0.26662188210116, 0.2759022990556, 
    0.28556624730579, 0.29480708462016, 0.30456967512758, 0.31395612492558, 
    0.32329276496356, 0.33326347598545, 0.34268624904613, 0.35219220290182, 
    0.36180194357856, 0.37113344471811, 0.38120718832171, 0.39044404602793, 
    0.40043413556831, 0.40972510432694, 0.41970989764208, 0.42925378522222, 
    0.43892249257114, 0.44873662614939, 0.45842148877597, 0.46807455927703, 
    0.47819857551531, 0.48768295938013, 0.49767508446009, 0.50734274736237, 
    0.51729279855467, 0.52735409813122, 0.53700290204236, 0.54708299037619, 
    0.55694856391684, 0.56699000342907, 0.57703620101968, 0.58725397801415, 
    0.59707194105657, 0.60719871348338, 0.61728749811494, 0.62743646917052, 
    0.63764899689771, 0.64785349639382, 0.65813763883871, 0.66841854056796, 
    0.67872144987979, 0.68882354810291, 0.69918626965175, 0.70978398808797, 
    0.72002560915511, 0.7306865500576, 0.74105471615123, 0.75154226846515, 
    0.76216216930036, 0.77274905080086, 0.78344612402845, 0.79406018902422, 
    0.80472504452426, 0.81561052353014, 0.82630835084622, 0.83715592001192, 
    0.84805971689746, 0.85905331460087, 0.87001219356389, 0.88107176268588, 
    0.89213063385275, 0.90325356407534, 0.91439379676487, 0.92564951588122, 
    0.93694703294269, 0.94828700908031, 0.95966422338794, 0.97109789853578, 
    0.98262934278611, 0.99419818175889,
  -0.99421642496958, -0.98267699808688, -0.9711925246546, -0.95976810057493, 
    -0.94841262475728, -0.93707178400761, -0.92580349254361, 
    -0.91459943328533, -0.90341056667412, -0.89228658514113, 
    -0.88121880235834, -0.87023673969545, -0.85922690183917, 
    -0.84825225119121, -0.83744016777961, -0.82648044224781, 
    -0.81578009966307, -0.80489416882235, -0.79432167075137, 
    -0.78367866701729, -0.77292009964277, -0.7624169502814, 
    -0.75165973902075, -0.74122941248434, -0.73075086714513, 
    -0.72028845907705, -0.70977771675008, -0.69940174483359, 
    -0.68900375715163, -0.67884805672964, -0.66845097689503, 
    -0.65819240969951, -0.64809448776088, -0.63776341181923, 
    -0.62767622262561, -0.61741451614409, -0.60734081165188, 
    -0.59744052977224, -0.58743394910287, -0.5769793868624, 
    -0.56723215156826, -0.55714377952453, -0.54722646880313, 
    -0.53726066268904, -0.5275177066002, -0.51745553406907, 
    -0.50745728639218, -0.49766267607664, -0.48807660639447, 
    -0.47837905779245, -0.46845464503022, -0.45879066412707, 
    -0.44874297557274, -0.43892101944123, -0.42977288748049, 
    -0.41960779614093, -0.41003158980117, -0.4005027929899, 
    -0.39085861783356, -0.38105635597937, -0.37147648087465, 
    -0.36212196703677, -0.35270609981133, -0.34263713496652, 
    -0.33337736934776, -0.32349840260859, -0.31428470485885, 
    -0.30482063944116, -0.29542013347616, -0.28553868710423, 
    -0.27631163724038, -0.26708984383325, -0.25720317141167, 
    -0.24800440414292, -0.23857517759493, -0.22911934018865, 
    -0.21973527085041, -0.20994790411234, -0.20102386920687, 
    -0.19156192748837, -0.18214118460378, -0.17276283660098, 
    -0.16348409430114, -0.15410235587434, -0.14440658606895, 
    -0.13497634122608, -0.12583869737883, -0.11667022191445, 
    -0.10709092697409, -0.098174468975968, -0.088699231444342, 
    -0.079184379277988, -0.07000434746975, -0.060527361028561, 
    -0.051413889827166, -0.041928955296586, -0.032641328955176, 
    -0.023306686391601, -0.014004413870231, -0.0046369801067137, 
    0.0046473789548154, 0.013592568149253, 0.02358666069326, 
    0.032573474215179, 0.041747778812909, 0.050986187381164, 
    0.060491905358201, 0.070096991122873, 0.079023573921517, 
    0.088437690098182, 0.09769760705388, 0.10741254801968, 0.11677616137248, 
    0.12570414462295, 0.13529492164423, 0.14478581977493, 0.15384865373197, 
    0.16321266129427, 0.17270067104143, 0.18215465527731, 0.1915734447879, 
    0.20100493973831, 0.21034949240829, 0.21939769442633, 0.22917867320066, 
    0.23836266422212, 0.24800891512771, 0.25718153911544, 0.26735437043322, 
    0.27616800756132, 0.285775131883, 0.29556583794186, 0.30469900330478, 
    0.31413064851155, 0.32410579573778, 0.33369335183447, 0.34314852658816, 
    0.35257164779278, 0.36223962523308, 0.37194505536479, 0.38137560032748, 
    0.39111152299521, 0.40049116186057, 0.41062958204392, 0.42001968077641, 
    0.42982057201234, 0.43950806559959, 0.44928668355554, 0.45890858494868, 
    0.46870862085588, 0.4785405225696, 0.48816200096827, 0.49816954294128, 
    0.50783501336292, 0.51778890356719, 0.52775056610322, 0.53773895855097, 
    0.54765905659523, 0.55773570077404, 0.56767950587914, 0.57738111214719, 
    0.5878642093098, 0.59781736339719, 0.60763598857895, 0.6179384741455, 
    0.62796323000214, 0.63801229669669, 0.64843650876823, 0.65861941851042, 
    0.66904081289228, 0.67895313344373, 0.68966883925179, 0.69969480086547, 
    0.71027147638849, 0.72063982456496, 0.73106932352779, 0.74151197360634, 
    0.75211441252194, 0.76273606982984, 0.7730491145944, 0.78389026787059, 
    0.79448426642924, 0.80518257477883, 0.81603597569055, 0.8267132837189, 
    0.83755585515874, 0.84844422061573, 0.85937176830804, 0.87028421598998, 
    0.88139017316367, 0.89239753484895, 0.90351244680379, 0.91464470027569, 
    0.92584513549151, 0.93712345328833, 0.94842344847546, 0.95978443043431, 
    0.97120822163406, 0.98267596617302, 0.99421334019315,
  -0.99424931431646, -0.98277598067815, -0.971347811775, -0.95999626043258, 
    -0.94869696794532, -0.93739382086505, -0.92616487626895, 
    -0.91507150922534, -0.90387206602345, -0.89286921225654, 
    -0.88175424428342, -0.87079968863305, -0.85991585177801, 
    -0.8490031535427, -0.8381533392863, -0.82724642178297, -0.81658923088645, 
    -0.8058694310891, -0.79498106476549, -0.78440912805579, 
    -0.77381868038151, -0.76321972902524, -0.7527067682303, 
    -0.74216296671471, -0.73164014224743, -0.72134362523081, 
    -0.71073982824875, -0.70045205842479, -0.69017977639727, 
    -0.67986007460619, -0.66934291145791, -0.65925309169848, 
    -0.64904862795512, -0.63891885302344, -0.62875391485532, 
    -0.61876126659401, -0.60831519621653, -0.59823145834429, 
    -0.58822719867591, -0.57811762974814, -0.5682666355674, -0.558370425808, 
    -0.54839910960353, -0.53839611587806, -0.52865615404632, 
    -0.51855049697431, -0.50863849789026, -0.49887018903215, 
    -0.48896881162779, -0.47888162818409, -0.46919002314488, 
    -0.45949062841517, -0.44995172041338, -0.44013268937665, 
    -0.43049023723005, -0.42061935806867, -0.4109519699175, -0.4014474258136, 
    -0.39174340219456, -0.38221156164341, -0.3726276580818, 
    -0.36289955553962, -0.35303802844342, -0.34376945965115, 
    -0.33424877017296, -0.32449611301569, -0.31534744889593, 
    -0.30503002466658, -0.29578271168097, -0.28639495039337, 
    -0.27679925137779, -0.26772001305369, -0.25788092829155, 
    -0.24876344281308, -0.23923684754712, -0.22994111196672, 
    -0.22031225626241, -0.21080742489877, -0.20114049358518, 
    -0.19185742116578, -0.18229214660345, -0.17346643873959, 
    -0.16382106894757, -0.15422266288726, -0.14503860716955, 
    -0.13576499153773, -0.12642402414314, -0.11680876379808, 
    -0.10714476366239, -0.097768209867257, -0.08899432973517, 
    -0.079742592780115, -0.070177925241469, -0.060388894280756, 
    -0.05161921079014, -0.042014843635409, -0.032731984383266, 
    -0.02342431895954, -0.014317119980273, -0.0047495046013329, 
    0.0046203014061155, 0.014036935128751, 0.023216768873361, 
    0.032971068288317, 0.041802456183631, 0.051035402133244, 
    0.060826671706355, 0.070266179010138, 0.079494741453807, 
    0.088596083749867, 0.098232968312594, 0.10731145157025, 0.11699937051374, 
    0.1260647267345, 0.13567414028055, 0.14488315912344, 0.15429923090248, 
    0.16372856641823, 0.17328211741694, 0.1828000681246, 0.19232475370551, 
    0.20151911263023, 0.21075815010324, 0.22024362881999, 0.22944315238236, 
    0.23909482958608, 0.24859046851031, 0.25799893412361, 0.26756455945489, 
    0.27702878168101, 0.2862777822908, 0.29606796921253, 0.30580919136637, 
    0.31501332557509, 0.32498279489344, 0.33432960128975, 0.34387809955203, 
    0.35351380810594, 0.36304996530772, 0.37273820355343, 0.38212018578515, 
    0.39203133289111, 0.40165942435804, 0.41126160507664, 0.42093587867876, 
    0.43069121432815, 0.4405058584869, 0.45013900729927, 0.46015998769594, 
    0.4696232579892, 0.47959240114619, 0.48913677454977, 0.49932714328634, 
    0.50912483599491, 0.51893268518482, 0.52887017328341, 0.53874702979143, 
    0.54859888360637, 0.5587740856701, 0.56844376449854, 0.57848655063942, 
    0.58871671630347, 0.59870821121239, 0.60894636008398, 0.61891522046214, 
    0.6292466293242, 0.63913582511481, 0.64923474485709, 0.65964282375277, 
    0.66998483670563, 0.68011811590707, 0.69047852235919, 0.70089968146225, 
    0.71122169778669, 0.72166177719997, 0.73198123497634, 0.74259731981591, 
    0.75299352258602, 0.7635584228581, 0.77394059074541, 0.78470847182878, 
    0.79526516660233, 0.806015137033, 0.81676385591864, 0.82748595325286, 
    0.83824685518143, 0.84911705175744, 0.86007016478077, 0.87095203721816, 
    0.88188493125436, 0.89296457708918, 0.90393801680094, 0.91507791814118, 
    0.92624055222682, 0.93746748128738, 0.94869660084625, 0.96000166682271, 
    0.97135955213085, 0.98277958526447, 0.99424930771495,
  -0.99430634197987, -0.98295162000288, -0.97164154646308, -0.9603763679286, 
    -0.94915520558661, -0.93799416520564, -0.92691257072531, 
    -0.91580106204792, -0.90472830876656, -0.89381260923444, 
    -0.88275092431576, -0.87193725556815, -0.86101702560656, 
    -0.85022115475504, -0.83935985743161, -0.82868478594646, 
    -0.81789957464081, -0.80730455667561, -0.79653315295223, 
    -0.78586976807908, -0.77539079951587, -0.76490603357738, 
    -0.75437163697116, -0.74383382729712, -0.73347622624743, 
    -0.72291201017156, -0.71255201939589, -0.70221864632429, 
    -0.6920217097992, -0.68175804287465, -0.67136431720491, 
    -0.66091764503654, -0.65108897331843, -0.64076256746659, 
    -0.63064954207517, -0.62024736934758, -0.61058439652751, 
    -0.6001237725224, -0.59007502448117, -0.5801347399477, -0.57011442431354, 
    -0.56021038798635, -0.5500301059579, -0.54030706479916, 
    -0.53026151080558, -0.52035109429504, -0.51038853515839, 
    -0.50070013248617, -0.49095202177635, -0.48107291822328, 
    -0.47126426597782, -0.46129505601005, -0.45165197912562, 
    -0.44191505929844, -0.43233094696365, -0.42232347523838, 
    -0.41262047549036, -0.40284601359672, -0.39342121087812, 
    -0.38354810113665, -0.37423035268043, -0.36431973848436, 
    -0.35450201209232, -0.34524789549932, -0.33558670633291, 
    -0.3260427351283, -0.31613624232163, -0.30678341625757, -0.2974655245129, 
    -0.28760535238699, -0.27797220472454, -0.26855046365306, 
    -0.25915122003276, -0.24971727500201, -0.24025107103374, 
    -0.2305009368004, -0.22131195489954, -0.21207924931299, 
    -0.20227801156795, -0.19304679406627, -0.18331634360047, 
    -0.17407865640251, -0.16422569373969, -0.15499456613157, 
    -0.14551545217424, -0.13627076872706, -0.12707322113344, 
    -0.11771808386951, -0.10775237805711, -0.098610572924102, 
    -0.089249443745026, -0.079913674498641, -0.07015445982204, 
    -0.061153540949916, -0.051490511455509, -0.042113493050161, 
    -0.032898304666665, -0.023570958896532, -0.014266129203678, 
    -0.0047265532209215, 0.0045504524422807, 0.01445759711161, 
    0.023111897184934, 0.033055582429277, 0.042369053171878, 
    0.051311487533126, 0.061301733717625, 0.070259041673835, 
    0.079593967116836, 0.089264377697746, 0.09850685313927, 0.1079978847908, 
    0.11733670702894, 0.12696638065519, 0.13645164111251, 0.14544667307708, 
    0.15521507045068, 0.16443325081648, 0.1738133012063, 0.1836031342901, 
    0.19309677936805, 0.20225611942098, 0.2118546511741, 0.2211657110985, 
    0.23095847577034, 0.24033450039411, 0.24980494578068, 0.25943860706705, 
    0.26848834086858, 0.27811208514196, 0.28784666291846, 0.29754844300343, 
    0.30705450381164, 0.31654678061825, 0.32607406433797, 0.33583188314667, 
    0.34534619212722, 0.35514750191762, 0.36442586195984, 0.37418737321286, 
    0.38374587254972, 0.39353535466127, 0.40348498537474, 0.41289324699861, 
    0.42253429612127, 0.43255061935433, 0.44207534702114, 0.45205870138032, 
    0.46156031132776, 0.47175853874938, 0.48126184782557, 0.49099849859508, 
    0.50103874106008, 0.51101361694382, 0.52067629006998, 0.5305601751385, 
    0.54071873921472, 0.55065016773471, 0.56036428671948, 0.57044159393232, 
    0.58052046154142, 0.59056344831433, 0.60064968706825, 0.61067107197081, 
    0.62088004947517, 0.63085130009972, 0.64118910393533, 0.65114255608096, 
    0.66152238937978, 0.67177059293592, 0.68183668322635, 0.69237865479621, 
    0.70258918926621, 0.71286816258296, 0.72338989282718, 0.73366271174521, 
    0.74418269202735, 0.75454665486398, 0.76516799569499, 0.77566170590003, 
    0.7861335994355, 0.796891358741, 0.80739607621761, 0.81807869143308, 
    0.82876816071832, 0.83962988111883, 0.85030712266117, 0.86115277980007, 
    0.87202975900925, 0.88289404837164, 0.89383785442936, 0.90482219827481, 
    0.91586480605567, 0.92693154029008, 0.93800918424433, 0.94920640020177, 
    0.96039921483301, 0.97165132351759, 0.9829523261113, 0.99430954611146,
  -0.99436147859516, -0.98309326014785, -0.97188309504717, -0.96071118777791, 
    -0.94965810065917, -0.93842991539483, -0.9274629429066, 
    -0.91655349419729, -0.90546328430936, -0.89449281421528, 
    -0.88363396984465, -0.87296190156888, -0.86199387630175, 
    -0.85121211494371, -0.8403657197855, -0.82974101096279, 
    -0.81901758508118, -0.80865845986484, -0.79780487002505, 
    -0.78743252736147, -0.77678333569564, -0.76618132932959, 
    -0.75556400619882, -0.7452101040881, -0.73516056035895, 
    -0.72476671120587, -0.7141130068722, -0.70370396246786, 
    -0.69367639526603, -0.68325698081773, -0.67284002716742, 
    -0.66297053826952, -0.65213410311896, -0.64243184297046, 
    -0.6325963242213, -0.6221721973227, -0.61203723764068, -0.60187401125718, 
    -0.59180115213336, -0.58178510902209, -0.57175930683802, 
    -0.56228757819371, -0.55155224883191, -0.54141333526097, 
    -0.53181764060178, -0.52149121162657, -0.51228879920643, 
    -0.5023562392617, -0.49245002135755, -0.48237548727082, 
    -0.47274685338191, -0.46284864805042, -0.45310389896329, 
    -0.44346431555298, -0.43377713530918, -0.42413852593964, 
    -0.41424299433465, -0.40426984334792, -0.39424399095994, 
    -0.38455032321542, -0.37513505739172, -0.3656921879995, 
    -0.35642118878459, -0.34665508171002, -0.33667999463894, 
    -0.32678536829296, -0.31718045443065, -0.3077701755891, 
    -0.29864653810034, -0.28882046015865, -0.27902684062604, 
    -0.26963939829358, -0.25929913503742, -0.25058090417206, 
    -0.24108735238729, -0.23224004019907, -0.22284341204786, 
    -0.21286204262361, -0.20300609429039, -0.19371496242784, 
    -0.18374661556822, -0.17502514143461, -0.1654511434631, 
    -0.15615644558763, -0.14610414873291, -0.13661910389254, 
    -0.12748610711208, -0.11809419422728, -0.10879585694361, 
    -0.098590194604498, -0.08963704132022, -0.079337002636273, 
    -0.070508531866368, -0.061484876059518, -0.052549564450715, 
    -0.042156139465707, -0.032984933523671, -0.023083861982779, 
    -0.01362881748123, -0.005003984852613, 0.0041809643630659, 
    0.013369508777692, 0.022887942391359, 0.033219176732831, 
    0.042522712953304, 0.051656798297832, 0.06167454596144, 
    0.071269243625689, 0.079790882706026, 0.089303441409566, 
    0.098133016950736, 0.10822604600969, 0.11828882816627, 0.1276608676031, 
    0.1373040331286, 0.14690265663639, 0.15570491814726, 0.16527887813989, 
    0.17458624460631, 0.1843109213848, 0.19326448101596, 0.20306119516596, 
    0.21243479663251, 0.22236310877508, 0.23230295688093, 0.24159792896134, 
    0.25070417467186, 0.25970515656488, 0.2698585540201, 0.27961654292286, 
    0.28887075077778, 0.29850290032987, 0.30856627772086, 0.31749787345068, 
    0.32690500097511, 0.33649635508842, 0.34637161815573, 0.35681426656836, 
    0.3663046489225, 0.37522402549434, 0.38539504912266, 0.39469094233054, 
    0.40454933949899, 0.41446535123223, 0.42420764522796, 0.4341173924689, 
    0.44353071173853, 0.45290251201805, 0.46314960544581, 0.47257858065213, 
    0.48247975045245, 0.49303196569634, 0.50285388647669, 0.51321710453301, 
    0.52289666903899, 0.53257524973952, 0.54193473650253, 0.5515283278004, 
    0.56168622393412, 0.57239125505411, 0.58231526303819, 0.59202977512188, 
    0.60276730124492, 0.61285095977214, 0.62313729642699, 0.63240312566524, 
    0.64224594204384, 0.65256336609225, 0.66308804950108, 0.67324487817372, 
    0.68316850676878, 0.69375860619489, 0.70456110083942, 0.71443322596272, 
    0.72468656479403, 0.73494590947657, 0.74553882180287, 0.7559122946338, 
    0.76649797941883, 0.77687733041148, 0.78732834050471, 0.79827874130712, 
    0.80880217264332, 0.81909533520407, 0.83010532787814, 0.84065021964052, 
    0.85131764606045, 0.86203977177828, 0.87315058151136, 0.88385663766548, 
    0.89457196613208, 0.90555009967332, 0.91645080872072, 0.92756231963116, 
    0.93845333350425, 0.94957984001517, 0.9607750855043, 0.97196715087634, 
    0.98307678070874, 0.99435517187429,
  -0.99439904926956, -0.98323198994658, -0.97209515657678, -0.96101156428462, 
    -0.94997080780342, -0.93892107121605, -0.9279871847249, 
    -0.91702511430118, -0.90610390602154, -0.89527221836646, 
    -0.88441797072888, -0.87366777119888, -0.86282591824353, 
    -0.85223344534903, -0.84139886924231, -0.8307832777233, 
    -0.82019125187984, -0.80953726988213, -0.7989423564946, 
    -0.78845062967106, -0.77805627757235, -0.76744544381576, 
    -0.75698826652858, -0.74658152530664, -0.73617574838888, 
    -0.72577176097992, -0.71556033961805, -0.70512247640639, 
    -0.69491008383642, -0.68453582155601, -0.6744076387907, 
    -0.66409152399933, -0.65404767883829, -0.64383903709654, 
    -0.63364693585198, -0.62345702355481, -0.61339029940653, 
    -0.60328128337538, -0.59313398348592, -0.5833207520026, 
    -0.57335146802234, -0.56321842479585, -0.55341666230921, 
    -0.5432296525173, -0.53347102617932, -0.52351122699942, 
    -0.51357636756676, -0.50366284676488, -0.49364584028448, 
    -0.48388668189088, -0.47423752323281, -0.46424661812142, 
    -0.45444004596881, -0.44455103708988, -0.43483086251072, 
    -0.42532587318565, -0.41526872330119, -0.40580025052985, 
    -0.39584822817863, -0.38618497353314, -0.37670497355293, 
    -0.36704327654258, -0.35706622213089, -0.34738595367867, 
    -0.33777394393649, -0.32839727495493, -0.31869136470253, 
    -0.30893613049739, -0.29934146378579, -0.28983293745136, 
    -0.28027464103507, -0.27076075873487, -0.26115194109548, 
    -0.25143966086732, -0.24170817137025, -0.23251417523518, 
    -0.22290274005908, -0.21356945293565, -0.20391789268773, 
    -0.19407562466887, -0.1849564965357, -0.17525566932111, 
    -0.16553564588858, -0.15650637747763, -0.14664676093396, 
    -0.1373456667263, -0.12789836288461, -0.11821530050894, 
    -0.10875685558549, -0.099605419349012, -0.089943592333238, 
    -0.080525838326542, -0.070887938001412, -0.061563874711003, 
    -0.051964997497856, -0.04249080931722, -0.033285500375899, 
    -0.023590535491053, -0.014208888050695, -0.0049588711669808, 
    0.0047018712841762, 0.014317665420956, 0.023694097312339, 
    0.033130244569612, 0.042571369095951, 0.051736667768447, 
    0.06145902077397, 0.070944963570238, 0.080545195382347, 
    0.089832810668695, 0.099033079760305, 0.10891448674369, 0.11853458593473, 
    0.12794093896078, 0.13739727148167, 0.14670432685982, 0.15613198711589, 
    0.16601849668103, 0.17538861766104, 0.18482803999778, 0.19418454507634, 
    0.20382357520911, 0.21352790902325, 0.22305108336864, 0.23260701917515, 
    0.24201765135921, 0.2515176227117, 0.26104593025297, 0.27078558678699, 
    0.28024504653586, 0.28983100461037, 0.29965468963198, 0.30923313613453, 
    0.31865849305571, 0.32846309248907, 0.33823756440082, 0.3477226046624, 
    0.3575644663654, 0.36708758821671, 0.37681730719327, 0.38627743608181, 
    0.3961678977535, 0.4059310911135, 0.41546202217855, 0.42549019416427, 
    0.43521294230949, 0.4451280658311, 0.45471836319259, 0.46466946881886, 
    0.47439434794862, 0.48412127963107, 0.4942079959951, 0.50385822395364, 
    0.51408207553442, 0.52364252411123, 0.53344581830509, 0.54378498511918, 
    0.55380844952666, 0.56348096830137, 0.57350512512208, 0.58374035116979, 
    0.59357617906109, 0.60366362147044, 0.61373947847281, 0.62382966106692, 
    0.63402164897336, 0.64421387644094, 0.65415128117623, 0.6645682322027, 
    0.67468869047341, 0.68487099878949, 0.69520325877599, 0.70540290769595, 
    0.71577302027608, 0.72603892400887, 0.73646489225983, 0.74692892793895, 
    0.75721901015814, 0.76766803949615, 0.77808501840461, 0.78866559118745, 
    0.79918821859567, 0.80973799657268, 0.82028121399642, 0.83097745629932, 
    0.84158523652953, 0.85226409436522, 0.86302885929463, 0.87372060790459, 
    0.88451976475151, 0.89533824776534, 0.90618068243834, 0.91709641958207, 
    0.92800496607974, 0.93900441196835, 0.94998061849698, 0.96102783651601, 
    0.97210248501111, 0.98323710832028, 0.99440261149313,
  -0.99445789767919, -0.9833955754781, -0.97237707555025, -0.96138462577007, 
    -0.95042042622952, -0.9395006892548, -0.92860291951417, 
    -0.91775294078273, -0.90693582570261, -0.89615063130276, 
    -0.88537692882692, -0.87466033422771, -0.86399075347689, 
    -0.85329070081302, -0.84265548810334, -0.83198007034898, 
    -0.82155811067215, -0.81096367867164, -0.80036033995601, 
    -0.78981936401849, -0.77954147961392, -0.7689945204773, 
    -0.75857655011288, -0.74818995376657, -0.73784928773484, 
    -0.72755621536939, -0.71708042652907, -0.70691186348548, 
    -0.69656024234319, -0.68627983231969, -0.67614460660175, 
    -0.66625334043402, -0.65568327143163, -0.64542683221991, 
    -0.6355660560936, -0.62544521111351, -0.61527485268056, 
    -0.60504501452774, -0.59522711632238, -0.58516194890756, 
    -0.57512973087157, -0.5649603844319, -0.55523391251726, 
    -0.54503707687388, -0.53540814251631, -0.52522481596165, 
    -0.5154496828455, -0.50541740989651, -0.49552519764037, 
    -0.48575028019272, -0.47582367868972, -0.46604450537023, 
    -0.45623882585119, -0.44654612873175, -0.43646009482788, 
    -0.42664530546893, -0.4170522052861, -0.40740757940172, 
    -0.39747235058388, -0.38801748961656, -0.37816743502045, 
    -0.36832158441541, -0.35879276805525, -0.34898152684862, 
    -0.33936694610736, -0.32933717932601, -0.32024910588746, 
    -0.31025563895243, -0.30064839209842, -0.29118797627523, 
    -0.28176180237005, -0.27183557003054, -0.2620455240192, 
    -0.25267986434171, -0.24291405686408, -0.23355012027905, 
    -0.22410405916006, -0.21411133855532, -0.20457013425604, 
    -0.19514344032946, -0.18561624442478, -0.17609602684689, -0.166557005821, 
    -0.15717666176404, -0.14767708808567, -0.13769836380164, 
    -0.12860298601077, -0.11869499425204, -0.1093041263969, 
    -0.09963368044839, -0.090353899388669, -0.080863477513715, 
    -0.071414057119391, -0.061543523360279, -0.052684780834147, 
    -0.042619325928507, -0.033159761347002, -0.023803614170474, 
    -0.014241752244506, -0.0047009033045126, 0.004758265854377, 
    0.014164722418878, 0.023522191291047, 0.033196084890342, 
    0.042769402198949, 0.052298606001766, 0.06169528691937, 
    0.071464404778275, 0.080795230323709, 0.090389918737446, 
    0.099473431265921, 0.10948922584412, 0.11906340723926, 0.12822768677731, 
    0.13820523886492, 0.14707646155134, 0.15698227433662, 0.16670874623116, 
    0.17587864136947, 0.18562599204192, 0.19534214829448, 0.20490768568128, 
    0.21422102634916, 0.22389423782414, 0.23342900634144, 0.24337536393601, 
    0.2525834984718, 0.26247127087126, 0.27176777084189, 0.28154351957341, 
    0.29135799221083, 0.30085131282626, 0.31048039707906, 0.31992338765344, 
    0.32995428539751, 0.33957224177339, 0.34930524317866, 0.35888958767915, 
    0.36834988560237, 0.37834568256962, 0.38813390996944, 0.39768635592122, 
    0.40755230830563, 0.41722463069847, 0.42710675087597, 0.43695623887475, 
    0.4466831482043, 0.45657460899596, 0.46633579262701, 0.47603470839878, 
    0.48580025068913, 0.49587663604897, 0.50591915518219, 0.51560577875984, 
    0.52566760745431, 0.53545929679673, 0.54538860527873, 0.55547124922926, 
    0.56532505231381, 0.57551598966071, 0.58541924982786, 0.59545288250258, 
    0.60542023125074, 0.61572321060936, 0.62564975318889, 0.63570206148759, 
    0.64588907482181, 0.65613258331492, 0.66627774618677, 0.67650619469948, 
    0.68658381230773, 0.69682363393096, 0.70719474401998, 0.71740787890057, 
    0.7277001594253, 0.73811527588219, 0.74840857519318, 0.75882109475639, 
    0.76926508364896, 0.77968709903157, 0.79003483425966, 0.80055951722945, 
    0.8111176753731, 0.82163241595815, 0.83219776380535, 0.84276764448123, 
    0.85339800067127, 0.86411371849269, 0.87470125510134, 0.88549087238961, 
    0.89621987273609, 0.90697375161093, 0.91784227987949, 0.92863426213329, 
    0.93951709927661, 0.95045715504474, 0.96138263845494, 0.97237954879926, 
    0.98339905660795, 0.9944589251991,
  -0.99447463443406, -0.98343771900447, -0.97246970846643, -0.96148994249118, 
    -0.9504862813677, -0.93969767427837, -0.92879871466352, 
    -0.91796284482383, -0.90719083738494, -0.89644344685067, 
    -0.88561760469727, -0.87491168246505, -0.86431728744369, 
    -0.85355254723212, -0.84304295287152, -0.83253523774241, 
    -0.82189397899793, -0.81117186531766, -0.80082298467281, 
    -0.79029296218653, -0.77987794451532, -0.76951352653632, 
    -0.75914367821334, -0.74849015704982, -0.73834378148739, 
    -0.72827998703053, -0.71767321366027, -0.70712932891626, 
    -0.69713287840009, -0.68689440847467, -0.6766549369697, 
    -0.66665950023949, -0.65628929972404, -0.64609877138886, 
    -0.63590372940018, -0.62578263529155, -0.61549554975348, 
    -0.6059037027088, -0.59600962724744, -0.58595372512721, 
    -0.57552778609528, -0.56561077290992, -0.55558798964008, 
    -0.54558655773009, -0.53575537365909, -0.52574198683008, 
    -0.51576958600733, -0.50596897940158, -0.49646030955422, 
    -0.48609462119251, -0.47644843923097, -0.46666560192457, 
    -0.45669121870457, -0.44711065312542, -0.43702564712687, 
    -0.4272495283222, -0.41773448173656, -0.407872922689, -0.39807964557422, 
    -0.38849284638607, -0.37853181772333, -0.36864516382131, 
    -0.35910431483564, -0.34916117945349, -0.33966703411351, 
    -0.32990074607531, -0.32043707303548, -0.31098509319239, 
    -0.30137229092556, -0.29135416171217, -0.28182596697092, 
    -0.27198896387454, -0.26236625748551, -0.25322476745103, 
    -0.24337688428693, -0.23355154545729, -0.2241199730811, -0.2148642242953, 
    -0.20504039524756, -0.19513059625264, -0.18632352067593, 
    -0.17640458476107, -0.16631576073229, -0.15731439628623, 
    -0.14796809935196, -0.13807156370861, -0.12872887264103, 
    -0.11937283576991, -0.10933076308644, -0.099592215101843, 
    -0.090732964553521, -0.080375680903218, -0.071303592959978, 
    -0.062029453209631, -0.052583723346454, -0.042675211953286, 
    -0.033221154715665, -0.023622860666799, -0.01438753471544, 
    -0.0049437236473273, 0.004859737288195, 0.014414228705433, 
    0.023361101450393, 0.03300757125059, 0.042819746772015, 
    0.052473708712933, 0.062238491688205, 0.071442702208196, 
    0.080716709595509, 0.090569776044454, 0.09958413260582, 0.10959659589578, 
    0.11893481890824, 0.12853885861027, 0.13810787142069, 0.14735860153996, 
    0.15714523661542, 0.16641693734936, 0.17611502781702, 0.1865929338277, 
    0.19524110286009, 0.20475555906831, 0.21424532291302, 0.22476069194699, 
    0.23440786515686, 0.24378930319735, 0.25298096899619, 0.26226813707239, 
    0.27247986216546, 0.28163275668998, 0.29157692859196, 0.30104710951813, 
    0.31102153431203, 0.32079805136903, 0.33016675789595, 0.33974942575581, 
    0.34940825473039, 0.35924794602506, 0.36907824870899, 0.37880766611436, 
    0.38871312425165, 0.39805960275949, 0.40805963123674, 0.41788953417705, 
    0.42714334355706, 0.43762890110246, 0.44738607531732, 0.45704819660284, 
    0.46674544940505, 0.47645279757409, 0.48648489517961, 0.49641616094052, 
    0.5066344785747, 0.51610970251285, 0.52611449186752, 0.53607264653, 
    0.54563589248994, 0.55554958035552, 0.56626358049178, 0.57595171461427, 
    0.5859123175485, 0.59576714993825, 0.60615727377159, 0.61627435286039, 
    0.62641353136943, 0.63638988016217, 0.64646346294068, 0.65656962089879, 
    0.66672816494503, 0.67683685915247, 0.68720498268863, 0.69763913190485, 
    0.70763993929075, 0.71771556694281, 0.7284316145157, 0.73842557617301, 
    0.74889777736508, 0.759448478637, 0.76968670892302, 0.77995258525842, 
    0.79044021373149, 0.80082388795218, 0.81163346389543, 0.82200224523177, 
    0.83271591153174, 0.84315241806556, 0.85364191733068, 0.86425042173238, 
    0.87513605214023, 0.88581281367337, 0.89640203581038, 0.90720705460383, 
    0.91806745628714, 0.92879634982631, 0.9396741175265, 0.95059137983226, 
    0.96149979441197, 0.97246060257781, 0.98345368356487, 0.99447546926949,
  -0.99452960578125, -0.98360889577503, -0.97271523544007, -0.96185941944786, 
    -0.951021701907, -0.94021786716039, -0.92943753588871, -0.9187180942672, 
    -0.9079705244462, -0.8973159705137, -0.8866016194477, -0.87606816146364, 
    -0.86536074205544, -0.85478259739285, -0.844242978942, -0.8336990533491, 
    -0.82330781768825, -0.81266078891249, -0.80226325372263, 
    -0.79192826576508, -0.78142923339584, -0.77102727105034, 
    -0.76065840179957, -0.7503423619468, -0.74007237107233, 
    -0.72977775344116, -0.71947254402069, -0.70910109638361, 
    -0.69888897061828, -0.68877013702827, -0.67850377432435, 
    -0.66834969406754, -0.65818787980231, -0.64822481588849, 
    -0.63809269110217, -0.62764358524463, -0.61785967873455, 
    -0.6076347798788, -0.59761847568273, -0.58749671892924, 
    -0.57769197889808, -0.56766521604056, -0.55765869153973, 
    -0.54763202003226, -0.53762687998534, -0.52768306740508, 
    -0.51787154796537, -0.50802711432871, -0.49799623055155, 
    -0.48790772010766, -0.47822832841374, -0.46830883836088, 
    -0.45872415734236, -0.44876172670249, -0.43879212577425, 
    -0.42924623562334, -0.41921607528875, -0.40944396487346, 
    -0.39965318765404, -0.38991030422658, -0.3802289654319, 
    -0.37046964558971, -0.36053627841958, -0.35089930430752, 
    -0.34147739685728, -0.33141420159936, -0.32170497395366, 
    -0.31250548114988, -0.3024003896871, -0.29279501314327, 
    -0.28285218505533, -0.27362772178807, -0.26385750627166, 
    -0.25424816365544, -0.24429182592743, -0.23504471371816, 
    -0.22503698041807, -0.21563071122452, -0.20602673648462, 
    -0.19615663800786, -0.18698281994979, -0.1771349616864, 
    -0.16777802058348, -0.15776078433333, -0.14850918487775, 
    -0.13894329747176, -0.12934426826596, -0.11941139517841, 
    -0.1099966788228, -0.10056189476464, -0.090564064045371, 
    -0.081429688319104, -0.071788059410548, -0.062174766714661, 
    -0.052568973627041, -0.042944753973538, -0.033450152665878, 
    -0.02381151009257, -0.014518171891813, -0.0050304289307575, 
    0.0046844342529685, 0.014295937141958, 0.023941755936199, 
    0.033360252203402, 0.043234463023584, 0.052782217225736, 
    0.061846534499421, 0.071644653207838, 0.081470224773199, 
    0.091012928117635, 0.10041274625561, 0.10979873205953, 0.11959297926089, 
    0.12923605804717, 0.13864777213861, 0.14832970712179, 0.15808754468775, 
    0.16761169918689, 0.17726924405103, 0.18673367226743, 0.19662098183327, 
    0.20591777069391, 0.21567476708507, 0.22526148279761, 0.23479467814888, 
    0.24448382422614, 0.25422166855743, 0.26391926904482, 0.27360308779347, 
    0.28295496213738, 0.2931392786951, 0.30245506238534, 0.31228287032747, 
    0.32184490947916, 0.33169405665786, 0.34130125826902, 0.35111993679436, 
    0.36075970537855, 0.3706170082528, 0.38030214476628, 0.38992849162951, 
    0.40002792400799, 0.40986465334731, 0.41951957026136, 0.428876785044, 
    0.43910652154132, 0.44895606302514, 0.45869314732007, 0.46878114013047, 
    0.47828219144635, 0.48840031489557, 0.49832213064134, 0.50811829085444, 
    0.51812915142603, 0.52786178619149, 0.53773389378253, 0.54774064610843, 
    0.55787977742542, 0.56795773241662, 0.57784756837928, 0.5878674392421, 
    0.59790581836889, 0.6079018008041, 0.61802439064354, 0.62804831684057, 
    0.63815730548292, 0.6481817655084, 0.65841595614835, 0.66855039061548, 
    0.67890406981023, 0.68893446981688, 0.69919504013269, 0.70935228206988, 
    0.7197277670923, 0.72991567335776, 0.74018833190839, 0.75053597425951, 
    0.76096684105884, 0.77109801137225, 0.78159237235694, 0.79201728505248, 
    0.80238579184951, 0.81288772500463, 0.82333159974706, 0.83386632429616, 
    0.84436922776514, 0.85486129427781, 0.86551599627448, 0.87604276830634, 
    0.88673321521062, 0.89738452199814, 0.90800791788897, 0.91874534084238, 
    0.92947534763746, 0.94024704141133, 0.95104989844161, 0.96186549402941, 
    0.97272182514129, 0.98361213264907, 0.99453281129984,
  -0.99455451351286, -0.98368231296517, -0.97282816834625, -0.9619981053986, 
    -0.9512202590778, -0.94046377556648, -0.92971361367452, 
    -0.91899949660051, -0.90834717590323, -0.89771254723265, 
    -0.88702879986175, -0.87642444898536, -0.86588896674972, 
    -0.85527610087499, -0.84477503799043, -0.83430694246646, 
    -0.82375014426901, -0.81337929705273, -0.80287905866042, 
    -0.79246569419315, -0.78210975066536, -0.77179542163068, 
    -0.76133514983743, -0.75103538291982, -0.74078338726074, 
    -0.73038150760946, -0.72016815176099, -0.70989063924374, 
    -0.69979584175334, -0.68948557798832, -0.67928536201692, 
    -0.66924332468239, -0.65898651400246, -0.64890760427767, 
    -0.6386404385834, -0.62877125658922, -0.61847935479935, 
    -0.60856236925158, -0.59853772331612, -0.58834659311772, 
    -0.57843158492589, -0.56827282184661, -0.55846086515271, 
    -0.54845776938848, -0.53857082248011, -0.52842523531202, 
    -0.51874679637985, -0.50884009489587, -0.49868508886065, 
    -0.48880791612714, -0.47907637599628, -0.46913810964452, 
    -0.45924599958579, -0.44963141102392, -0.43957867713155, 
    -0.42988244389197, -0.419992085452, -0.41021688382216, -0.40030145476471, 
    -0.39054544515616, -0.38087178415081, -0.37124818672594, 
    -0.36139231153116, -0.35158765917757, -0.34202480705229, 
    -0.33239065970573, -0.3221912985502, -0.31279443405834, 
    -0.30302812761889, -0.29326677864213, -0.28374137790792, 
    -0.27399837362688, -0.26431125579974, -0.25457766820598, 
    -0.24494963624592, -0.23538903865935, -0.22573265261358, 
    -0.21611365520151, -0.20629363281318, -0.19690916650524, 
    -0.18717390855571, -0.17759949982516, -0.16776962006999, 
    -0.15831814584327, -0.14859512384183, -0.13924073348782, 
    -0.12917283322036, -0.11997492525366, -0.11033767700292, 
    -0.10076142835627, -0.091218307528523, -0.081548840426013, 
    -0.071822582896568, -0.062213695056727, -0.052653382671737, 
    -0.043270133254296, -0.033592994139049, -0.023930053268477, 
    -0.014273489405191, -0.0049010381634801, 0.0046539053578047, 
    0.014385044956439, 0.024078948783663, 0.033406207129382, 
    0.043185483376191, 0.052564668475081, 0.062485075862679, 
    0.071866598059781, 0.08152745974242, 0.090874038179939, 0.10060109683528, 
    0.11030734211183, 0.11997555764052, 0.12923186158282, 0.1392149470975, 
    0.1488549284968, 0.15825179843189, 0.16793088266197, 0.17749606047168, 
    0.18700400124266, 0.1968395218033, 0.20653902872373, 0.21623606220818, 
    0.2258231767703, 0.23518938014857, 0.24499262885211, 0.25485895713377, 
    0.26451682616115, 0.27406403752957, 0.28354470244406, 0.29341595412259, 
    0.30301028371345, 0.31291602857139, 0.32261413569643, 0.33214466671104, 
    0.3419345010592, 0.35189557482523, 0.36154824423802, 0.37142147051423, 
    0.38087074402248, 0.39074841390897, 0.40051895175998, 0.4104377493737, 
    0.4201290844425, 0.43010412067791, 0.4396873414139, 0.44957540599169, 
    0.45949689099521, 0.46947269840108, 0.47905406024354, 0.48927201746739, 
    0.49884370656692, 0.50892412931944, 0.51873414013155, 0.52882929199708, 
    0.53877455001135, 0.54870347485734, 0.55855060042374, 0.56873663246922, 
    0.57854009283144, 0.58866007003344, 0.59868715114704, 0.60867251436681, 
    0.61885641260621, 0.62878151222084, 0.6390459217128, 0.6490913006171, 
    0.65918682639507, 0.66941912987874, 0.67953471616052, 0.68963269477872, 
    0.69981852479806, 0.71017416902069, 0.72033620569213, 0.73060778486533, 
    0.74097189798657, 0.75118254527723, 0.76158879766302, 0.77183127222974, 
    0.78222632982446, 0.79262983326572, 0.80301193707816, 0.81348419833905, 
    0.82389361310084, 0.83438127148895, 0.84484845938293, 0.85537315003763, 
    0.86593512173228, 0.87651456119994, 0.88709434578163, 0.89773730541039, 
    0.90837178138545, 0.91906685025912, 0.92974782225723, 0.94048492688338, 
    0.95123166724477, 0.96202760877792, 0.97283580374074, 0.98368336413989, 
    0.99455640658608,
  -0.99457498404921, -0.98374253446119, -0.97292445073923, -0.96213666529453, 
    -0.95142394554129, -0.94067183639868, -0.92996686172737, 
    -0.91933114991742, -0.90861534097938, -0.89805678541829, 
    -0.88739427372304, -0.87688895777876, -0.86626895823107, 
    -0.85571813294366, -0.84526535229129, -0.83475243152953, 
    -0.82425080551888, -0.81390535969684, -0.80344221936281, 
    -0.79301924863373, -0.78277818135828, -0.77231415511456, 
    -0.76200648783273, -0.75167956286442, -0.7413780177477, 
    -0.73126761145878, -0.72086864023411, -0.71069379553892, 
    -0.70037959568865, -0.69009797733589, -0.68003124574089, 
    -0.66982892772523, -0.65995504839097, -0.64958490521462, 
    -0.63952663937236, -0.62929235215173, -0.61925421419686, 
    -0.60943345537613, -0.59924339554714, -0.5892977976, -0.57913574415444, 
    -0.56906210582431, -0.55920056276376, -0.54931018355174, 
    -0.53912025495245, -0.52925430731447, -0.51928943908253, 
    -0.50938873036104, -0.49980031014586, -0.48964884524928, 
    -0.4796241470218, -0.46985741467233, -0.45999671090354, 
    -0.45014207272743, -0.44022905556939, -0.43054017343832, 
    -0.42071950890501, -0.41095125176151, -0.40113334518793, 
    -0.39129521537528, -0.38139422083334, -0.37174178675617, 
    -0.3619575932628, -0.35226649706875, -0.3425087019104, -0.33261971237724, 
    -0.32300671848192, -0.31320921737681, -0.30352913386365, 
    -0.29389764423672, -0.2840916101445, -0.27469749951973, -0.26470552316, 
    -0.25506049171962, -0.24536056701111, -0.23573775169639, 
    -0.22614842986286, -0.21630338764659, -0.20676523028233, 
    -0.19722209536767, -0.18753053999067, -0.17792769429667, 
    -0.16817172477193, -0.15836152492517, -0.14912408135451, 
    -0.13934330050526, -0.1299381419647, -0.12003071003094, 
    -0.11022620918878, -0.1007638596174, -0.091397477712906, 
    -0.081673965027087, -0.072028181203816, -0.062679533153892, 
    -0.052708212381724, -0.043349185753553, -0.033732571319795, 
    -0.023826735339745, -0.014290398402215, -0.004757576475607, 
    0.0046978087148598, 0.014415746140079, 0.024309254036235, 0.033265045363, 
    0.043143086120777, 0.05285644987675, 0.062315635694467, 
    0.071953940337774, 0.08160118552353, 0.091532148634819, 0.1009512295049, 
    0.11034344288235, 0.12017124479312, 0.12976830097045, 0.13923037567385, 
    0.14903453485635, 0.15882699844132, 0.16841307487528, 0.17809004034251, 
    0.18740291851085, 0.19710689364743, 0.2065118596593, 0.21631679259402, 
    0.22635967405734, 0.23588056574664, 0.24515317943433, 0.25513944398731, 
    0.26508131814931, 0.27456007187063, 0.28408099851413, 0.29390759658137, 
    0.30381360396509, 0.31329218135459, 0.32312254362377, 0.33301794970312, 
    0.3425870795461, 0.35222861760229, 0.36189687265707, 0.3718969569269, 
    0.38161543675026, 0.39146665842973, 0.40126122633271, 0.41103197312069, 
    0.42068874725745, 0.43055114756859, 0.44036468234924, 0.45035425561515, 
    0.4603347176588, 0.47002442001378, 0.4799851809375, 0.48967984767385, 
    0.49963708462436, 0.50967117773409, 0.51952183346474, 0.52951571768953, 
    0.53948588835333, 0.54931302621819, 0.55924735902734, 0.56930030558263, 
    0.57942656000163, 0.58950362084474, 0.59935303088544, 0.60930225174609, 
    0.61948147541803, 0.6297569163864, 0.63964030745983, 0.64974624856581, 
    0.66004075194565, 0.66992043636144, 0.68028147774895, 0.69044585731232, 
    0.70057725535366, 0.71077417669954, 0.72102952481121, 0.73120959559247, 
    0.74149832613869, 0.75188833894761, 0.76217543905725, 0.77257143286153, 
    0.78268370652831, 0.79321223465446, 0.80358898284098, 0.81391077342201, 
    0.8244027494833, 0.83488048160654, 0.84531970586134, 0.8557948840288, 
    0.86641243131426, 0.87690166616322, 0.88743888801255, 0.89807939317263, 
    0.90868265745267, 0.91931839296785, 0.92999325443932, 0.94070514194873, 
    0.95140839179013, 0.96216986032944, 0.97293901144764, 0.98374208851838, 
    0.99457629102952,
  -0.99458447538467, -0.98377570670719, -0.97296827305685, -0.96218264727051, 
    -0.95146740072793, -0.9408068562361, -0.93018126173055, 
    -0.91930818794432, -0.90883598582182, -0.89829856471433, 
    -0.8876111345279, -0.87696040189505, -0.86623041020403, 
    -0.85600073596476, -0.84566004896667, -0.83505649449923, 
    -0.82433341124468, -0.81444053368703, -0.80374379109339, 
    -0.79294667812858, -0.7827819068993, -0.77238483534087, 
    -0.76225387577065, -0.7523154036806, -0.74181672336098, 
    -0.73172619812253, -0.72131639757712, -0.7107779464387, 
    -0.70075433104726, -0.69048821953588, -0.6801421633043, 
    -0.67036152473104, -0.66037537194094, -0.64997922034136, 
    -0.63987326056837, -0.62971464706218, -0.61948846922454, 
    -0.6095797414513, -0.59947520120705, -0.58958193381434, 
    -0.57941697321204, -0.56980967437758, -0.55982574639897, 
    -0.54970465522377, -0.53947390908776, -0.52918775106638, 
    -0.5197241434846, -0.50934096637172, -0.49995733447559, 
    -0.49066924408216, -0.47998330194305, -0.4699178556018, 
    -0.46012824612038, -0.45078223317737, -0.44084141243222, 
    -0.43111505236308, -0.42089966684484, -0.41081083441822, 
    -0.40098014941901, -0.39151127425004, -0.38224583725011, 
    -0.37230239533481, -0.36236029746301, -0.35234736906458, 
    -0.34259937153161, -0.33267747178277, -0.32295132303617, 
    -0.3136631291509, -0.30411472269193, -0.29440921072742, 
    -0.28489909628074, -0.27444297232588, -0.26469045547225, 
    -0.25465537493945, -0.24523751301155, -0.23631838138564, 
    -0.22657574951878, -0.21685827441545, -0.20716169617602, 
    -0.19730890955488, -0.18686696908541, -0.17761864895145, 
    -0.1687971870021, -0.15915638418749, -0.14887411461727, 
    -0.13905261379173, -0.1298005170771, -0.12010344289143, 
    -0.11047935628395, -0.1010356744822, -0.09150433337277, 
    -0.081805285319023, -0.071762916599249, -0.062568026546156, 
    -0.05280341967643, -0.043584981927262, -0.033894094699488, 
    -0.024332761679733, -0.013761045959436, -0.0051471249815337, 
    0.0050323990041739, 0.014306997789216, 0.023460337659608, 
    0.033235100652951, 0.043928164541773, 0.052621989906725, 
    0.062867263949513, 0.07302045056289, 0.082061836947797, 
    0.091093512078286, 0.10070857106505, 0.10954736309654, 0.12044777722817, 
    0.12979369001427, 0.13938673626046, 0.14883537063114, 0.15883331273442, 
    0.1684007680295, 0.17800421668138, 0.1877349360782, 0.19742082994113, 
    0.20646731004259, 0.21694174943518, 0.22599698317679, 0.2355463914085, 
    0.24552292901153, 0.25574769099568, 0.26555850085716, 0.27484231162821, 
    0.28425552732179, 0.29401739957143, 0.30410531858285, 0.31361335047766, 
    0.32404767657233, 0.33319864264154, 0.34343745402379, 0.35230020910462, 
    0.36205979452472, 0.37203270190312, 0.38165128924418, 0.39148421492082, 
    0.40124307119668, 0.41196700998657, 0.42143307931458, 0.43090893959518, 
    0.44082582911368, 0.45033156195553, 0.46054719602015, 0.47079552904188, 
    0.48021304909177, 0.48974781289535, 0.49970077760597, 0.50983124231819, 
    0.52048424849519, 0.52979336488985, 0.53982906081875, 0.54930549653588, 
    0.55962107616866, 0.56976644343119, 0.57953985474192, 0.58994331229281, 
    0.60000681854082, 0.60969220248884, 0.61993931388395, 0.62928338094101, 
    0.63982311814346, 0.6502140114614, 0.66049969714065, 0.67048000646022, 
    0.68041914648505, 0.6905858139453, 0.70075652656758, 0.71139801697225, 
    0.72138824023574, 0.73170030743648, 0.74182328277634, 0.75179928139856, 
    0.76244237863337, 0.77281269217634, 0.78320905496696, 0.79367395377584, 
    0.80353018504837, 0.81410142246256, 0.82447191588701, 0.83507072175105, 
    0.84573333895831, 0.85593644533064, 0.86664234420962, 0.8770678751775, 
    0.88769890995325, 0.89823364524937, 0.90872058761506, 0.91942561586755, 
    0.93018487393556, 0.94079035828976, 0.95146120391654, 0.96222967311185, 
    0.97300248808473, 0.98378297742914, 0.99458466083269,
  -0.9946105761352, -0.98384963430977, -0.97311894884911, -0.96239795468308, 
    -0.95171012411064, -0.94103726332746, -0.93041334942145, 
    -0.91976867636833, -0.90919960722866, -0.89860568906562, 
    -0.8880681488201, -0.87752496307334, -0.86705294897207, 
    -0.85653065965505, -0.84606770715343, -0.83567557111181, 
    -0.82520430884751, -0.81480130179076, -0.80447517126888, 
    -0.79401399149173, -0.78378799768529, -0.77331179237359, 
    -0.76319363078268, -0.75287659717659, -0.74247321609991, 
    -0.73223261875974, -0.72206664475815, -0.71191049382382, 
    -0.70159102340445, -0.69145888785729, -0.68131659420719, 
    -0.67120064613804, -0.66093439708658, -0.65089832912606, 
    -0.64078124619117, -0.63078232675115, -0.62052879497333, 
    -0.61063501009779, -0.60054199569783, -0.59054251751088, 
    -0.58061778700175, -0.57034975387952, -0.56057525152576, 
    -0.55057232172015, -0.54043719935125, -0.53048283604075, 
    -0.52074796923366, -0.51054986669217, -0.5009343223802, 
    -0.49083052289753, -0.4811078097357, -0.4710478518515, -0.46119404724834, 
    -0.45157066033586, -0.44157254698337, -0.43169391201349, 
    -0.42185748736755, -0.41205605746918, -0.40218584651515, 
    -0.39225172552493, -0.3827763772826, -0.37290258746969, 
    -0.36313415229613, -0.35340087242053, -0.34336595172965, 
    -0.33355352190115, -0.32391043076645, -0.31432425752579, 
    -0.30455504048651, -0.29485634379958, -0.28494019865697, 
    -0.27536605748618, -0.26559849638593, -0.25603993038519, 
    -0.24614892021957, -0.2364340778205, -0.22671280260312, 
    -0.21729293177603, -0.20738937687548, -0.19768728626738, 
    -0.18808256227557, -0.17852347685187, -0.16881994654392, 
    -0.15916970911794, -0.14926041374596, -0.13974612406452, 
    -0.1301317528641, -0.12056611183428, -0.11091067179835, 
    -0.10106322614202, -0.091665999703822, -0.081867445229998, 
    -0.072354551608579, -0.062451693132287, -0.052998717825438, 
    -0.043485443969047, -0.03372559826771, -0.023866699372138, 
    -0.014450708594861, -0.0046441975714963, 0.0047623887974062, 
    0.014415834086454, 0.024212902037009, 0.033634991841378, 
    0.043421195119473, 0.052972570526477, 0.062663412781951, 
    0.071973394741824, 0.081984430561053, 0.091635405379215, 0.101177355224, 
    0.11087673226288, 0.12058145611802, 0.13007015559284, 0.1399211745846, 
    0.14940345446859, 0.15911804619713, 0.16858093410544, 0.178720465582, 
    0.18823263299606, 0.19781103149528, 0.20741480766375, 0.21706481377905, 
    0.2268208379662, 0.23660432715022, 0.24629124201814, 0.25581106616597, 
    0.26575888457796, 0.27561584965841, 0.28501605700851, 0.29482882898273, 
    0.30453511612466, 0.314295157788, 0.32424922050193, 0.33382621200122, 
    0.34343837569084, 0.35329536130345, 0.36318980557271, 0.37293202412017, 
    0.38280688718941, 0.39237280635028, 0.40228959137181, 0.41200426681239, 
    0.42208120839644, 0.43188370444195, 0.44168106792677, 0.45137889935873, 
    0.46140318893072, 0.47121365713576, 0.48115598393662, 0.49096702220761, 
    0.50091306816755, 0.51078091020913, 0.52089955351777, 0.53066866149071, 
    0.54064220311513, 0.55065989359881, 0.56059991636443, 0.57068314080531, 
    0.58061902639512, 0.59071030788969, 0.60055381360435, 0.61067519682419, 
    0.62077393285712, 0.63081233383122, 0.64100233881643, 0.65095840768646, 
    0.66117139874534, 0.67125948201171, 0.68143486184418, 0.69155956757315, 
    0.7017365237072, 0.71200920801511, 0.72213686880061, 0.73238090738168, 
    0.74267933140147, 0.75289679641947, 0.7631555443398, 0.77350938139931, 
    0.78381564066444, 0.79413333986556, 0.80455664779399, 0.81490377990576, 
    0.82524533998858, 0.83572632100922, 0.84609803431682, 0.85661628496047, 
    0.86709971092123, 0.87755830977029, 0.88813322693742, 0.89864987725327, 
    0.90919040494315, 0.91981962086756, 0.93041861276448, 0.94105057428264, 
    0.95172330180396, 0.96240502128534, 0.97311683479431, 0.98385308916177, 
    0.99461475082506,
  -0.99462751354075, -0.98389455902745, -0.97319460207098, -0.96251117242599, 
    -0.95184131755388, -0.94120398989051, -0.93056400991061, 
    -0.92002445483771, -0.90942329873333, -0.89887747836207, 
    -0.88831782347852, -0.87786920701954, -0.86735731624156, 
    -0.85693004589218, -0.84639667280453, -0.83598300762014, 
    -0.82567571342095, -0.81523747015856, -0.80487674875851, 
    -0.79453310761589, -0.78411388359585, -0.77393198124264, 
    -0.7636283459078, -0.75326414433443, -0.74308093623235, 
    -0.73279607980637, -0.72258857934687, -0.71237640641331, 
    -0.70230695457831, -0.6919461019001, -0.68187087890678, 
    -0.67172570685958, -0.66158046333211, -0.65150685863961, 
    -0.64134076392983, -0.63133131806899, -0.62115031627664, 
    -0.61119640807261, -0.60111393678455, -0.59115709849548, 
    -0.58112357828728, -0.57101730474619, -0.56104275730412, 
    -0.55100243014191, -0.54122263331665, -0.53114435959003, 
    -0.52130664992856, -0.51121420634022, -0.50139900337622, 
    -0.49134619685382, -0.48154904776738, -0.47183548541449, 
    -0.46165785884157, -0.45205250852928, -0.44206459256694, 
    -0.43229065479913, -0.42236034377361, -0.41255331056288, 
    -0.40268578236907, -0.39295794142869, -0.38301293928038, 
    -0.37315245938103, -0.36364320486271, -0.35379363911668, 
    -0.34396176781864, -0.33440177450873, -0.32420808414271, 
    -0.31456835060606, -0.3049793360503, -0.29507356250157, 
    -0.28517967870599, -0.27586007588424, -0.26617958029793, 
    -0.25640112306782, -0.24656882450469, -0.23688775285367, 
    -0.2270611937515, -0.21732945045422, -0.20767673145147, 
    -0.19815258640501, -0.18833738949703, -0.17858917812225, 
    -0.16904555333322, -0.15940052002226, -0.14963099590492, 
    -0.13991311969813, -0.13057342162895, -0.12052025027542, 
    -0.11097936133883, -0.10123748494955, -0.091735042268223, 
    -0.082083689818324, -0.072266300204522, -0.062594028902759, 
    -0.053102436439266, -0.043472904689758, -0.033758447909117, 
    -0.024184025575797, -0.014488062072569, -0.0048126616126913, 
    0.0048765472610116, 0.014684779768193, 0.024149286260626, 
    0.033829820226883, 0.043290714377886, 0.053021946891683, 
    0.062858108084925, 0.072268365286128, 0.08210221097194, 
    0.091430432357104, 0.10144195038116, 0.11123868761117, 0.12052112456543, 
    0.13041640919841, 0.13986237684919, 0.14975741636874, 0.15941576070798, 
    0.16920994332644, 0.17880493162203, 0.1883624759653, 0.19822583330265, 
    0.20752442283105, 0.21731193096512, 0.22728280607165, 0.23673990908135, 
    0.24676413109956, 0.25626887164537, 0.26610599259483, 0.27588561948767, 
    0.28560192838653, 0.29528534341001, 0.30464494169239, 0.31485962587846, 
    0.32434279298673, 0.33445138673094, 0.34392117527792, 0.35384309299228, 
    0.36370790088961, 0.37315022451189, 0.38329127010479, 0.39277001424096, 
    0.40292583408922, 0.41247727717043, 0.42255116070791, 0.43220276570277, 
    0.44235787930991, 0.45198462374323, 0.46186159360929, 0.47164285252844, 
    0.48167642153869, 0.491678192483, 0.50144057787405, 0.51131386417394, 
    0.52145389872857, 0.53134856644976, 0.54103370788956, 0.55123366100676, 
    0.56114854501599, 0.57117318637859, 0.58131732905401, 0.59128103942297, 
    0.6011577800037, 0.61129881496675, 0.62122839589347, 0.63137590448126, 
    0.64147323217957, 0.65156738849436, 0.66172102242741, 0.67184102084042, 
    0.68201081830513, 0.69210019000354, 0.70218985145368, 0.71248389165857, 
    0.72260227316728, 0.73294434691455, 0.74314506810519, 0.7533942558701, 
    0.76362215540393, 0.77395249108995, 0.78429425437086, 0.79453195315338, 
    0.80495762309886, 0.81524460720214, 0.82568470827429, 0.83610525889713, 
    0.84647671620629, 0.85694721612007, 0.86740339226967, 0.8778825485601, 
    0.88839455434752, 0.89889332405486, 0.90946005158928, 0.91999249188814, 
    0.93059160773571, 0.94124092965955, 0.9518498604153, 0.96251455248019, 
    0.97319572162579, 0.9839028828287, 0.99462675785017,
  -0.99469092635842, -0.98408920743749, -0.9735009466213, -0.96292987112019, 
    -0.95238186419643, -0.94183246937722, -0.93137403557665, 
    -0.92084893635198, -0.91032650851478, -0.89992503851444, 
    -0.88950645776352, -0.87911233400868, -0.8685548011744, 
    -0.85842636064651, -0.84795635899322, -0.83749142551477, 
    -0.82713277141515, -0.81683098282413, -0.80681238138587, 
    -0.79643074831245, -0.7859597565006, -0.77572197715394, 
    -0.76546071956773, -0.75511780902235, -0.74510921941585, 
    -0.73479712753155, -0.72476617185124, -0.71443781639875, 
    -0.70432996883537, -0.69430426695113, -0.68420879942254, 
    -0.67411261364618, -0.66384975247807, -0.6535989014755, 
    -0.64363267976369, -0.63372409577576, -0.62349134558992, 
    -0.61342263079764, -0.6033902421022, -0.59339465656055, 
    -0.58362511427892, -0.57317323876854, -0.56330658661396, 
    -0.55376158992706, -0.54358298283527, -0.53372995259811, 
    -0.52366833437824, -0.51326449695486, -0.50362154755688, 
    -0.49407901983075, -0.48362124038237, -0.47363592993655, 
    -0.46399291403421, -0.45399634976179, -0.44416546058545, 
    -0.4345552894268, -0.4243133182612, -0.41439896333976, -0.40460458057753, 
    -0.3950049552969, -0.38511686162397, -0.37550786126842, 
    -0.36552073767501, -0.35586776585298, -0.34580668561997, 
    -0.33587345412359, -0.32627372576258, -0.31592215945308, 
    -0.30659319693459, -0.29699647939988, -0.28731510475092, 
    -0.27693001822582, -0.26754013460597, -0.25752310256149, 
    -0.2479060305883, -0.23784266484479, -0.2285642266184, -0.21878307439752, 
    -0.20892723132277, -0.19921484407767, -0.18960526864557, 
    -0.17951322100211, -0.16995232501437, -0.16058972893387, 
    -0.15034569956014, -0.14077649758772, -0.13124356800131, 
    -0.12154728338863, -0.11161464018268, -0.10197503651613, 
    -0.091722153020422, -0.082511927023184, -0.073139501453696, 
    -0.062678699466092, -0.053416153134404, -0.043707497899784, 
    -0.034026128436198, -0.02406950832317, -0.014635944109401, 
    -0.0051907629946582, 0.0049629152539146, 0.014579569890734, 
    0.024352629458038, 0.034082216863869, 0.043424163593307, 
    0.053799440652784, 0.06296532641886, 0.072798496799094, 
    0.082447442388533, 0.092124994200256, 0.10178333698757, 0.11187950550036, 
    0.12139424648475, 0.13119492774726, 0.14113976229258, 0.15068470255501, 
    0.16036297684325, 0.17039068075883, 0.17947145148048, 0.18973098151478, 
    0.19942017713591, 0.20899169508221, 0.21834962486085, 0.2285315913887, 
    0.23835881476234, 0.24781242926122, 0.25787035397957, 0.26755587776702, 
    0.2772980071775, 0.28717293345997, 0.29682929866431, 0.30631745821991, 
    0.31651010910147, 0.32602064398483, 0.33616769920942, 0.34607257759395, 
    0.35554455611384, 0.36529213580254, 0.37528097699826, 0.38546280316543, 
    0.39482430213156, 0.40452251706875, 0.41449955336019, 0.42464529689147, 
    0.43440403727538, 0.44417174712138, 0.45421210887418, 0.46382360153559, 
    0.4739504904175, 0.4839639281522, 0.49360884835337, 0.50363387159299, 
    0.51381592862228, 0.52348584915925, 0.53352427884654, 0.54347759605786, 
    0.553436157701, 0.56331752797077, 0.57350520794927, 0.58348298386121, 
    0.59342812849216, 0.60329354085265, 0.61361025401764, 0.62337929396299, 
    0.63356208807355, 0.64358229176357, 0.65377066586027, 0.66392165732424, 
    0.67382714209238, 0.68416641460464, 0.69427093429711, 0.70415199235768, 
    0.71454492112019, 0.72473657774497, 0.73498343965599, 0.74505085832868, 
    0.75525620442676, 0.76551506438444, 0.77581726489745, 0.78596880422871, 
    0.79636057969503, 0.80648384000231, 0.81704532121335, 0.82712978429415, 
    0.8374905601967, 0.84796247713375, 0.85832182509902, 0.86860330626787, 
    0.87907787063202, 0.88940576185085, 0.90006218388474, 0.91028050276959, 
    0.92084895706685, 0.93137445936652, 0.94185392400516, 0.9523782362907, 
    0.96291861722157, 0.97352475626005, 0.98409076813265, 0.99469074992061,
  -0.99473512060186, -0.98421751253281, -0.97371692329485, -0.96323321203323, 
    -0.95276430715864, -0.94230932977902, -0.93187440957577, 
    -0.9214349933336, -0.9110471782001, -0.90065457713777, -0.89025043465387, 
    -0.87994115527928, -0.86956694168316, -0.85925868941899, 
    -0.84889189570779, -0.83860207495195, -0.82835840270852, 
    -0.81804031420838, -0.80781656026021, -0.79751749190167, 
    -0.78734066914584, -0.77710112241876, -0.76683142149649, 
    -0.7567319837443, -0.74649989484086, -0.73636983302484, 
    -0.72611371331452, -0.71594107504871, -0.70599775147351, 
    -0.69569375562272, -0.68561787165407, -0.67560572320973, 
    -0.66539123407979, -0.65538613726496, -0.64523691202604, 
    -0.63521359184232, -0.62517852827972, -0.61509711680657, 
    -0.6052484633265, -0.59510231608592, -0.58493486148257, 
    -0.57506684691117, -0.56506046039639, -0.55517846448755, 
    -0.54509077407742, -0.53505640247196, -0.52508737983819, 
    -0.51538937761555, -0.50520440068364, -0.49530219438732, 
    -0.48544364551061, -0.47542402378522, -0.46569888378356, 
    -0.45563300935691, -0.44566523464217, -0.43594558330166, 
    -0.42593258614543, -0.41611638580936, -0.40612685630182, 
    -0.39643046079154, -0.38641790223236, -0.37661216335639, 
    -0.36675316328476, -0.35673790205947, -0.34727151667795, 
    -0.33733754339302, -0.32738711592068, -0.31763798263929, 
    -0.30770328519054, -0.29794462069304, -0.288076425326, -0.27833453272108, 
    -0.26847448325138, -0.25878534149655, -0.24896483602101, 
    -0.2391132251219, -0.22936405157964, -0.21949653654276, 
    -0.20983210377773, -0.19989343921621, -0.19026685269261, 
    -0.18028119466708, -0.17067400460923, -0.16097932330649, 
    -0.15112903179127, -0.14139648634156, -0.13164365933829, 
    -0.12175280841665, -0.11222775065498, -0.10226757751652, 
    -0.092720207740553, -0.082757623577485, -0.073136039350143, 
    -0.063345145435632, -0.053386185688507, -0.04388047388398, 
    -0.03411486335646, -0.024276486324513, -0.014656826289238, 
    -0.0050700623519281, 0.0049485547913363, 0.014675714391013, 
    0.024533752779094, 0.034180722775662, 0.043995753126284, 
    0.053689428778789, 0.063415514994279, 0.073032547176514, 
    0.082939330308453, 0.092732604903494, 0.10212654237223, 0.11211184777779, 
    0.12203653931434, 0.13155997944061, 0.14164351614261, 0.15111493849726, 
    0.16092882465898, 0.17066672636632, 0.18046600434902, 0.19044001335112, 
    0.19994362567939, 0.20979541509498, 0.2195929670124, 0.22930616496614, 
    0.23914161868248, 0.24890198558142, 0.25887980961401, 0.26848056446884, 
    0.27846315128522, 0.28799953935566, 0.29795289344712, 0.30768417919036, 
    0.31754185859428, 0.3274850455544, 0.33723813287694, 0.3471272972117, 
    0.35679928869297, 0.36684870701711, 0.37645897599898, 0.38652570509073, 
    0.39629080640485, 0.40623866639538, 0.41601585269813, 0.42581255421508, 
    0.43595464725713, 0.44560021293108, 0.45559177288262, 0.46541476676523, 
    0.47562149101909, 0.48537701699133, 0.49524223459822, 0.50518375372051, 
    0.51508647211949, 0.52519539070313, 0.53505776740833, 0.54499149476035, 
    0.55496426971128, 0.56495327173643, 0.57507227391427, 0.58504312340457, 
    0.59505026130562, 0.60505001363245, 0.61503211536972, 0.62510756059281, 
    0.63516981727114, 0.64517519823373, 0.65530979867434, 0.66537044220303, 
    0.67547835097873, 0.68555418683794, 0.69578371236691, 0.70577235111827, 
    0.71596590490794, 0.7261456409957, 0.73623289731886, 0.74640054986091, 
    0.75672500658593, 0.76680939186532, 0.77706454498894, 0.78728101470189, 
    0.79752580231018, 0.80775909676235, 0.81804156693441, 0.8282847578922, 
    0.8385957452459, 0.84887918191897, 0.85924660950319, 0.86953564276158, 
    0.87990580388492, 0.89024646383178, 0.90064790931514, 0.91103859285909, 
    0.92143579725695, 0.93186474825126, 0.94230609562977, 0.95275732543638, 
    0.96323003934846, 0.97371890198666, 0.98421894884424, 0.99473633156981,
  -0.99476876826366, -0.98431548745676, -0.97387786385562, -0.96345114965064, 
    -0.95303297117925, -0.94264207722404, -0.93225542685973, 
    -0.92189698106669, -0.9115393873315, -0.90118070642116, 
    -0.89088853432902, -0.88053295671888, -0.87025427203751, 
    -0.85994746710375, -0.84969976249759, -0.8393990918776, -0.8291661137896, 
    -0.81891911229731, -0.80869044614113, -0.79844937349009, 
    -0.78829180502173, -0.77808647114775, -0.76790453972345, 
    -0.7577166916476, -0.74745980284065, -0.73749261131965, 
    -0.72721514754756, -0.71708733656063, -0.70707133115509, 
    -0.69680161496042, -0.68685438340755, -0.67671087579873, 
    -0.6666448975222, -0.65657530574338, -0.64649545627937, -0.63638522105, 
    -0.62642425897562, -0.61634343712554, -0.60635074122582, 
    -0.59625049619596, -0.58636429778843, -0.57622679994488, 
    -0.56627576283153, -0.5563017230952, -0.5462730451251, -0.5363949149924, 
    -0.52643202718039, -0.51637270644769, -0.50648265641338, 
    -0.49653084601181, -0.48660133738151, -0.47649432578707, 
    -0.46681873240269, -0.45672447455714, -0.4469570082422, 
    -0.43693148753748, -0.4271649652895, -0.4172314782942, -0.40735410598552, 
    -0.3973179055689, -0.3875655045276, -0.37750967619972, -0.36778877602432, 
    -0.35793758686469, -0.34811086828266, -0.3381823678708, 
    -0.32833623484682, -0.31853432766321, -0.30855877597365, 
    -0.29878233005728, -0.28890835990816, -0.27925139119017, 
    -0.26924507939448, -0.25951640191347, -0.24956275846963, 
    -0.24001363850995, -0.2299535376287, -0.22015624596711, 
    -0.21046400013053, -0.2007258728261, -0.19073396919472, 
    -0.18098917128351, -0.17125433359538, -0.1613046137821, 
    -0.15162907895956, -0.14174853936116, -0.13207297007701, 
    -0.12231830202925, -0.11244972358896, -0.10268519914205, 
    -0.092762771352443, -0.083122825051886, -0.073381121147759, 
    -0.063511247915251, -0.053610769848571, -0.04394923106372, 
    -0.034369377195802, -0.024435388468419, -0.014606272338042, 
    -0.0047539894821064, 0.0047482965900173, 0.014644762504942, 
    0.024563929893025, 0.034226166539545, 0.044004570743725, 
    0.053646589471321, 0.063563617583275, 0.073348293593391, 
    0.083104949350445, 0.093029216783111, 0.10259395329605, 0.11249962133352, 
    0.12235308856536, 0.13205698045839, 0.14187830769312, 0.15160561609548, 
    0.16120990350236, 0.171246849593, 0.18105178348519, 0.19074080204635, 
    0.20058335399463, 0.21035261039883, 0.22036188000447, 0.22996610129041, 
    0.2397421774369, 0.24966849542351, 0.25949757146741, 0.26924636998749, 
    0.27903089891692, 0.28900941287689, 0.29874405263371, 0.30854278925677, 
    0.3183096805742, 0.32844890359849, 0.33807764405415, 0.34792708263813, 
    0.35780261728415, 0.36783617168911, 0.37749455684309, 0.38745257682084, 
    0.39746409861099, 0.40708624017164, 0.41708540971088, 0.42699392399184, 
    0.43702997609982, 0.44669435652022, 0.45661578386291, 0.46660116341346, 
    0.47660532394003, 0.48641768539398, 0.49643662892918, 0.50643179561634, 
    0.51627258103735, 0.52628309073082, 0.53619840652281, 0.54614290563947, 
    0.55623922320147, 0.56625131586308, 0.57619100726247, 0.58618157174621, 
    0.59619706465889, 0.60626229352947, 0.61615822086788, 0.6263133519218, 
    0.63637952588663, 0.64640709682225, 0.65642613011052, 0.66652322633247, 
    0.67666162078027, 0.68671112966867, 0.69677248025424, 0.70695070028188, 
    0.71703955114655, 0.72721164756776, 0.7373168506974, 0.74755132460287, 
    0.75760127183179, 0.76782288301306, 0.77804333134012, 0.78820601625115, 
    0.79846052548327, 0.80866381418095, 0.8188543234004, 0.82911066338471, 
    0.83939571494184, 0.8496426462767, 0.85998084610242, 0.87022172374674, 
    0.88054210693732, 0.89083511844801, 0.90120107883747, 0.9115183325964, 
    0.92189567920081, 0.93227160390469, 0.94263877389819, 0.9530473142911, 
    0.96344910565013, 0.97387575835141, 0.98431588422019, 0.99476792325594,
  -0.99479598262382, -0.98439186940278, -0.97399493261641, -0.96364140304449, 
    -0.95331522469188, -0.94287093048416, -0.93256613105337, 
    -0.92218056173158, -0.91197375271097, -0.90155386578388, 
    -0.89135127134142, -0.88098353781024, -0.87082060269764, 
    -0.86076866651722, -0.85013986339417, -0.83993265073726, 
    -0.8298219268206, -0.81948556244229, -0.80930019016394, 
    -0.79917809874372, -0.78908400073793, -0.77910494376384, 
    -0.76867751239245, -0.75847748583392, -0.74812504899009, 
    -0.7381480423976, -0.72812267346783, -0.71793263902884, 
    -0.70794005927982, -0.6980084860901, -0.68773696456683, 
    -0.67759215739967, -0.66744727818441, -0.65728262505675, 
    -0.64695668095526, -0.6376703473862, -0.62763422358536, -0.6176649866311, 
    -0.60722621960636, -0.59729698435029, -0.5870629664549, 
    -0.57714648976924, -0.56701935481604, -0.55759205628954, 
    -0.54742769016452, -0.53760188367358, -0.52697022336095, 
    -0.51752717556932, -0.50757797364322, -0.49748875179484, 
    -0.48723743078734, -0.47731373077316, -0.46751429689835, 
    -0.45769284521219, -0.44814923548036, -0.43772473296219, 
    -0.42795797122614, -0.41775339406122, -0.40790999941767, 
    -0.39859888402232, -0.38832266498577, -0.37872418767606, 
    -0.36876625599155, -0.35845303445027, -0.34822615207755, 
    -0.3393204008665, -0.32920558460447, -0.31932449309772, 
    -0.30921690350509, -0.29942652188567, -0.28961828862072, 
    -0.27941386737044, -0.27007903778696, -0.26027491480148, 
    -0.2498262662113, -0.24049028847568, -0.23031796727678, 
    -0.22064306842425, -0.21127676351476, -0.20143565636557, 
    -0.19101002166707, -0.18142859796567, -0.17118955714343, 
    -0.16157127377343, -0.15197586464912, -0.14274396028338, 
    -0.13246032053667, -0.12257528013649, -0.11234545406437, 
    -0.10235063754066, -0.093078043754877, -0.08364644251133, 
    -0.074117633220154, -0.064081617631207, -0.054197946122042, 
    -0.043836530016882, -0.034269952239421, -0.024148273062856, 
    -0.01462965071551, -0.0048792797280057, 0.0047861899274601, 
    0.014780213968061, 0.024355654484508, 0.034235430520428, 
    0.044170428470207, 0.054067139641607, 0.064006897692807, 
    0.073154460600507, 0.083093725750373, 0.093164465663429, 
    0.10242592284138, 0.11285064962484, 0.12290963381789, 0.13199132002375, 
    0.14171824112591, 0.15180451244621, 0.16193885970001, 0.1720505769209, 
    0.18120928038096, 0.19102162141853, 0.20128851569272, 0.21080833682448, 
    0.22062916887461, 0.23055566047934, 0.24031843465615, 0.25033519251306, 
    0.25982142039604, 0.26988261031196, 0.27980425443389, 0.28944210046542, 
    0.29922286842595, 0.3096415802008, 0.31895581073727, 0.32848906942036, 
    0.33882617567, 0.34862436590891, 0.35812869027966, 0.3688468308294, 
    0.37824112355797, 0.38819000033096, 0.39804434496742, 0.40806023449368, 
    0.41806913710327, 0.42800917435732, 0.43802663421674, 0.44785245158406, 
    0.45762870689437, 0.46711883351853, 0.47743624909378, 0.48744885893761, 
    0.49682322862452, 0.50746638654448, 0.5172669492442, 0.52699655450283, 
    0.53750774629761, 0.54716100740153, 0.55735235449891, 0.56674808808742, 
    0.57690594118051, 0.58681073356556, 0.59724934475666, 0.6076753896039, 
    0.61746510221303, 0.62729436167203, 0.63691036671814, 0.64695458996876, 
    0.65711856528211, 0.6675053578672, 0.67745175544789, 0.68805988099185, 
    0.69797876402868, 0.70776923038763, 0.71785912745745, 0.72785081228534, 
    0.73808032217303, 0.7482922930742, 0.75821027295971, 0.76861825390442, 
    0.77899410556813, 0.78903674866442, 0.79914225860776, 0.80912888935751, 
    0.81931518153176, 0.82989962697063, 0.84031716488264, 0.85014482509877, 
    0.86030317466967, 0.87069907064913, 0.88108942785, 0.89141459535684, 
    0.90148131398204, 0.91196826524743, 0.9221634488731, 0.93262749906194, 
    0.94292689161608, 0.95326275829241, 0.96360786792956, 0.97400809039498, 
    0.98438830804078, 0.99479413446585,
  -0.99481539476866, -0.984453467515, -0.97410545700448, -0.96376717541333, 
    -0.9534417665889, -0.9431193293308, -0.93281685391816, -0.92251761032303, 
    -0.91222848706661, -0.90195041558882, -0.89171839782984, 
    -0.88143534551293, -0.87120629472449, -0.86098890001966, 
    -0.85071625859011, -0.84053912598641, -0.83037468104101, 
    -0.82009998210587, -0.809967326549, -0.79975091042257, -0.7896455090535, 
    -0.77943231572053, -0.76931703259544, -0.75915791343805, 
    -0.74904162200505, -0.73890668656437, -0.72881729742396, 
    -0.71865552598358, -0.70862281621269, -0.698460968725, -0.68847244899948, 
    -0.67837865857897, -0.66828014129033, -0.65816146910509, 
    -0.64819468633497, -0.63815631070994, -0.62806961702488, 
    -0.61806912564703, -0.60807646354393, -0.5979689854046, 
    -0.58796134417746, -0.5780600816709, -0.56800959275759, 
    -0.55808170289444, -0.54804741261338, -0.53801471163815, 
    -0.52802358746089, -0.51809953881806, -0.5081362070278, 
    -0.49820781540722, -0.48826002802202, -0.47828212268334, 
    -0.46836962619743, -0.45835891645004, -0.44853382605027, 
    -0.43859013844825, -0.42866924601513, -0.41867907619542, 
    -0.40880754660187, -0.39886532833984, -0.38898670128674, 
    -0.37915774583845, -0.36908238183539, -0.35928958861576, 
    -0.34948860000779, -0.33958655433367, -0.32959757424625, 
    -0.31971954419902, -0.30994111000252, -0.30003833558139, 
    -0.29012879194414, -0.28025356425013, -0.27041139998564, 
    -0.26055647204814, -0.25083840140334, -0.24085617358505, 
    -0.23104489048446, -0.2211767907564, -0.21130984516508, 
    -0.20155518975138, -0.19162047531731, -0.18187464099276, 
    -0.17195359875677, -0.16201903310608, -0.1523964905342, 
    -0.14225779425026, -0.13272362276122, -0.12291330602452, 
    -0.11295520540957, -0.10305397688607, -0.093236468262237, 
    -0.083624609734114, -0.073574713706473, -0.063899904272252, 
    -0.054014485216111, -0.044138499483049, -0.034513247636585, 
    -0.024553201970004, -0.014685776092655, -0.0050681673984137, 
    0.0048675167203559, 0.014828985239833, 0.024331152876121, 
    0.034447519983365, 0.044124177850805, 0.053999143463851, 
    0.063709538483557, 0.073581552078832, 0.083535522840581, 
    0.093173580886807, 0.1032033323696, 0.11280392329752, 0.12268530180951, 
    0.13262443444143, 0.14233683583567, 0.15237272874445, 0.16200028651891, 
    0.17184192493625, 0.1815368869116, 0.19161640513998, 0.20142179336526, 
    0.21122725381173, 0.22100945320628, 0.23086844363685, 0.24088415941745, 
    0.25056012230299, 0.26046166599729, 0.27033286842397, 0.28007082680185, 
    0.29018666354208, 0.29994515874872, 0.30974190829057, 0.31961113178144, 
    0.32942913872128, 0.33941326668405, 0.349273181116, 0.35912994519465, 
    0.36906277675596, 0.37892232572965, 0.38892194396347, 0.39866091650599, 
    0.40870008676477, 0.41856658701944, 0.42843752469589, 0.43848171728287, 
    0.44829383661231, 0.45823978145053, 0.46812474589593, 0.47814542621183, 
    0.4880399107709, 0.49801810743097, 0.50806439405361, 0.51792152322168, 
    0.52784787839772, 0.53788158013296, 0.5478647936261, 0.55785755543564, 
    0.56785842352264, 0.57783879119671, 0.5878554912592, 0.59785111674793, 
    0.60790019132553, 0.61795896977369, 0.62789562884044, 0.63797174556992, 
    0.64800272942679, 0.65809853924111, 0.66812789806928, 0.67826847444713, 
    0.68831560380887, 0.69836520239287, 0.70848600691215, 0.71860704975269, 
    0.72869645934722, 0.738784359813, 0.74897679105704, 0.75910398650232, 
    0.76920155922331, 0.77938629972308, 0.78954197835294, 0.79969325469291, 
    0.80990635768261, 0.82007454092775, 0.83026799550065, 0.84050050321533, 
    0.85070191571075, 0.86095415567635, 0.87116084765719, 0.88142788257943, 
    0.89167922918918, 0.90194515333353, 0.91222307105524, 0.92250983522346, 
    0.93279961468984, 0.94311404749876, 0.95343030147334, 0.96376349890174, 
    0.97410246022672, 0.98445455159026, 0.99481513868677 ;

 alpha =
  0.94195441308895, 0.8912235988041, 0.85769716219964, 0.82877634869549, 
    0.80246037175108, 0.77744040054658, 0.75176573729612, 0.73428500593946, 
    0.71992869283302, 0.70285142043492, 0.68484349517288, 0.66612383475999, 
    0.64917648785851, 0.63367460959231, 0.61946309796364, 0.60175614708102, 
    0.58908729772107, 0.57622502932073, 0.56162985620631, 0.54521469138437, 
    0.53381614265002, 0.51822093902309, 0.50841477321566, 0.49762157213528, 
    0.48571494728655, 0.47656385080381, 0.46447548235123, 0.45169821212411, 
    0.44015139490439, 0.42913122833793, 0.41490533230739, 0.40226541434342, 
    0.39056953167031, 0.38180592209905, 0.36634834264059, 0.35833536996177, 
    0.34785469909939, 0.33934327744965, 0.32912162322336, 0.31993110577429, 
    0.30947161626283, 0.30030939134654, 0.29330685617601, 0.27994895838948, 
    0.27397192920687, 0.26376934543045, 0.25247862402982, 0.24335307306076, 
    0.23650232093532, 0.22646774915947, 0.2209090856225, 0.21148426708444, 
    0.20270349175863, 0.19732138357503, 0.18645498044729, 0.18121285114406, 
    0.17138295012222, 0.16452226618348, 0.15577872867468, 0.15091144671662, 
    0.14325996664625, 0.13695326281733, 0.13107597161799, 0.12311064312162, 
    0.1176151020175, 0.11183552369394, 0.10334088706977, 0.097782524692833, 
    0.092206756490468, 0.088339081136087, 0.08162014858039, 0.07754474608176, 
    0.072117408147238, 0.067361562546303, 0.061688884779009, 
    0.057411771221266, 0.052678287753141, 0.048812630827792, 
    0.044702250687332, 0.04071274647943, 0.03638952362988, 0.033067220269872, 
    0.029507853111923, 0.026330386003588, 0.023443323517307, 
    0.020623798143854, 0.018374943228259, 0.016564466367349, 
    0.013139705302423, 0.011717982015915, 0.0090739605131293, 
    0.007317664766833, 0.0054203519838957, 0.0041364802435113, 
    0.0029855720148419, 0.0019210936541214, 0.0013599915300892, 
    0.00065936834684549, 0.00027081761926095, 0.00014281983789054, 
    2.5501686417858e-06, 0.0001335279420248, 0.00060098759745357, 
    0.00087916143035995, 0.0015789502743379, 0.0023187588810699, 
    0.003595249546695, 0.0049848524213758, 0.0062255904281196, 
    0.007643966648257, 0.0096587581570991, 0.01142724354083, 
    0.013654920922939, 0.015983772714607, 0.019062795466457, 
    0.021846424190017, 0.025226088908656, 0.027348668907127, 
    0.031543595666465, 0.035046141123906, 0.038161892839298, 
    0.042962162915112, 0.04704501175878, 0.050925522186992, 
    0.057229026379377, 0.062026023719332, 0.065556070884545, 
    0.069092006406984, 0.075749130995997, 0.082713599770704, 
    0.085441245241851, 0.092655464424019, 0.097848285194601, 
    0.10084475756958, 0.10697287870702, 0.11533678373415, 0.12114695891193, 
    0.12923156716223, 0.13535250173864, 0.14007585781116, 0.14739476969566, 
    0.15187661172062, 0.16226736772862, 0.16996435920716, 0.17670374297507, 
    0.18394882122922, 0.19229936158365, 0.1981379438932, 0.21115941919899, 
    0.21528496778808, 0.22728130276065, 0.23718569545067, 0.24485304190955, 
    0.25153483354235, 0.26316624125973, 0.26822462426964, 0.27857249795682, 
    0.28734446404056, 0.30305108951354, 0.30912209685846, 0.3189588683647, 
    0.33010336800903, 0.33865441539985, 0.34751713882251, 0.36147358277584, 
    0.37273689935379, 0.38240294212218, 0.3939806206846, 0.40272989637556, 
    0.41616325374678, 0.42638895785398, 0.43915907640997, 0.44787066563961, 
    0.45947538299784, 0.47206214751194, 0.48534910517202, 0.49945655669226, 
    0.51223182599757, 0.52252873959096, 0.53214691225532, 0.55046196890945, 
    0.56330882813386, 0.57756610415366, 0.58997435506576, 0.60553350152345, 
    0.62066469507055, 0.63678393782657, 0.64981265479303, 0.66723360454719, 
    0.68572903121053, 0.70099323691237, 0.72046543781335, 0.7387394618946, 
    0.75130942264139, 0.77483707434749, 0.794937531571, 0.82776806916157, 
    0.85618157485264, 0.88969318992959, 0.94399168668066,
  0.97943908745933, 0.95074254086926, 0.92839545656601, 0.90739489760613, 
    0.89035298081012, 0.87229111072011, 0.85671829694803, 0.84178519398772, 
    0.82635663973134, 0.81093104790105, 0.79703340928385, 0.78155975935244, 
    0.76866546861975, 0.75580260443486, 0.74237599679307, 0.72968530000359, 
    0.71537706908596, 0.70564332737296, 0.69028237142268, 0.67872239475734, 
    0.66698900581836, 0.65436868002035, 0.64248187014893, 0.62987629131486, 
    0.61849247123857, 0.6078849124856, 0.59393515090492, 0.58487280710845, 
    0.57101400792172, 0.55919113940978, 0.54678852761319, 0.53396992605326, 
    0.52454585158788, 0.5124513800612, 0.49954657844075, 0.48731941626665, 
    0.47877727097497, 0.46602520929964, 0.45357902180662, 0.44355311524133, 
    0.43074644087363, 0.41918662804787, 0.40805783250641, 0.3980536473437, 
    0.38789627506948, 0.37632201617599, 0.36626489450767, 0.35474346695212, 
    0.34264740346806, 0.33353637966825, 0.32407590654797, 0.31206192548638, 
    0.30149384213587, 0.29036203422836, 0.28072137966676, 0.26958114144386, 
    0.26022097113717, 0.25052925370182, 0.24096333062522, 0.23173050668673, 
    0.22111288738361, 0.21019281689813, 0.20094976067792, 0.19201519960417, 
    0.18319853291139, 0.17249242631124, 0.16005074516254, 0.15664103425436, 
    0.14532140879351, 0.13690591637793, 0.12873172969782, 0.12080860655666, 
    0.11370317738619, 0.10793919184227, 0.098750978665107, 0.091192147362782, 
    0.085971554083718, 0.079816485659105, 0.072127400738318, 
    0.065934272049139, 0.059898473878358, 0.053099883617924, 
    0.049177310619978, 0.042557087554042, 0.039071196371352, 
    0.034036032754088, 0.029605846758106, 0.025369632524447, 
    0.021879476633589, 0.018680185423684, 0.014928915491535, 
    0.012567749845112, 0.0095480649953898, 0.0072568410221632, 
    0.005559667017303, 0.0033046599013513, 0.0023026304873163, 
    0.0012414963319779, 0.00048626563133276, 6.7549589857968e-05, 
    1.0989883267052e-05, 0.00021807720589111, 0.00055653822517714, 
    0.001635172786507, 0.002686345832305, 0.0042897301065713, 
    0.0063081865459722, 0.0082043349016712, 0.011041765124365, 
    0.013862270797102, 0.017555588320333, 0.020013206671308, 
    0.023410331633441, 0.02679715379183, 0.031289802516901, 
    0.036348120910583, 0.040883524624225, 0.047670410471142, 0.0524405046808, 
    0.058921798233212, 0.064516047184387, 0.071652766244012, 
    0.077385473348574, 0.083103928437873, 0.091031054518102, 
    0.09839236719717, 0.10615370944919, 0.11420634018848, 0.12072277488576, 
    0.12795122376751, 0.13565799042504, 0.14624983462043, 0.15494555520066, 
    0.16144944918466, 0.17040799771102, 0.17726493888379, 0.1869776720333, 
    0.19858128201691, 0.20810327709012, 0.21692007940096, 0.22470169825054, 
    0.23724349091774, 0.24843566212022, 0.25561804049459, 0.26576447798492, 
    0.27636593868771, 0.28792779103085, 0.29671530492436, 0.30808125829188, 
    0.32047253973796, 0.33170628260698, 0.34259279645856, 0.35248602390604, 
    0.36258543374326, 0.37284909386804, 0.38442495363304, 0.39519581591073, 
    0.40547071339777, 0.41601636850228, 0.43005513721049, 0.44012874603241, 
    0.45000053443008, 0.46094489789671, 0.47233667257922, 0.48445313279332, 
    0.49899287662674, 0.51168874738581, 0.52397726920662, 0.53432679231199, 
    0.5473276434247, 0.55700463157799, 0.56889816295099, 0.58263588847359, 
    0.59265098760052, 0.6059596523357, 0.61761164620546, 0.63036140362724, 
    0.64013881557334, 0.65489557532102, 0.66522459667585, 0.68001068898494, 
    0.69195085753636, 0.7052845280302, 0.7154633128217, 0.72792758996119, 
    0.74221215173172, 0.75568154436623, 0.76848216181265, 0.78280287089648, 
    0.79612209278583, 0.81086597822275, 0.82571915633538, 0.84042385122234, 
    0.85578595564629, 0.87209702548863, 0.88649336586099, 0.90678513151019, 
    0.92770664523111, 0.95056592323693, 0.97926589439077,
  0.99040717517716, 0.97384847455979, 0.95886026546621, 0.94473384881914, 
    0.93154362833745, 0.91871143253411, 0.90658486934121, 0.89472902290218, 
    0.88316823969293, 0.87162542237259, 0.8599547669105, 0.84870644965986, 
    0.83700919281671, 0.82524452871168, 0.81424674534255, 0.8033449416378, 
    0.79268993270279, 0.78113730586237, 0.77092843485293, 0.75975651492902, 
    0.74834618452196, 0.73778912617403, 0.72737175400742, 0.71661168437585, 
    0.70539718054737, 0.6944264240949, 0.68423690806716, 0.67420263152516, 
    0.66164812687067, 0.65138521561693, 0.64010835767076, 0.62878902134739, 
    0.61636831328409, 0.60600541437952, 0.59497520810976, 0.58383228453575, 
    0.57047912421806, 0.55990498250094, 0.54967514489499, 0.53707623706869, 
    0.52531612149459, 0.51467140134326, 0.50231062877813, 0.4910134528168, 
    0.47936067117967, 0.46638647891603, 0.45500859324021, 0.44498502599015, 
    0.4323307611444, 0.42083305088022, 0.4079648459035, 0.39578957271628, 
    0.38323384828653, 0.37229776062579, 0.36232232174947, 0.34973900693342, 
    0.33694342320181, 0.32428240564961, 0.31422978655262, 0.30034663724867, 
    0.29036559967288, 0.27702749115294, 0.26581869398444, 0.25668246880379, 
    0.24554426342577, 0.23382473955461, 0.2206523691645, 0.21078849100072, 
    0.19758573758318, 0.18876261425072, 0.17737559673818, 0.16825750403548, 
    0.15714078558948, 0.14798407458333, 0.13731884639827, 0.12855776037428, 
    0.11896146715894, 0.10972079648386, 0.10191830326303, 0.092112291704843, 
    0.08570638569647, 0.07650956298659, 0.068210433012264, 0.062293525508378, 
    0.055881513155605, 0.048038494748639, 0.042828532972795, 
    0.036433498610989, 0.03106974800888, 0.026168050922678, 
    0.021432231869599, 0.017872991724814, 0.013325229673063, 
    0.010349376894484, 0.0079271954145349, 0.0051056554882046, 
    0.00324044042344, 0.0018490635212454, 0.00065055514933001, 
    7.7600013232e-05, 1.6321682481712e-05, 0.00043370858760566, 
    0.0013173897104553, 0.0026237800605261, 0.0042160970630017, 
    0.006389282207362, 0.0089689920660163, 0.012265190539956, 
    0.016388594152662, 0.020256496857686, 0.024059900449334, 
    0.029463473435591, 0.034140810421562, 0.039959628454923, 
    0.045674754577435, 0.052129617074341, 0.060310893981769, 
    0.067439653144307, 0.074461670090775, 0.083302000968878, 
    0.090410808515019, 0.098613304213677, 0.10747085016743, 0.11539258662306, 
    0.12530251964731, 0.13659720387755, 0.14531663644965, 0.15392518346227, 
    0.16332977807307, 0.173264903236, 0.18496209681608, 0.19748708067766, 
    0.2063150470774, 0.21900525956937, 0.23048904003328, 0.24014991380915, 
    0.25414565245394, 0.26515776485502, 0.27672512080733, 0.28769625387585, 
    0.2994056253248, 0.31060495504381, 0.32230776605977, 0.33368119391392, 
    0.34676730915794, 0.35841702400829, 0.37156088188304, 0.38333943337256, 
    0.39545105773677, 0.40843484645935, 0.42038463761087, 0.43214518719187, 
    0.44316577763721, 0.45614338205902, 0.46594225045649, 0.47871952037644, 
    0.48943144372379, 0.50207684440766, 0.51189015522002, 0.52499989704381, 
    0.53691426900937, 0.54670676843899, 0.55885021890824, 0.56977323910087, 
    0.58268410437801, 0.59448795535339, 0.60594204278978, 0.61598076062504, 
    0.62881029727663, 0.63878627892214, 0.65077707938071, 0.66146494698388, 
    0.67235119332272, 0.68301015622629, 0.69266777390693, 0.7041572785786, 
    0.71595439327041, 0.72672711529714, 0.73795819954038, 0.74903897837855, 
    0.76020871206718, 0.77051000241042, 0.78187103417172, 0.79272065022579, 
    0.8031741956519, 0.81392926110609, 0.82446898557577, 0.83609686277084, 
    0.84725801749509, 0.85848359330061, 0.87003273598379, 0.88204727535934, 
    0.89371174747534, 0.90586073387707, 0.91779414830834, 0.9309199674478, 
    0.94424663509014, 0.95874684065868, 0.97355670069284, 0.99041215988346,
  0.99436425591938, 0.98368881487758, 0.97316746477717, 0.96296232430699, 
    0.95294059930763, 0.94360775021582, 0.93408359756903, 0.92474823989375, 
    0.91547213692663, 0.90650177687499, 0.89694586519343, 0.8878503745531, 
    0.87861860542433, 0.86924543372599, 0.8597865438524, 0.85046874137555, 
    0.84094940292897, 0.83242211594966, 0.82273543242427, 0.8134550398599, 
    0.80436796763397, 0.79455460299558, 0.7857129580972, 0.77572714657041, 
    0.76674836043386, 0.75626054645803, 0.74687938016776, 0.73723347593899, 
    0.72624250821699, 0.71747445166696, 0.70625251411695, 0.69575285730699, 
    0.68605694349796, 0.67408601728928, 0.66420834930002, 0.65423782484289, 
    0.64202068956726, 0.63331084076019, 0.62164162751172, 0.61078110239279, 
    0.60005528910529, 0.58726879680069, 0.57621864529655, 0.5639123894213, 
    0.55136030719143, 0.54096089472212, 0.52932928187709, 0.51663468431925, 
    0.50558183137764, 0.49372986912408, 0.4800399640877, 0.46891568790658, 
    0.45500337313406, 0.4425315712353, 0.43074163678676, 0.4171663283125, 
    0.40440336192396, 0.3903436182594, 0.37859049612188, 0.36503624909215, 
    0.35388958886427, 0.33867977332714, 0.32751162925786, 0.31175492133345, 
    0.30093209587185, 0.2877114588985, 0.27427691430442, 0.26261090110606, 
    0.25059897678211, 0.2364218405401, 0.22368848253544, 0.21071242994679, 
    0.19954975987675, 0.18697279007278, 0.17591586619061, 0.16465343731047, 
    0.15186589886099, 0.14161899852806, 0.13175387945151, 0.12021378072832, 
    0.10978893337063, 0.099140873322759, 0.089173811872823, 
    0.079405871582335, 0.071679798806779, 0.063648090422589, 
    0.055637568250918, 0.047110388423063, 0.040885830646514, 
    0.033988712457871, 0.028417836418778, 0.022776682599804, 
    0.017940404015489, 0.014004872775548, 0.0095784706040396, 
    0.007042418073128, 0.0039337141620506, 0.0023903643079923, 
    0.00092040293414124, 0.00014841300187594, 2.7606527102254e-05, 
    0.00058172145017622, 0.0019028535864964, 0.0033095781672174, 
    0.0060344806443129, 0.0084000319265425, 0.013046093741936, 
    0.016811458228225, 0.020849667336289, 0.027184678344496, 
    0.032459521575237, 0.040213099735131, 0.045004975838564, 
    0.053640638150022, 0.06181590214393, 0.069305421630971, 0.07834910399267, 
    0.087321586840576, 0.095976717400332, 0.10710865402279, 0.11790060105703, 
    0.12681938834423, 0.1381103307044, 0.14850357536248, 0.16138962030485, 
    0.17100956954856, 0.18310991735309, 0.19627849602982, 0.20826858627663, 
    0.22212016955375, 0.23479141483977, 0.24410813882063, 0.25831369857501, 
    0.27287504618783, 0.28533979490185, 0.29641035646499, 0.30990619062075, 
    0.32177469194379, 0.33423654864177, 0.34809725586854, 0.3627860879296, 
    0.37656682785142, 0.38917467894034, 0.40193433190886, 0.4135364193391, 
    0.42846091133314, 0.43992648796868, 0.45317233143602, 0.46478104724676, 
    0.47885202522671, 0.49181216009654, 0.50499311312407, 0.51500043747507, 
    0.52789662233236, 0.53951914368312, 0.55208831930912, 0.56406254498802, 
    0.57480548936645, 0.58565215425525, 0.5980037539066, 0.60887873902349, 
    0.62054671779684, 0.63229137399177, 0.64161336305031, 0.65297745657258, 
    0.66378303581941, 0.6741061617853, 0.68558091047296, 0.69518259870016, 
    0.70561082092265, 0.7159097357388, 0.72633391744152, 0.73685391368367, 
    0.74672724498549, 0.75612852402014, 0.7664257999312, 0.7754320603984, 
    0.78510307863078, 0.79442743801328, 0.80411295866475, 0.81246819755092, 
    0.82276034706812, 0.8316918122308, 0.84186675587337, 0.85071716835061, 
    0.8596727990409, 0.86878029711861, 0.8779492187528, 0.88706627959499, 
    0.89572913134328, 0.905127654533, 0.91467956816482, 0.92399485097377, 
    0.93348672644508, 0.94311843731206, 0.95279124601896, 0.96272769194206, 
    0.97276963955034, 0.9834672925179, 0.99434791217827,
  0.9962159341973, 0.98860463888137, 0.98089277141944, 0.97319465675762, 
    0.96559788234228, 0.9582010689882, 0.95069224127825, 0.94313770292084, 
    0.93544712297776, 0.92820740527588, 0.92047493870803, 0.91274075428912, 
    0.9046585119688, 0.89736716685839, 0.88988227457498, 0.88165112199684, 
    0.87380411039231, 0.86548876606453, 0.85730287197207, 0.85017217875342, 
    0.84231394537551, 0.83390395706478, 0.82514173445959, 0.81656287611549, 
    0.80831624841078, 0.79987291502027, 0.79026430841021, 0.78150181088536, 
    0.77251285709304, 0.76288835802958, 0.75435691712239, 0.74409112550595, 
    0.7352022545518, 0.7253247398147, 0.71671900127811, 0.70595651233357, 
    0.69629121678146, 0.68551871314144, 0.67366254759839, 0.66406133073927, 
    0.65426242123794, 0.64258607769289, 0.63469055832594, 0.62246015011335, 
    0.60910431504865, 0.59812137103405, 0.58698609552871, 0.57553430220487, 
    0.56511637715626, 0.55290024393827, 0.53940143961895, 0.52516031171594, 
    0.51270429547966, 0.49970786951789, 0.48846345025128, 0.47601867650952, 
    0.46209488447155, 0.44804724760458, 0.43422681053937, 0.42088747797683, 
    0.40730011160265, 0.3935651696864, 0.37946702700495, 0.36686491685071, 
    0.34997090723859, 0.33687063053385, 0.3223790016369, 0.31002422497317, 
    0.29458907447795, 0.28190500431983, 0.26891239973641, 0.25381136035968, 
    0.23863534345618, 0.22595771626048, 0.21172821200881, 0.1987475603828, 
    0.18628491148707, 0.17333811871756, 0.15759993209082, 0.14719256617816, 
    0.13334438882582, 0.12166186715055, 0.11048507785422, 0.1001591238354, 
    0.088123537766072, 0.077992081684805, 0.068222089844679, 
    0.058358826637098, 0.050827568267845, 0.042249109945647, 
    0.035329432643867, 0.028109071385324, 0.022727614961546, 
    0.016548380439445, 0.012118202260824, 0.008041152647725, 
    0.0050614710399178, 0.0028844952321092, 0.0011265597238475, 
    0.00019326612654024, 2.7602770903472e-05, 0.00068695206589238, 
    0.0020728472180884, 0.0042117649562697, 0.0077114237650604, 
    0.010881440767846, 0.014947670734085, 0.02101212002037, 
    0.025754534787779, 0.033088164289316, 0.039762157648355, 
    0.048386369170836, 0.056521501424868, 0.066561665610855, 
    0.075072883474586, 0.085870189932235, 0.097174982187383, 
    0.10777633458405, 0.11812378750999, 0.13087750221778, 0.14258810424765, 
    0.15453254344782, 0.17054691265132, 0.18068548436493, 0.19307996936963, 
    0.20769442036181, 0.22129660516041, 0.23436813371539, 0.24752049906093, 
    0.26434719148034, 0.27779191553293, 0.29286656365457, 0.30636689424102, 
    0.3228011054306, 0.33556759198127, 0.34807219265221, 0.36389037898326, 
    0.37746848999497, 0.39200044205314, 0.40547948730275, 0.41464934692249, 
    0.4324974909999, 0.44671927939199, 0.45857702039396, 0.47302886241223, 
    0.48662577031883, 0.49770420240098, 0.51373194052424, 0.52554362220407, 
    0.53792315485284, 0.54840151882379, 0.56208468258745, 0.57526263662315, 
    0.58808696332832, 0.59855874357677, 0.60938104871727, 0.62095362196973, 
    0.63141377248197, 0.64306220043627, 0.65444727386663, 0.66555030012088, 
    0.67642433407481, 0.68695954518384, 0.6962426005875, 0.70631722986234, 
    0.71720690780776, 0.726470744556, 0.73591094646396, 0.74556095567603, 
    0.75546156063126, 0.76601764319725, 0.77257213932335, 0.78200655250617, 
    0.79153435458105, 0.80020943357078, 0.80911000539308, 0.81641702083836, 
    0.82554608862827, 0.83313257556344, 0.84206584298429, 0.85007389858261, 
    0.85862469027989, 0.86632500159008, 0.87380826130746, 0.88185030566143, 
    0.8896343708564, 0.89748971574779, 0.90496851284243, 0.91235807369474, 
    0.9203513999934, 0.92769042571456, 0.93520416426904, 0.94296522824161, 
    0.95017363477191, 0.95768579715058, 0.96534297695168, 0.97303512152194, 
    0.98078475513143, 0.98854537540612, 0.99619823749139,
  0.99717553720749, 0.99139275892645, 0.98570339746122, 0.97959038447131, 
    0.97334307615437, 0.96750905355371, 0.961171660163, 0.9550383519463, 
    0.94886458535162, 0.9426544543528, 0.93606423640333, 0.92972834253205, 
    0.92324009758543, 0.91701960663092, 0.91026568764793, 0.90339146369024, 
    0.89687340217636, 0.88994560250217, 0.88317426849222, 0.87580827545021, 
    0.86877385838746, 0.86174358899047, 0.85500314631197, 0.8465798147946, 
    0.83944611492358, 0.83240956363656, 0.82292106148337, 0.81589740964407, 
    0.80696252892211, 0.79881115412403, 0.79003983207393, 0.78179626688836, 
    0.77476038809433, 0.76460830889086, 0.75676756042696, 0.74698192930786, 
    0.7371548994137, 0.72806790763631, 0.71893946069359, 0.7088791785387, 
    0.69939088828626, 0.69084361434497, 0.67838879188006, 0.66773196509423, 
    0.65632777030015, 0.64595369809865, 0.63341245372657, 0.62222070504042, 
    0.6117579379294, 0.60063839279268, 0.58772251173061, 0.5752050637798, 
    0.56484861532885, 0.55205232220923, 0.53576149558327, 0.52532971876578, 
    0.51195905100415, 0.49965157458438, 0.48282679510824, 0.4696124691917, 
    0.45672604319205, 0.44300202771463, 0.42553309632132, 0.41271310355054, 
    0.39841223998893, 0.38213933806203, 0.370340961634, 0.35127302104323, 
    0.33770805798514, 0.31950318382209, 0.30520718032299, 0.28976093572261, 
    0.27487019802551, 0.25982478473383, 0.24527229257892, 0.2302666610974, 
    0.21469245851967, 0.201353224596, 0.18770891976029, 0.171404885753, 
    0.15868053129159, 0.14481890053518, 0.12998156275358, 0.11683006256324, 
    0.10420907371091, 0.091757719054526, 0.08108525439779, 0.070450852803516, 
    0.06132607164001, 0.05051570173642, 0.042719430820306, 0.0337546289103, 
    0.027489810770584, 0.020913367310111, 0.014671142591351, 
    0.010319692017286, 0.0067872829841346, 0.0031185136788522, 
    0.0011033312622934, 0.00026963124598539, 2.7253902759244e-05, 
    0.00088123243524682, 0.0025339170315707, 0.0051146324867955, 
    0.009006032612033, 0.013770874977539, 0.018955070786418, 
    0.025470031136986, 0.032499236552512, 0.040793096114531, 
    0.048534842554317, 0.057712997998078, 0.067669339929102, 
    0.079424692426903, 0.090076759201285, 0.1033760128348, 0.11401392921398, 
    0.1273028527598, 0.14059125271867, 0.15502835069875, 0.16846841579749, 
    0.18305590160114, 0.20005052915016, 0.21323210406875, 0.22942406297665, 
    0.24386287801214, 0.25746095054387, 0.27413217258238, 0.28692081537921, 
    0.30441545842973, 0.32045242086416, 0.33397571318054, 0.35160603794492, 
    0.36645079339767, 0.38102990475889, 0.39579444157635, 0.40940421148908, 
    0.42427304184653, 0.44014785935004, 0.45394467971796, 0.46516279091042, 
    0.48219368779543, 0.49531434368554, 0.50799480538715, 0.52067439103864, 
    0.5368769670198, 0.54948362296081, 0.56220353500565, 0.57376631365222, 
    0.58667220864103, 0.59870780347244, 0.60949256251469, 0.6208125648111, 
    0.63426475212653, 0.6447704872929, 0.65603817709702, 0.66724014589223, 
    0.67845074693839, 0.68755838284039, 0.69833149253351, 0.70906105754233, 
    0.71755384408088, 0.72901149958955, 0.74050965276531, 0.74823045843879, 
    0.75724402689683, 0.76594613721187, 0.77545762582132, 0.78274304894841, 
    0.79187803066992, 0.80004807926714, 0.80800692078213, 0.81621051281452, 
    0.82477658606713, 0.83214697316486, 0.83933673731919, 0.84661792486106, 
    0.85442862756897, 0.86096428106464, 0.86877487215121, 0.87642655918638, 
    0.88248364078556, 0.89040570302434, 0.89679407388326, 0.90325918721482, 
    0.91034160346142, 0.91701186766087, 0.92318268639865, 0.92956558291689, 
    0.93553451875203, 0.94210059293212, 0.94813544077102, 0.95466468623267, 
    0.96115456845166, 0.96719346393486, 0.97325529382993, 0.97937186227931, 
    0.98542461837622, 0.9914327627175, 0.99717984530605,
  0.99814767151268, 0.99436237937845, 0.99030214330821, 0.98629629532357, 
    0.98226685773514, 0.97791476956081, 0.97373183980114, 0.96920274926398, 
    0.96490651915526, 0.96011812202593, 0.9553066947786, 0.95056163375291, 
    0.9459899394931, 0.94121745720897, 0.9364675217681, 0.93119443713546, 
    0.92604684246711, 0.92057043785842, 0.91508121859473, 0.90977599988474, 
    0.90360741697002, 0.89832804181807, 0.89258975818077, 0.88612117011953, 
    0.88025552542148, 0.87324914177577, 0.86747203094202, 0.86185479795716, 
    0.85418867268671, 0.84786535678711, 0.84129922261042, 0.83302983232809, 
    0.82695252063462, 0.81895134312987, 0.81069963655719, 0.80433833494169, 
    0.79557376359017, 0.78899439386147, 0.77999509504305, 0.77166761581334, 
    0.7629735855639, 0.75410944910188, 0.74536757839113, 0.73402447863296, 
    0.72526932700721, 0.71508782502136, 0.70443720885345, 0.69476153964096, 
    0.68408516028705, 0.67466432351808, 0.66305921187525, 0.65151269613066, 
    0.63936111343916, 0.62651022400069, 0.61433761883621, 0.60178467026351, 
    0.58865285440175, 0.57646342905389, 0.56210971505399, 0.54725940637426, 
    0.53385550514938, 0.51909495728489, 0.50427247410184, 0.48825582132383, 
    0.47114337230353, 0.45847658384388, 0.4421506606671, 0.42419348927051, 
    0.41057438142925, 0.39402920005031, 0.37772489489736, 0.36088476750748, 
    0.34086312731382, 0.32406704771073, 0.30639732535079, 0.28781182040696, 
    0.27111782394653, 0.25629855149333, 0.23601504230726, 0.21917272873763, 
    0.20438469383336, 0.18753995934442, 0.17052773567277, 0.15461418461209, 
    0.13966364696506, 0.12297263786351, 0.10564346329938, 0.094571806135184, 
    0.07966376214628, 0.06802225294903, 0.056700830192037, 0.04724411353578, 
    0.035770055697272, 0.027533660864682, 0.020854338418746, 
    0.014039010505295, 0.008293288637883, 0.0044767245356427, 
    0.00184896342125, 0.00035771423354365, 6.6944183317897e-05, 
    0.0010830272343606, 0.0035027761531408, 0.0071007272492944, 
    0.012491134969965, 0.020168183049715, 0.026938960295738, 
    0.03477320676591, 0.043930814450867, 0.055079915940247, 0.06545992864019, 
    0.078170394167561, 0.090687064021479, 0.10452986482272, 0.12000716214232, 
    0.13603867060723, 0.14988911054579, 0.16902471705807, 0.18495917469684, 
    0.20171856243428, 0.21781762899176, 0.23598247096572, 0.25324586465811, 
    0.26976738127686, 0.28835616201797, 0.30590578725657, 0.32526857581348, 
    0.34023396790844, 0.3586831136763, 0.37664962604872, 0.39296683611456, 
    0.40825234453398, 0.42425770088787, 0.44175227485849, 0.45712634867968, 
    0.47333744369772, 0.49044478494073, 0.50347406874454, 0.51952228574478, 
    0.53404337807394, 0.54781828569063, 0.56141274379161, 0.57481175899015, 
    0.58804842181862, 0.59951580185355, 0.61614079323691, 0.62613353525021, 
    0.63950612995254, 0.65094143783431, 0.66346412174564, 0.67382701915613, 
    0.6845785072031, 0.69455625097286, 0.70518379457829, 0.71671623996613, 
    0.7270751057588, 0.73480429284925, 0.74505927612041, 0.75479412582426, 
    0.76388549944567, 0.77200943159109, 0.77937588972915, 0.78898558884133, 
    0.79783249678416, 0.80538025692611, 0.81195140497581, 0.82121087283158, 
    0.82713668990389, 0.83469351891067, 0.84265132357043, 0.84839389846692, 
    0.85534099930267, 0.86224757676428, 0.86885385165479, 0.87492359938616, 
    0.88077404822145, 0.88608319743704, 0.89282537276507, 0.89847832989526, 
    0.90397648959042, 0.90964680230626, 0.91545747849343, 0.92040968696688, 
    0.92557433268418, 0.93067426531609, 0.93582076010815, 0.94082299209339, 
    0.94564117361287, 0.95013064303473, 0.95512371733482, 0.96003607501063, 
    0.96430610586099, 0.96863059904762, 0.97327369285972, 0.97758888381524, 
    0.98200010285032, 0.98617964030686, 0.99031601309416, 0.99428166693502, 
    0.99813214287104,
  0.99861285056096, 0.99579573675831, 0.99285695591306, 0.9898289477994, 
    0.98676184266498, 0.98356824595431, 0.98028070949945, 0.97687077150761, 
    0.97344548328058, 0.96994052459658, 0.96629303109131, 0.96254238372357, 
    0.95885313703154, 0.95494594846363, 0.95100617889723, 0.94691040867458, 
    0.94292716393148, 0.93866808198418, 0.9342589710786, 0.92980905487631, 
    0.92532277617306, 0.92083910481231, 0.9161542637924, 0.91121186733643, 
    0.90622987884636, 0.90104717440007, 0.89551268518715, 0.89014927891393, 
    0.88508079162233, 0.87910902640213, 0.87322067885306, 0.86694052809627, 
    0.86144427639458, 0.85484525578622, 0.84871353017601, 0.84164652644703, 
    0.83458370003946, 0.82806282014793, 0.82071753355297, 0.81369859907521, 
    0.80575302082242, 0.79829322097971, 0.78987126075566, 0.78218337342601, 
    0.77286425073257, 0.76432484480167, 0.75482664884361, 0.74605293053455, 
    0.73588624467986, 0.72609199816029, 0.71660201887697, 0.70549301944266, 
    0.69409856034974, 0.68260851443545, 0.67201747279352, 0.6591842453287, 
    0.6471651011693, 0.6344716778049, 0.62262208056535, 0.60785423042409, 
    0.59428217123206, 0.58120672104262, 0.56612702849962, 0.55147938655528, 
    0.53665564290403, 0.51944317567534, 0.50478955739758, 0.48713585699242, 
    0.46922348539958, 0.45348908972015, 0.43478702463537, 0.41680090860968, 
    0.40053973364723, 0.38162178815623, 0.36276809945047, 0.3433090877686, 
    0.32194395207012, 0.30605084613263, 0.28531243948376, 0.26530070970908, 
    0.24428724652468, 0.22572522793263, 0.20755398049667, 0.18652194596069, 
    0.16957739526824, 0.15100161578534, 0.13346283272174, 0.11601713215583, 
    0.10047721557673, 0.085087171127906, 0.07027850419727, 0.057688380779929, 
    0.046015224299702, 0.034649774586023, 0.024391128768841, 
    0.017243750680987, 0.009941962762961, 0.0054365365464599, 
    0.0020271102206002, 0.0002722925761981, 0.00016298084470819, 
    0.0016542202993721, 0.0049320427157751, 0.0093678906657911, 
    0.015719183369698, 0.023614607639094, 0.032564638833096, 
    0.04411383615914, 0.054606999051734, 0.067916394559018, 
    0.083931171626956, 0.098111144095082, 0.11393612261289, 0.13116139164703, 
    0.14954377381334, 0.16673486031797, 0.18610649584522, 0.20444644413843, 
    0.22420450820261, 0.24460057094337, 0.26313099703875, 0.28261630158186, 
    0.30195988472037, 0.32221003787189, 0.34230955883759, 0.36077723053401, 
    0.37934536689506, 0.39730631212251, 0.41703498713469, 0.4338435359101, 
    0.45169000618676, 0.46998301288415, 0.48685905882474, 0.50440019857394, 
    0.51793435454658, 0.53546805014006, 0.55092247312571, 0.5655824985703, 
    0.58056837153105, 0.59546019972053, 0.60881708343617, 0.62324041835294, 
    0.63565178798481, 0.64707782944582, 0.65981895521275, 0.67173953254062, 
    0.68290800064246, 0.69491918194153, 0.70619746422367, 0.71638633905058, 
    0.7267342739858, 0.73677837733865, 0.74613642769859, 0.75541353990489, 
    0.76413884525885, 0.77272274798252, 0.78178758853823, 0.7907756027346, 
    0.79789561747717, 0.80620275111461, 0.81361985030674, 0.82171073331228, 
    0.82812501692496, 0.83545815669711, 0.84186501171618, 0.84895864115516, 
    0.85546727403311, 0.86211003481425, 0.86790349886409, 0.87396024998004, 
    0.87981433239759, 0.88535497531267, 0.89080309377288, 0.89592547158453, 
    0.90106022121119, 0.90632617708295, 0.91140994780061, 0.91579756345994, 
    0.92079630612194, 0.92542814086553, 0.92974399614676, 0.9342184071492, 
    0.93827185765925, 0.94253699863816, 0.94658520195014, 0.95043286928781, 
    0.95457506879766, 0.95842579158668, 0.96208040206372, 0.96591642805823, 
    0.9694520651278, 0.97307600905369, 0.97655131450298, 0.97993310044288, 
    0.98327225156045, 0.98658288490861, 0.98977580542617, 0.99283074659729, 
    0.995801174843, 0.99862632757229,
  0.99877620744331, 0.9962603704026, 0.99368110738028, 0.99104171230556, 
    0.98825755116173, 0.98542741552047, 0.98260469988992, 0.97949691723977, 
    0.97647762474483, 0.97327284329383, 0.97018866228677, 0.96685755803692, 
    0.96334974488356, 0.95988965560425, 0.95621971463044, 0.95271469109595, 
    0.94856703289541, 0.9451619689001, 0.94148751781086, 0.93733175765709, 
    0.93275458572773, 0.92824903430556, 0.92441964712193, 0.91970278401325, 
    0.91543078251904, 0.91077383617248, 0.90605389240802, 0.90069654483491, 
    0.89595491261365, 0.89114348513505, 0.88552563144891, 0.87956389149666, 
    0.87370170181975, 0.86885357233387, 0.86289774792493, 0.85584371704065, 
    0.84959036963256, 0.84340904063602, 0.83596289291252, 0.8297117076278, 
    0.82175744085402, 0.81540700935752, 0.80774506044502, 0.79930915751691, 
    0.79159861488289, 0.78295117236049, 0.77573002123268, 0.76564106472631, 
    0.75546677708705, 0.74721307046634, 0.73919782586778, 0.7284778868106, 
    0.71711260954228, 0.70710656680237, 0.69471311206015, 0.68512126749975, 
    0.66937860403931, 0.66039799248614, 0.64640573070245, 0.6349388982875, 
    0.61938173459707, 0.606385798567, 0.59374044676283, 0.57786774431157, 
    0.56115344560806, 0.54613400431589, 0.52905024113387, 0.51231773828764, 
    0.49498996283696, 0.47730069746716, 0.46323450822794, 0.44314925294789, 
    0.42553446060339, 0.40426255425534, 0.38649078399174, 0.3653252407611, 
    0.34854960942663, 0.32645301981949, 0.30670039678029, 0.28534518300372, 
    0.26569214261194, 0.24358608734915, 0.22569411500661, 0.2039434964931, 
    0.18494066326243, 0.1650694877768, 0.1487741500631, 0.12753762131154, 
    0.11044410047884, 0.093017633567466, 0.077897979534659, 
    0.063902522949163, 0.052053818210419, 0.038726255912392, 
    0.027488314881832, 0.01870460292136, 0.011262100383302, 
    0.0061379322412716, 0.0022495262302987, 0.0003676554813297, 
    0.00019816943204844, 0.0020296999777056, 0.0054047378451474, 
    0.010425941230234, 0.017440953716275, 0.028122106118051, 
    0.037897538906734, 0.048829689639568, 0.060670505050691, 
    0.074728660062746, 0.092000646793786, 0.10862209595049, 0.12402126513138, 
    0.14361503926423, 0.16422102871193, 0.18410423559238, 0.20357366847706, 
    0.22222279459958, 0.24067156895229, 0.26280537109167, 0.28635478620123, 
    0.30359168465881, 0.3241026359308, 0.34593253666328, 0.36483727747419, 
    0.38405597328889, 0.40266773355779, 0.42035444027472, 0.44234931899092, 
    0.46153051958943, 0.4779632895002, 0.49716655406714, 0.51381847786916, 
    0.53105213476226, 0.54783206201247, 0.5623839463891, 0.5768264787839, 
    0.58977494054114, 0.60602299173973, 0.62123895684308, 0.63511035491462, 
    0.64633839808733, 0.65704555199018, 0.6717706488238, 0.68454916807967, 
    0.69485653989723, 0.70530364164291, 0.71740632017118, 0.72743096088005, 
    0.73726356518663, 0.7467105780811, 0.75602955457166, 0.76502228373732, 
    0.77572267156361, 0.78375413509076, 0.79159532157452, 0.79959582291457, 
    0.8073957076582, 0.81543747232768, 0.82308291991509, 0.83028772544697, 
    0.83724774533908, 0.84422194711666, 0.85022304537461, 0.85640447688527, 
    0.86255990513911, 0.86889824366049, 0.87470680764178, 0.88062318474729, 
    0.88607767840465, 0.89085404513857, 0.89605206099068, 0.90145148032981, 
    0.90616409722688, 0.91111094871267, 0.91512179589105, 0.91998703797275, 
    0.92436260259661, 0.92880412735687, 0.93269258346476, 0.93676773533469, 
    0.94120543598777, 0.9447991785271, 0.94841006925951, 0.95226076984016, 
    0.95592750640989, 0.95936982874141, 0.96276692055429, 0.96615405754384, 
    0.96960573134261, 0.97285805473321, 0.97608937697825, 0.9791107860723, 
    0.98220601845629, 0.98517017594302, 0.98816108987677, 0.99094069019018, 
    0.99368154997527, 0.99627852384561, 0.99878074599733,
  0.9988986954209, 0.99666679009305, 0.99435651925821, 0.99194741759502, 
    0.9894809199522, 0.98696453028972, 0.98434592611469, 0.98162947409644, 
    0.97893475145833, 0.97594832003283, 0.97315196629002, 0.96999772293683, 
    0.96700040249519, 0.96387929985783, 0.96059705047633, 0.9572150282039, 
    0.95391761703782, 0.95031607203944, 0.94671688813128, 0.94311161622011, 
    0.93945904015592, 0.93546655766849, 0.93155860091228, 0.9276486623518, 
    0.92331726964922, 0.91917026498092, 0.9146920234996, 0.90967101123437, 
    0.90535105186212, 0.90053901826278, 0.89521023525373, 0.8904946493747, 
    0.88495533966871, 0.87973866497319, 0.87427048950301, 0.86849881043191, 
    0.86248301010286, 0.8561432734497, 0.84993568434742, 0.84353564138667, 
    0.83696459171324, 0.82943371738704, 0.82283253239855, 0.81556053193954, 
    0.80711418586006, 0.7997950770537, 0.79179699814498, 0.78254196292157, 
    0.77385478560023, 0.76565295101492, 0.75604598172568, 0.7465210387468, 
    0.73607905290364, 0.72594399014843, 0.71530724793278, 0.70381140192774, 
    0.69286578955141, 0.68120476103672, 0.66874933481304, 0.65556423671754, 
    0.64205206436972, 0.62901145603972, 0.61543872888414, 0.60063679743901, 
    0.58582357121403, 0.57013775232267, 0.55386928474917, 0.53692728450572, 
    0.52125487970737, 0.50429543649298, 0.48347630119107, 0.46657102646498, 
    0.44797307493907, 0.42893444059672, 0.40808863351177, 0.38873904844642, 
    0.37006662121177, 0.34708810889496, 0.3269094455893, 0.30609488667998, 
    0.28408534785971, 0.26314331234441, 0.24123989672946, 0.21947318357471, 
    0.20013797976564, 0.17714909533965, 0.15754397243357, 0.13782935034262, 
    0.12129141786185, 0.1014001566081, 0.084780865347584, 0.068580645788001, 
    0.05522833730704, 0.04185781863054, 0.029902365901849, 0.021557159870983, 
    0.01257889247301, 0.0063519855054893, 0.0023835046895358, 
    0.00037007354614865, 0.00017967765369593, 0.0019545352058555, 
    0.0060065295570897, 0.011455002005796, 0.019617220962084, 
    0.029194443743698, 0.039882922526259, 0.053764241065387, 
    0.068698656433083, 0.082252763630146, 0.099694049668901, 
    0.11698366871575, 0.13700364181035, 0.15481083005862, 0.17582213029076, 
    0.19593760317835, 0.21830663210907, 0.23879847638125, 0.25934168725973, 
    0.28360190755115, 0.30262392633957, 0.32493591498728, 0.34579841307716, 
    0.36660477758903, 0.3880137705043, 0.4082867975045, 0.4282235583296, 
    0.44659941401636, 0.46749750725358, 0.48327027400112, 0.50180913524636, 
    0.52082084201033, 0.53721185121411, 0.5531233224264, 0.56944055279145, 
    0.58536056108565, 0.59956635796899, 0.61492260616937, 0.62896992556441, 
    0.64311694039133, 0.65591011788791, 0.66746472672448, 0.68093071871523, 
    0.69274426889308, 0.70489510350209, 0.71532314256459, 0.72661726445601, 
    0.73685149477052, 0.7472931471236, 0.75566064217877, 0.76555819417338, 
    0.77445174190755, 0.78295854155464, 0.79237151522495, 0.80055926547643, 
    0.80785324263924, 0.81589804713378, 0.82290837291432, 0.83036229084783, 
    0.83694614784656, 0.84393154393367, 0.84991596159299, 0.85647559143616, 
    0.86321446015652, 0.86847703625672, 0.87451223300155, 0.88003835036133, 
    0.88497591937454, 0.89018282914397, 0.89591825757472, 0.90079345858254, 
    0.90538385705081, 0.91010865425977, 0.91447658025555, 0.91875163951767, 
    0.92306341966339, 0.92748738005878, 0.93125481281765, 0.93537681537094, 
    0.93899951917315, 0.94298491254314, 0.94632828871357, 0.94992331071679, 
    0.95353754859109, 0.95684424372439, 0.96013434886719, 0.96344077606306, 
    0.96652909209885, 0.96961275647352, 0.97268372674107, 0.97563417607018, 
    0.97851758128088, 0.9813821528057, 0.98408099583994, 0.98673166509019, 
    0.98935470207358, 0.99189454563474, 0.99431487380711, 0.99667679290915, 
    0.99890455252486,
  0.99908924657294, 0.99725952522584, 0.99531230560407, 0.99337138799659, 
    0.99125799274003, 0.98910180696998, 0.98697874819151, 0.98487073209134, 
    0.9824783192631, 0.98007520614549, 0.97766458855261, 0.97516716646397, 
    0.97239755997642, 0.96998187160214, 0.96701149640263, 0.9641403323999, 
    0.9614838634038, 0.95844790865143, 0.95547863459667, 0.9524041674845, 
    0.94885282604555, 0.94575971694891, 0.94249108660855, 0.93898996080088, 
    0.9354757763982, 0.93141029446915, 0.92793798396925, 0.92379528156376, 
    0.91990625039591, 0.91522367152558, 0.91098134294061, 0.90677605494885, 
    0.9024670645535, 0.89759034126896, 0.89273921441991, 0.88744506024035, 
    0.88220879461534, 0.87640022914358, 0.87111228420168, 0.86548774709256, 
    0.85934090599455, 0.85376386041592, 0.84750327265746, 0.84113038643884, 
    0.833476479692, 0.82648018554852, 0.81983153187295, 0.81041278082904, 
    0.80363406395476, 0.79627440569506, 0.78676221681651, 0.77785881325409, 
    0.76874935193652, 0.75992977853683, 0.74944864838148, 0.73810758749719, 
    0.72857602660406, 0.71668591969059, 0.70540498816302, 0.69377361211052, 
    0.6813519783344, 0.66883741526378, 0.6550597666261, 0.640719257648, 
    0.62672844355037, 0.61238637363019, 0.59595531725267, 0.58019735820175, 
    0.56250825476394, 0.54466189061671, 0.52739295898696, 0.50914645731433, 
    0.49152587877129, 0.47179797119335, 0.44956601979179, 0.43035606289132, 
    0.40641152443831, 0.38653981178058, 0.36260772205307, 0.34158118142011, 
    0.31844045371072, 0.2944208470987, 0.2739322287363, 0.25173311314936, 
    0.22565308805416, 0.20340747127288, 0.18307083522446, 0.16113233553025, 
    0.14036027515088, 0.1193015682008, 0.097702954380163, 0.080083776909903, 
    0.064537113303247, 0.048993595022275, 0.035417428149556, 
    0.022977490896104, 0.014136726825853, 0.0078884223060174, 
    0.002688830851535, 0.00025266936611423, 0.0002054123251789, 
    0.0024819826692761, 0.0075423341419045, 0.014111420048125, 
    0.023235931461428, 0.033713461799235, 0.046819302954625, 
    0.063906280771745, 0.08071416927138, 0.097415070482305, 0.11603155822584, 
    0.13450907092228, 0.15815440287648, 0.17956602450329, 0.20137741084402, 
    0.22281699332278, 0.247868867418, 0.27109872605076, 0.29267293439832, 
    0.3170854532343, 0.34003742609072, 0.3633537725398, 0.38611399440606, 
    0.40550669866219, 0.42701295883425, 0.4483598197472, 0.46877461020971, 
    0.48969022419444, 0.50838660088367, 0.52432445419761, 0.54512305030785, 
    0.56327518442421, 0.58140939192035, 0.59530789556687, 0.61056777456494, 
    0.62522592448252, 0.64165542623018, 0.65562751494762, 0.66827252630267, 
    0.68166535373692, 0.69311416001672, 0.70554441337111, 0.718354934017, 
    0.72843768003973, 0.73855344120321, 0.74936731068738, 0.75936464471792, 
    0.76886861438763, 0.77818130543651, 0.7877365451852, 0.79551054942137, 
    0.80386877339106, 0.81151963341274, 0.81911152823112, 0.8270945394198, 
    0.83500497604076, 0.84101366229417, 0.84740349240648, 0.85443549507653, 
    0.86056124043295, 0.86623761135825, 0.87109012383126, 0.87703496378757, 
    0.8822715469431, 0.8882459377691, 0.89294877256325, 0.89781243321274, 
    0.90203026237684, 0.90694792505882, 0.91176898678937, 0.91593069501146, 
    0.91989501618575, 0.92383090983004, 0.92745260869478, 0.93076910955472, 
    0.93499199996422, 0.93882569694302, 0.9418901685638, 0.94553021076872, 
    0.94820447189301, 0.95188159888282, 0.9553189038853, 0.95823508579767, 
    0.96111345508103, 0.96400635459119, 0.96675714644206, 0.96947230568973, 
    0.97207407033479, 0.97467629709201, 0.97718122007843, 0.97976909638071, 
    0.9821117915204, 0.98463858757947, 0.98687917407654, 0.98904131715136, 
    0.99118358565757, 0.99328968884453, 0.99532305422748, 0.99724495348898, 
    0.99909111896233,
  0.9992208299603, 0.99763546286272, 0.99601861184038, 0.99437321904702, 
    0.99264659941441, 0.99075200864622, 0.98888143616418, 0.98699220185897, 
    0.98506973510033, 0.98295330639267, 0.98086449497745, 0.97880492782488, 
    0.97660962075607, 0.97420284352931, 0.97162327340479, 0.96938291100541, 
    0.96673358095466, 0.96442924394336, 0.96189004327382, 0.9590114805556, 
    0.95636639884192, 0.95346731290747, 0.95054140191457, 0.94740381337954, 
    0.94452342935108, 0.94099838407581, 0.93770081475132, 0.9341734910054, 
    0.9305817101063, 0.92662774953506, 0.92330385854595, 0.91955992446217, 
    0.9154114133142, 0.91066976084544, 0.90672953607532, 0.90243699583312, 
    0.89809618577002, 0.89287244404335, 0.8872411866953, 0.88239094781806, 
    0.87664501463466, 0.87151790213511, 0.86562551454189, 0.85970553213109, 
    0.8539246045718, 0.84757948501696, 0.84102992418408, 0.83322717704771, 
    0.82568059381584, 0.81812402780636, 0.81121915382828, 0.80347854707084, 
    0.7950423918828, 0.78621700977026, 0.77579229096582, 0.76726369403268, 
    0.75728551753152, 0.74561558463244, 0.73587746927806, 0.72459881898192, 
    0.71203388594586, 0.70104148802516, 0.68626539293571, 0.67429084796871, 
    0.66141076018292, 0.64832558459386, 0.63087264817104, 0.61326355368815, 
    0.60038441667072, 0.58219936196231, 0.56674503703561, 0.54424232865193, 
    0.52572041182366, 0.50837640945422, 0.48786616854057, 0.46731333752455, 
    0.44398950470329, 0.42213974425074, 0.39939915382439, 0.37420115564337, 
    0.35155781998736, 0.32851977082203, 0.30361919165654, 0.27890709107929, 
    0.25141841931813, 0.22689106912135, 0.20518037164704, 0.18022311391072, 
    0.15671542581141, 0.13179307053381, 0.11132626830963, 0.090854621756679, 
    0.072659147806143, 0.056779492489789, 0.040315487622113, 
    0.027439183745195, 0.016887218940027, 0.0084083166898326, 
    0.0032498203588929, 0.00052365125935483, 0.00026542263321509, 
    0.0031513301291744, 0.0079318832596368, 0.016341770705387, 
    0.026176114930837, 0.038796645331059, 0.053687373278434, 
    0.072137633342046, 0.090524807776533, 0.11062262402812, 0.13334311028638, 
    0.15288007865224, 0.17813803725267, 0.20167037809664, 0.22981338212895, 
    0.25097523139452, 0.27591126603319, 0.30187282717746, 0.32428499385518, 
    0.34880447465702, 0.37356293209636, 0.39701784884286, 0.41919081763308, 
    0.44299659292628, 0.46324123152752, 0.48772955893568, 0.50687944884232, 
    0.52653744958662, 0.5459037383176, 0.56423605007117, 0.5810440205862, 
    0.59887498782169, 0.61519506190303, 0.63146284454231, 0.6457356614303, 
    0.6598603141904, 0.67430012068153, 0.68922117995366, 0.69996139615013, 
    0.7135349799498, 0.72470931381189, 0.73709689716547, 0.74811820506993, 
    0.756656950183, 0.76793725692974, 0.77726954053962, 0.78682995744589, 
    0.79450789349287, 0.8028142050663, 0.811691057624, 0.81892515026349, 
    0.82709253900516, 0.83334153490156, 0.83969428743895, 0.84712912017684, 
    0.8531423981317, 0.8612062399438, 0.86672550646455, 0.87223450391911, 
    0.87747211161438, 0.88265659922983, 0.88789023432227, 0.89308056333085, 
    0.89810520460498, 0.90263672786431, 0.90605996284701, 0.91080744303087, 
    0.91518476942536, 0.91904286995379, 0.92296575942325, 0.92715958229852, 
    0.93038176580524, 0.93419339049621, 0.93743945690566, 0.94059371501929, 
    0.94375496399952, 0.94721394807476, 0.95023574549642, 0.95312338596511, 
    0.95565965030321, 0.95853351057205, 0.96128199755769, 0.96407034989122, 
    0.966666788187, 0.96916120771637, 0.97141348888654, 0.97368616272246, 
    0.9762970679672, 0.97846298934495, 0.98055819133116, 0.98269376596357, 
    0.98482799882212, 0.98682133641632, 0.98877457836107, 0.99065390340643, 
    0.99249108007623, 0.99431677582229, 0.99600528074094, 0.99766333693285, 
    0.99922829633766,
  0.99932118903704, 0.99795070436907, 0.9965281240534, 0.99505498868699, 
    0.99354454974144, 0.99197376850312, 0.99031254369763, 0.98866585810565, 
    0.9869329421259, 0.98519174323628, 0.98337508670757, 0.98143996906086, 
    0.97955388353184, 0.97756527199509, 0.97542023855394, 0.97335808303524, 
    0.97109751528443, 0.9688484015235, 0.9667053503409, 0.96417992178606, 
    0.96180824226159, 0.95904866619441, 0.95664003938465, 0.95390613669823, 
    0.95112762373411, 0.94811334066891, 0.94508461703086, 0.94195431860925, 
    0.93884727118993, 0.93580085399502, 0.93231084819054, 0.92873386547019, 
    0.92524022981103, 0.92146015569303, 0.91747668160318, 0.9135305261456, 
    0.90939268576277, 0.90510527510766, 0.900572975577, 0.89583509729056, 
    0.89073762672556, 0.88566412019246, 0.8805210317901, 0.87528698539281, 
    0.86978682869631, 0.86383289587607, 0.85728637537965, 0.85140690623285, 
    0.844865277865, 0.83767804282743, 0.83078219747936, 0.82334763928464, 
    0.81490501467553, 0.80673513300808, 0.79881685657572, 0.79003280334135, 
    0.78072435410256, 0.77002298678832, 0.76040490628793, 0.75007060171205, 
    0.73865697939201, 0.72796480016744, 0.71528317706075, 0.70148753193914, 
    0.68993998371157, 0.67642615588208, 0.66068421876471, 0.64514729810713, 
    0.62978471628319, 0.61355706706067, 0.59458397790104, 0.57800328413883, 
    0.55933303524983, 0.53971533038651, 0.51846917438011, 0.49910795425926, 
    0.47497913353425, 0.45274763218307, 0.43061140538936, 0.40619646343779, 
    0.38153993441082, 0.35469621436591, 0.33025523476685, 0.30481216022413, 
    0.27751287947527, 0.25250104857959, 0.22396151910473, 0.19886800851497, 
    0.17381061313516, 0.14976967560116, 0.12389901182519, 0.10425145977757, 
    0.081707071487237, 0.062653113667763, 0.046363124321486, 
    0.031105444134537, 0.019262995690838, 0.010125426201044, 
    0.0038350663091563, 0.00042510032693104, 0.00040506850224813, 
    0.0033175554931017, 0.0099404368744311, 0.018263734893068, 
    0.029468146825304, 0.044527124735294, 0.062361303005733, 
    0.080051970214578, 0.10041797662322, 0.12404791115417, 0.14822090103722, 
    0.17281440075739, 0.19758500559605, 0.22521043056811, 0.24955899386316, 
    0.27706531263799, 0.30307412423716, 0.3284415715341, 0.35298340088445, 
    0.37932926522903, 0.40423776021879, 0.42949701848463, 0.4521835129814, 
    0.47492502779332, 0.49554576975561, 0.51852320117998, 0.53964233687101, 
    0.55855151669911, 0.57777433965297, 0.59549772700198, 0.61244981058643, 
    0.62933338226012, 0.64548586258374, 0.66087938777823, 0.6745075635302, 
    0.68887517648105, 0.70177714660997, 0.71438003549059, 0.72806370546399, 
    0.73896375566832, 0.7504528435362, 0.76043272289415, 0.77119321637388, 
    0.7804601991061, 0.79034775955575, 0.79881762505844, 0.80778837678533, 
    0.81571890582949, 0.82352875101352, 0.83040795922537, 0.83834217865687, 
    0.84479460828417, 0.85185267731893, 0.85838811938507, 0.86441013778923, 
    0.86941853271594, 0.87584959871292, 0.88112290688088, 0.88586752982085, 
    0.89124788492476, 0.89594744579363, 0.90092209371432, 0.90491506431109, 
    0.90953561111234, 0.91382257548889, 0.91768401431689, 0.92142764075305, 
    0.92517700559538, 0.9287340501626, 0.93224803343564, 0.9354418879819, 
    0.93874575837852, 0.94155397568264, 0.94492003174714, 0.9477843658454, 
    0.95073637094827, 0.9535318805539, 0.95610735523059, 0.95883957016074, 
    0.96117583445248, 0.96377790571332, 0.96616543780291, 0.96840850756277, 
    0.97077497161007, 0.97289924802716, 0.97500945020583, 0.97716757171229, 
    0.97921677268565, 0.98110090630282, 0.98307792991792, 0.98497238588132, 
    0.98675361544295, 0.9885224965502, 0.99022138322957, 0.99190303802653, 
    0.99348998151729, 0.99503999577203, 0.99652579261658, 0.99795392758298, 
    0.99932210187598,
  0.9993980182726, 0.99818847232616, 0.99693331065357, 0.99563820205435, 
    0.99427040888939, 0.9929133008372, 0.99144898155048, 0.98996712090901, 
    0.98849634786151, 0.98681816913556, 0.9852214882016, 0.98358272909721, 
    0.98188857484029, 0.98006706889824, 0.97828005107426, 0.97633300536784, 
    0.97439262386544, 0.97235492628201, 0.97032814497532, 0.96817950719683, 
    0.96585184573056, 0.96375407088585, 0.96148725209338, 0.95897950332748, 
    0.95642852645741, 0.95394699546942, 0.95113866498573, 0.94841887413114, 
    0.9453421824165, 0.94255396811377, 0.93980972214572, 0.93645658624352, 
    0.93323039835443, 0.92952367260514, 0.9261476082911, 0.922494209644, 
    0.9190917673228, 0.91470214726508, 0.9105811398265, 0.90655155897109, 
    0.9021568686204, 0.89733006430215, 0.89263846616615, 0.88800357391811, 
    0.88237766809956, 0.87686880828675, 0.87131909322654, 0.86507692313049, 
    0.85901888471584, 0.85357584971923, 0.84550547723338, 0.83920798412965, 
    0.83286895671702, 0.82506841231126, 0.81730909886244, 0.80896436381137, 
    0.80039792937954, 0.79101043229916, 0.78098486662973, 0.77127602162882, 
    0.76142006849667, 0.74978205525493, 0.73845865322624, 0.72525640429889, 
    0.71424555302882, 0.6999691162964, 0.68665639425609, 0.6711468608356, 
    0.65654438991079, 0.64034110689975, 0.62394210213668, 0.60661573456916, 
    0.58727836103819, 0.56843699527546, 0.5469582991334, 0.52636283171524, 
    0.50378094535978, 0.48188894223637, 0.45788835832315, 0.43375290377556, 
    0.40921621391717, 0.38181885966436, 0.35576848550609, 0.32748573326546, 
    0.30167954651763, 0.2722083983499, 0.24632150481106, 0.21909452369407, 
    0.19258765423486, 0.16401883451098, 0.13897294918693, 0.11514159749815, 
    0.091557128112922, 0.0696979936275, 0.050469498233956, 0.035007555708209, 
    0.021302933842064, 0.011166489818349, 0.003783110271238, 
    0.00042957078594356, 0.00042471714685313, 0.0037319029912618, 
    0.010584053253882, 0.02104129501592, 0.034024515757891, 
    0.049437242417331, 0.068567272589111, 0.089227533550385, 
    0.11239546100836, 0.13717597708069, 0.16147935088768, 0.18829868762475, 
    0.21443705030898, 0.24474118784166, 0.27217230822667, 0.29830574713425, 
    0.32619153196423, 0.35505600105991, 0.38107782356642, 0.40747449163358, 
    0.43253417838019, 0.45819477870779, 0.48317210757418, 0.50448863880975, 
    0.52722254376378, 0.54720578849341, 0.56793352104452, 0.58841911139631, 
    0.60705104654892, 0.62326704234323, 0.63920052747558, 0.65581378795132, 
    0.67201146315092, 0.68643701095834, 0.70032746113263, 0.71351841723375, 
    0.72587710648706, 0.73843391378203, 0.74993505017252, 0.76075649878762, 
    0.77120194401318, 0.78118341599305, 0.7908181598594, 0.80025885327757, 
    0.80875778760355, 0.81724314316463, 0.82608233890409, 0.83295436484056, 
    0.84002197507878, 0.84677505540514, 0.85362510458335, 0.86014284093879, 
    0.86647385723131, 0.87200916541519, 0.87771590232001, 0.8833197963019, 
    0.88802068040973, 0.89267759686286, 0.8975196526146, 0.90217790177866, 
    0.90661690899644, 0.91073610055833, 0.9147317344472, 0.91865857880025, 
    0.92283106519597, 0.92611411634147, 0.92970351948128, 0.93301299029984, 
    0.9363176295978, 0.93927034334573, 0.94248707571672, 0.94527584514399, 
    0.94821285216789, 0.95084768717603, 0.9534399843097, 0.95595123836627, 
    0.95858154082966, 0.96098360504204, 0.9632958377344, 0.96547771422703, 
    0.96772012329635, 0.96990245203331, 0.97207876605069, 0.97410771878074, 
    0.97585524855362, 0.97795852042891, 0.97970461843695, 0.9815789728621, 
    0.98321313635466, 0.9850669759121, 0.98666589096294, 0.98828256844151, 
    0.98983776912446, 0.9913608646154, 0.99279835068055, 0.99424236627491, 
    0.99561245550582, 0.99691214309983, 0.99818779070659, 0.9993980705979,
  0.99950828754242, 0.99852368333019, 0.99750395080499, 0.99644554634985, 
    0.99536963588477, 0.99424556050328, 0.99307088909586, 0.99188271659078, 
    0.9906585059478, 0.98936728340029, 0.98805732974583, 0.98668605474253, 
    0.98529189717893, 0.98383787452434, 0.9823219950274, 0.98082747084528, 
    0.97918672204276, 0.97753223707668, 0.97587118306735, 0.97413962778324, 
    0.97223014200499, 0.97032371154907, 0.96850641365885, 0.96642250987534, 
    0.96438359930306, 0.96233285091386, 0.96003196501667, 0.9576103821409, 
    0.95537391842792, 0.95299509560169, 0.95014813759078, 0.94774208821759, 
    0.94493132043385, 0.94192437151353, 0.93914744837957, 0.93592017677968, 
    0.93273257846921, 0.92931363646796, 0.92615186639642, 0.92232684944729, 
    0.91854304133233, 0.91466749516139, 0.91055509151232, 0.90617868782, 
    0.90194726559014, 0.89726539470909, 0.89245677956044, 0.88728662369893, 
    0.88180241388552, 0.87667617726424, 0.87104578797067, 0.86473513114747, 
    0.85816197103613, 0.85188467900452, 0.84483124915905, 0.83747152610123, 
    0.82968745573958, 0.82174984764713, 0.81376358027974, 0.80460406294477, 
    0.79558098231045, 0.78475769784321, 0.77564836322062, 0.76266840206349, 
    0.75294654823703, 0.74047793464268, 0.72720363467293, 0.71413304179397, 
    0.70030015017109, 0.68445213980013, 0.6688183490948, 0.65261397645179, 
    0.63495604907959, 0.61590264990686, 0.59650032707952, 0.57483570507831, 
    0.55394755760663, 0.53263689833753, 0.50794315477207, 0.48503886805686, 
    0.45927820961215, 0.43079465213178, 0.40235463444501, 0.37377137527164, 
    0.34603427541905, 0.31354794132814, 0.28287611711544, 0.25423617258496, 
    0.22343497724218, 0.19235067003581, 0.16343041582936, 0.13440961926293, 
    0.10795196122992, 0.082982104339698, 0.062022338315166, 
    0.042258193550143, 0.026566563220862, 0.013685700119011, 
    0.0049977011184054, 0.00063481694910351, 0.00055940558508243, 
    0.0045131975639759, 0.013533874229394, 0.025228026115332, 
    0.040814541956113, 0.060033885489192, 0.081815717076627, 
    0.10659775675717, 0.13401799592832, 0.1615484363227, 0.19046876589179, 
    0.22082417763534, 0.25214624156197, 0.28249841877561, 0.31239829017953, 
    0.34115004256059, 0.37318098053388, 0.40044693264164, 0.42947427522065, 
    0.45514032142669, 0.48197921264153, 0.50747514290383, 0.53186936486501, 
    0.55380263639419, 0.57508379689101, 0.59541981852934, 0.61622028858232, 
    0.63455813135175, 0.65197060428324, 0.66800942908431, 0.68491189926803, 
    0.69892040282136, 0.71455725412324, 0.72805875072803, 0.74146769735102, 
    0.75280019767635, 0.76350644725615, 0.77553267746923, 0.78586281011881, 
    0.79565535847369, 0.80585361366006, 0.81438645468894, 0.82251872135502, 
    0.83104144576928, 0.83824897860508, 0.8462259932931, 0.85276642430192, 
    0.85975023619752, 0.86559250118101, 0.87181701780563, 0.877060115813, 
    0.88287515198705, 0.88829778842114, 0.89344248496884, 0.89803319716752, 
    0.90239258766255, 0.90686130941895, 0.91138970839261, 0.91518355799404, 
    0.91925630999194, 0.92269736241978, 0.92632644215125, 0.92956173899303, 
    0.93300314476133, 0.93616241207266, 0.93925037650437, 0.9422206679465, 
    0.94475137157379, 0.9476711730242, 0.95008988169717, 0.9526008223638, 
    0.95501286713269, 0.95746673917635, 0.9597154184633, 0.96187980577772, 
    0.96416672536639, 0.96606734266066, 0.9680994637184, 0.97006453263255, 
    0.97184931443603, 0.97373495707085, 0.9753873734816, 0.97715503681246, 
    0.97883713168961, 0.98043337455471, 0.98205916441186, 0.98355749986843, 
    0.98498274550127, 0.98643847441392, 0.98784861603722, 0.98915440948267, 
    0.99049649386241, 0.99176524649682, 0.99298451669849, 0.99417244668462, 
    0.99532580325673, 0.99643548424025, 0.9975019847861, 0.99852666590625, 
    0.9995092337894,
  0.99954909180101, 0.99864828240225, 0.99774358110474, 0.99679215904402, 
    0.99577800181685, 0.99473274884893, 0.99367525238539, 0.99259255403789, 
    0.99144065126587, 0.99028590571503, 0.98910506833846, 0.98778506919545, 
    0.98658768963159, 0.98530393406905, 0.98393670528119, 0.98244289447468, 
    0.9810538936495, 0.97956832041115, 0.97798067508149, 0.9762584254169, 
    0.97450772327418, 0.97279782295938, 0.97108194349934, 0.9693794845078, 
    0.96747067108056, 0.96526662530245, 0.96320977799599, 0.96124142130619, 
    0.95909018703833, 0.95678737974206, 0.95443305412643, 0.95199151775402, 
    0.94988124224481, 0.94677665545959, 0.94374535576137, 0.94094852994204, 
    0.93810692204309, 0.93482166691344, 0.9318843149594, 0.9285243495406, 
    0.92518369063102, 0.92124589371119, 0.91763403813205, 0.91363264260501, 
    0.90973033550333, 0.90488282972387, 0.90003672590467, 0.89626735904976, 
    0.89068939108387, 0.88549937554629, 0.8797868779612, 0.87431856874437, 
    0.86879367535147, 0.86282876007251, 0.85573590148054, 0.84926721288809, 
    0.84103886019389, 0.83357521164444, 0.82645503513823, 0.81748290155653, 
    0.80880040952978, 0.79936626173335, 0.79087182657526, 0.77992944060319, 
    0.76799092756599, 0.75697597171344, 0.74503627576186, 0.73162570622477, 
    0.71806162296064, 0.70363602835783, 0.68714195844775, 0.66896094422498, 
    0.65341186594349, 0.6372678419678, 0.61878574799224, 0.59780672533282, 
    0.57485814590718, 0.55469740883841, 0.53124233280267, 0.50554962730922, 
    0.47925136389356, 0.45138293939758, 0.42047371391752, 0.39351172113518, 
    0.36281080242179, 0.33331282575859, 0.30304018160768, 0.26900465255607, 
    0.24002184694207, 0.20583703251736, 0.17690933369537, 0.14577765081501, 
    0.11665194551086, 0.091451790217217, 0.066885631061746, 
    0.045967952970523, 0.029098808054381, 0.015094453213688, 
    0.0057875971852027, 0.00042991545863792, 0.00050394384889974, 
    0.0053214158845594, 0.013102818180905, 0.026038851172782, 
    0.043523321888511, 0.064573719688769, 0.089666424666633, 
    0.11667963893416, 0.14473709133299, 0.17272368503046, 0.20537867198671, 
    0.23805778902598, 0.26638647570355, 0.30106712689783, 0.33365012981758, 
    0.35988156116316, 0.39176245425434, 0.42126494498761, 0.45199184407345, 
    0.47812328387631, 0.50391154952326, 0.52583677399697, 0.5525761287216, 
    0.57656805172003, 0.59623171552207, 0.61717762628728, 0.6375072303593, 
    0.65400988741148, 0.67075354714776, 0.68738566223136, 0.70429972534813, 
    0.71853618550361, 0.73285832736687, 0.7438197001222, 0.75693907939295, 
    0.76946544281857, 0.77984618030082, 0.79161195538207, 0.80024572883464, 
    0.80975039514096, 0.81905380697995, 0.82645840256804, 0.83469874825725, 
    0.84277365780839, 0.85056837097875, 0.85735437512697, 0.8636248661342, 
    0.8700293933823, 0.87537483174607, 0.88126686700204, 0.88578520668003, 
    0.89178892203825, 0.89710586540774, 0.90145377476934, 0.90599487198162, 
    0.91047444331616, 0.91435234702993, 0.9178695769491, 0.92191993959787, 
    0.92540197571232, 0.92894777383077, 0.93224531620695, 0.93544721972171, 
    0.93850433888502, 0.9413052778592, 0.94408540993387, 0.94634251463545, 
    0.94981527434903, 0.95207818078267, 0.95419993271779, 0.95637839773459, 
    0.95893980523332, 0.96099036174177, 0.96313336018473, 0.9649537364908, 
    0.96702593214869, 0.96891987795711, 0.97083223244249, 0.97275460409152, 
    0.97439277048942, 0.97603844991106, 0.97761782857823, 0.97911891417453, 
    0.98058688766462, 0.98205378649934, 0.98350194737574, 0.98500403516496, 
    0.98629422480647, 0.98772292704229, 0.98892445285259, 0.99007262984877, 
    0.9912406094901, 0.99244351542716, 0.99361733972097, 0.99469451096484, 
    0.99573700677856, 0.99674069232343, 0.99770629138802, 0.99864841456529, 
    0.99955196945795,
  0.99958472022222, 0.99875617580304, 0.99790302980024, 0.99701571373087, 
    0.99610103137352, 0.99515502328224, 0.99418448984686, 0.99317841664794, 
    0.99212824101026, 0.99105378384256, 0.98996917405524, 0.98880739274877, 
    0.9876221459163, 0.98642623564133, 0.98518409082912, 0.98381170502903, 
    0.98249169205563, 0.98106374296266, 0.97969123040803, 0.97818361395141, 
    0.97663233372795, 0.97505996790139, 0.97338380381993, 0.97159780174967, 
    0.96999254029165, 0.9680337946301, 0.96615347141302, 0.9641972476451, 
    0.96215693410963, 0.96002986104123, 0.95786140585542, 0.9557068021779, 
    0.95315933094488, 0.95079471523751, 0.94821374125743, 0.94535279759852, 
    0.94288900035377, 0.9397767120554, 0.93690898921406, 0.93362340367548, 
    0.93038152345333, 0.92741658025104, 0.92360494658625, 0.9194742605277, 
    0.91598027324589, 0.91166703800301, 0.90767325847688, 0.90323374866076, 
    0.89876362215504, 0.89386521966757, 0.88846866721254, 0.8832917399862, 
    0.87765429474945, 0.87211052967427, 0.86560047478234, 0.85901190710888, 
    0.8522931117043, 0.84519921664891, 0.83743267471583, 0.82893788288316, 
    0.8210470875604, 0.8131519526838, 0.80263784150198, 0.7928784614552, 
    0.78229783280943, 0.77019378367757, 0.7596780467186, 0.74665683474692, 
    0.7332897204685, 0.719645423872, 0.70496365516578, 0.68927361585404, 
    0.67194437565266, 0.6550965491388, 0.63551569850014, 0.61582512036187, 
    0.59461263628707, 0.57135203872662, 0.5486328685272, 0.52377492013812, 
    0.50016113016437, 0.4726711255051, 0.4440767675013, 0.41277287795715, 
    0.38342868903239, 0.35116867648514, 0.3201931367775, 0.28668669667952, 
    0.25250176866025, 0.22216688409783, 0.18753512085686, 0.15493739731426, 
    0.12459104528691, 0.097759980613579, 0.071781875167938, 
    0.049327217513889, 0.031170457577859, 0.015651880476766, 
    0.0057589944668637, 0.00070878005346702, 0.0006013002900991, 
    0.0054257830467411, 0.015356969002958, 0.029556893448958, 
    0.048134580110359, 0.070098862065261, 0.095389111809129, 
    0.12243092243473, 0.15436792668265, 0.18587286703926, 0.21810982668683, 
    0.25175724989031, 0.28313160411301, 0.31760239009435, 0.34943244245697, 
    0.38107374384678, 0.41326497127073, 0.44064473000953, 0.47028273574653, 
    0.49661749720744, 0.52324098317385, 0.54884577658148, 0.57262097769923, 
    0.5955482878801, 0.61373784922523, 0.63651303249892, 0.6550977808342, 
    0.67202155413738, 0.68893907106728, 0.70425935785289, 0.71901624856121, 
    0.73488792457285, 0.74781987066311, 0.7603982356559, 0.77204957330668, 
    0.78234283433874, 0.79353139234393, 0.80411379841441, 0.81346635432654, 
    0.82169053488254, 0.83084000144602, 0.83834977762111, 0.84602749997208, 
    0.85319550344744, 0.860426385202, 0.86704842564337, 0.87289064473338, 
    0.87888004216978, 0.88449623451968, 0.88970753877301, 0.89454849930353, 
    0.89960680587631, 0.90397180361233, 0.90854088984023, 0.91288544430896, 
    0.91684298702888, 0.92035831473695, 0.92413793882122, 0.92756853084818, 
    0.93110726459495, 0.93397332178397, 0.93715636259045, 0.94025418448982, 
    0.94293942056886, 0.94582661049677, 0.948278974707, 0.95079090683689, 
    0.95316827498538, 0.9555137426888, 0.9578072111108, 0.95989228762735, 
    0.96198890027685, 0.9640457398275, 0.96593963953155, 0.96792004836485, 
    0.96954331105062, 0.97139277656636, 0.97305975815523, 0.97471312770833, 
    0.97626898904759, 0.97788912604429, 0.97935587621107, 0.98079314556395, 
    0.98220992610114, 0.98356994492599, 0.98486428439576, 0.98615324117272, 
    0.9874128087714, 0.98859995226659, 0.9897881755935, 0.99090128434228, 
    0.99201960183814, 0.99307741038738, 0.99410003137594, 0.99510905229948, 
    0.99606845474104, 0.99699539395189, 0.99789556559998, 0.99875447965642, 
    0.99958507360497,
  0.99964147505979, 0.99893326358365, 0.99820427376276, 0.99741324908164, 
    0.9966183037232, 0.9958046229403, 0.99498208458987, 0.99413483174929, 
    0.99328184440939, 0.99230541134567, 0.99135847445044, 0.99036549698867, 
    0.98936974730614, 0.98823971840374, 0.98719502048206, 0.98607130397794, 
    0.98485810205923, 0.98365801618755, 0.98249768611259, 0.98117283193867, 
    0.97977353405102, 0.97839909637378, 0.9768888831075, 0.97568474058862, 
    0.97414437739144, 0.97237477913373, 0.97063708159164, 0.96923524535346, 
    0.96725764301148, 0.96538683208181, 0.96348759190515, 0.96175447420721, 
    0.95955611783301, 0.95721956680606, 0.95492460026066, 0.95253867959545, 
    0.95028368773977, 0.94763225727507, 0.9452100170984, 0.94255770421585, 
    0.93947496614308, 0.93640455091594, 0.93287852345984, 0.93021680578974, 
    0.92667835939391, 0.92290745200672, 0.91941844456351, 0.91536413691863, 
    0.91112917924264, 0.9066382856281, 0.90181974273585, 0.89772537489235, 
    0.89231450443927, 0.8872798235963, 0.88161555489331, 0.87608395339823, 
    0.86980412688855, 0.86302988730412, 0.85590032900328, 0.84797922408935, 
    0.84092161562763, 0.83225575995832, 0.82412885819091, 0.81433397793075, 
    0.8059866950378, 0.79513421700658, 0.78473569504134, 0.77332386534385, 
    0.7607043578912, 0.74732272741939, 0.73425360544451, 0.72061482951629, 
    0.70307644554991, 0.68859199728541, 0.67008043025846, 0.64798055904391, 
    0.62934804528518, 0.60991182158152, 0.58512798309326, 0.5577804655735, 
    0.53147126667643, 0.50701011483097, 0.47726229416586, 0.4474942789931, 
    0.41762443230723, 0.3845020654134, 0.35177143397116, 0.31695038127035, 
    0.28314923418894, 0.24466987162873, 0.20838952060808, 0.17520177705304, 
    0.14250937187759, 0.10996970090122, 0.080190324578789, 0.054938629511495, 
    0.035113673469198, 0.018835514401481, 0.0068331464375787, 
    0.00077953003573895, 0.00069388523552366, 0.0066196262341174, 
    0.016842612360058, 0.033759462662802, 0.055430134900495, 
    0.081167621295699, 0.10976145335141, 0.13855355703304, 0.17471471860712, 
    0.20617971970118, 0.24268211511868, 0.28028110697435, 0.31322223028094, 
    0.34787274779048, 0.37985386016293, 0.41483785527578, 0.44911363715309, 
    0.47973523160962, 0.50488701206668, 0.53415692458494, 0.56054448146036, 
    0.58285041510347, 0.60711420366972, 0.62735054052547, 0.64869441354182, 
    0.6703134541337, 0.68670907479069, 0.70221289511991, 0.71844691728918, 
    0.734778154066, 0.74742444783088, 0.76148767643688, 0.77365259080384, 
    0.78687301568114, 0.79582728365041, 0.80615796588893, 0.81680981834603, 
    0.82478408236124, 0.83422202200782, 0.84240727298304, 0.84915417482157, 
    0.85732081246268, 0.86382930190221, 0.8704775389682, 0.87728426024021, 
    0.8832310391864, 0.88778148671435, 0.8934171256379, 0.89845884074391, 
    0.90396161702709, 0.90807184934745, 0.91201268855079, 0.91619535501481, 
    0.92010413583245, 0.9238212627459, 0.92684035739598, 0.93078708499571, 
    0.93353410328806, 0.93728655238456, 0.93966746310423, 0.94275450224102, 
    0.94523140633156, 0.94806592639122, 0.95027690194856, 0.95280304174195, 
    0.95534623848539, 0.95736092495897, 0.95946235707553, 0.96154004145279, 
    0.96342973945786, 0.96519699055729, 0.96731286979744, 0.96886279286618, 
    0.97052607960793, 0.97217147376592, 0.97372700045353, 0.97530519922658, 
    0.97677879891918, 0.97827921121683, 0.97950251076466, 0.98082382430404, 
    0.98225754938795, 0.98343426556998, 0.98469822673908, 0.98585786382079, 
    0.9869002975985, 0.98805328919114, 0.98917786483287, 0.99023360720808, 
    0.9911773985862, 0.99214616203489, 0.9930928181252, 0.9940079441623, 
    0.99494104115088, 0.99577910858166, 0.99660433202323, 0.99740518095612, 
    0.9982025856585, 0.99892037936158, 0.99963967727633,
  0.99968272668564, 0.9990544247714, 0.99841475157109, 0.997730181659, 
    0.9970390563028, 0.99634896248783, 0.99560434814275, 0.99481796914, 
    0.99403997298652, 0.993273357045, 0.99241145797064, 0.99152877224414, 
    0.99065332364093, 0.98974855003645, 0.98879454608639, 0.98778950927937, 
    0.9867574346528, 0.98562367482475, 0.98462332964501, 0.98348066559019, 
    0.98229768645743, 0.98105486868307, 0.97980426802955, 0.97849182099362, 
    0.9770983088594, 0.97570641280145, 0.97418966421078, 0.97277642302514, 
    0.97118755731379, 0.96952138900207, 0.96779261801226, 0.96614108932158, 
    0.9640564771269, 0.96219574786324, 0.96029950880327, 0.95813057125555, 
    0.95604770594615, 0.95381252707008, 0.95128711432299, 0.94870507945628, 
    0.94615869259291, 0.94343138163383, 0.94067785095822, 0.93786171312109, 
    0.93508709500565, 0.93174675433429, 0.92830494586438, 0.92435592345314, 
    0.92075414924922, 0.91722680322479, 0.91272346902162, 0.90868514257508, 
    0.90344919864238, 0.89965917517188, 0.8947620943462, 0.8887426518082, 
    0.88324875246697, 0.87740626578356, 0.87092475019607, 0.86459681471827, 
    0.85814304173901, 0.85041401961172, 0.8420103391611, 0.83327159333004, 
    0.82415935507677, 0.81508676589198, 0.80562460947469, 0.79403810072478, 
    0.78248744505058, 0.76998649349058, 0.75775921608065, 0.74390702788224, 
    0.72736296831166, 0.71246610743215, 0.69587912039965, 0.67745136453394, 
    0.65845981858779, 0.63751275363463, 0.61531927631877, 0.59060413437283, 
    0.56529140869031, 0.5380654745311, 0.50913364664317, 0.47984720760658, 
    0.44810116635647, 0.41491109814242, 0.37886052418948, 0.34535523289348, 
    0.30729447361021, 0.27059496763721, 0.23233925313957, 0.19399721366565, 
    0.15749113988831, 0.12420138202265, 0.092208551788558, 0.063218594742661, 
    0.039031849847487, 0.020749200436576, 0.0075241863122603, 
    0.00085164254689081, 0.00071264633319524, 0.0075227078915847, 
    0.020729419941756, 0.038140314118752, 0.060810856493205, 
    0.090824062098946, 0.12200556683712, 0.15247562053714, 0.19190197575064, 
    0.22937286401035, 0.26803654858095, 0.3047812923409, 0.3430469780218, 
    0.37706576885255, 0.41506484288889, 0.44661100947583, 0.48114184921538, 
    0.51043742768308, 0.53784598196171, 0.56434994905265, 0.59174271306598, 
    0.61513857914383, 0.63710525415982, 0.65761970317653, 0.67666054690858, 
    0.69581156896159, 0.71253586142287, 0.72954717147341, 0.74404478676077, 
    0.75889752248978, 0.77085367906909, 0.78359611710965, 0.7945669925215, 
    0.80599408746803, 0.81616619162224, 0.82589681612142, 0.83467091743466, 
    0.84222044543707, 0.85086762813545, 0.85907829334508, 0.86582989693601, 
    0.87224701847926, 0.87870304108238, 0.88431391270516, 0.89035551107283, 
    0.89487088847116, 0.90057149053987, 0.90449148149644, 0.90939839040385, 
    0.9137815292757, 0.91757141072494, 0.92132573586749, 0.92528851296783, 
    0.92900949413174, 0.93236385320362, 0.93512876520922, 0.9384366641981, 
    0.94119857263664, 0.94428718167055, 0.94684570089228, 0.94925790432795, 
    0.95133137825002, 0.95376030744561, 0.95632064305272, 0.95811806241738, 
    0.96020581929513, 0.96223721035834, 0.96421665035462, 0.96595941509805, 
    0.96786274463481, 0.96930237001717, 0.97086457219369, 0.97250821714154, 
    0.97405258692663, 0.97554751807255, 0.97674575641106, 0.97826008981602, 
    0.97955031762301, 0.9808331271723, 0.98201813382248, 0.98316784695653, 
    0.98433520709953, 0.98549747734281, 0.98654859772119, 0.98758410927297, 
    0.98847264649999, 0.98957082487012, 0.99048797963629, 0.99137361277201, 
    0.99224492934569, 0.99312721638155, 0.99399477316523, 0.99476889551193, 
    0.9955213012127, 0.99626913687093, 0.99702793391844, 0.99772867665605, 
    0.99839653424836, 0.99905068533938, 0.99968167647304,
  0.99971558608549, 0.99915436119907, 0.99857856174646, 0.99798173425619, 
    0.99736076117431, 0.99672663986431, 0.99607442193134, 0.99539510815158, 
    0.99469424109928, 0.99398503657191, 0.99321853696223, 0.99246902868637, 
    0.99164233656661, 0.99085064971603, 0.99001912158501, 0.98908992777479, 
    0.98817995109626, 0.98726416293486, 0.98629133279769, 0.98524961640222, 
    0.98420347933716, 0.9831278980157, 0.9819513546601, 0.98077050121734, 
    0.97956303088871, 0.97826271367079, 0.97707727232695, 0.97566928880049, 
    0.97409541703022, 0.97275609172032, 0.97126123006454, 0.96961233264894, 
    0.9679195406327, 0.96613121612652, 0.96440624662279, 0.9626001111894, 
    0.96051010751455, 0.95859343621537, 0.9562332904847, 0.95424312003143, 
    0.95153135197625, 0.94934792378559, 0.94673398090202, 0.94421365312681, 
    0.94125608193228, 0.9386024690362, 0.93552950942943, 0.93189963674383, 
    0.9288220533213, 0.9252615867519, 0.92174344778565, 0.91759603651088, 
    0.91341260396884, 0.90894803322584, 0.90411881769235, 0.89973001706162, 
    0.89422525281206, 0.88882434060149, 0.88332586436944, 0.87649326836797, 
    0.8702271160551, 0.86345282353931, 0.85649236559657, 0.84845792479486, 
    0.84124826132701, 0.83135298269031, 0.82166917597557, 0.8118834794951, 
    0.80028255979357, 0.78873670576574, 0.77764489122143, 0.76411922129093, 
    0.75048275094942, 0.73493607046605, 0.71906378216218, 0.70053622622051, 
    0.68083252710329, 0.66171245048813, 0.64130521843869, 0.61677880233456, 
    0.5921782434318, 0.56483350135389, 0.53957275396294, 0.50833750586813, 
    0.47521593349417, 0.442029486483, 0.40578765801567, 0.37025791856619, 
    0.33106969439303, 0.29126305746715, 0.25146308413346, 0.21399720701543, 
    0.17296808502086, 0.13551704056862, 0.10175395730279, 0.069491420765368, 
    0.043729776754901, 0.023037972814613, 0.0082918465805256, 
    0.0010903692591167, 0.00088981285433596, 0.0077539134174045, 
    0.021545700799002, 0.042890854670769, 0.068495760251257, 
    0.099873742878927, 0.13401861527575, 0.17144587426433, 0.21221524745017, 
    0.24931404893767, 0.2897197344767, 0.33098167570147, 0.36895917902531, 
    0.40684866466259, 0.44179418018405, 0.47479848042814, 0.50698370877413, 
    0.53775487258141, 0.56502382598378, 0.59280134995177, 0.61771219669216, 
    0.6393812194953, 0.66316043189543, 0.68339763458167, 0.70068530743749, 
    0.71972527860799, 0.73640999084706, 0.75054577060914, 0.76574820547503, 
    0.77894085554274, 0.7907344727231, 0.80161843573824, 0.81309041591774, 
    0.82269254076402, 0.83224494084134, 0.84143450736199, 0.84984147655724, 
    0.85747476222903, 0.86461589122633, 0.87158129388166, 0.87846642207059, 
    0.88420561457587, 0.89010892184005, 0.89540331167464, 0.90047590932351, 
    0.90531283184126, 0.91008619126488, 0.91434570676755, 0.9184690527053, 
    0.92216242097105, 0.92603993675191, 0.92932851704751, 0.93289208685541, 
    0.93599362021952, 0.93891025267091, 0.94186916577951, 0.94464389277822, 
    0.9473766115598, 0.94962824667703, 0.95191688417663, 0.95431449049932, 
    0.95658475376882, 0.95858274011813, 0.96063656175761, 0.96272532194638, 
    0.9643059556673, 0.96614375969315, 0.96790684132259, 0.96945194426789, 
    0.97100327030136, 0.9726179268747, 0.9740402622318, 0.97544435692917, 
    0.97671860132667, 0.97815509851768, 0.97932918544745, 0.9805629700303, 
    0.98171602280216, 0.98286213355886, 0.9839740422829, 0.98501512721598, 
    0.98598499571368, 0.98702686846572, 0.98802307209563, 0.98891873384868, 
    0.98978838914885, 0.99067824483385, 0.99150986551991, 0.99232768734997, 
    0.99311576510865, 0.99387610580222, 0.99461416970093, 0.99533936140189, 
    0.99602399205219, 0.99669553704176, 0.99733693005339, 0.99796746214299, 
    0.99856696392471, 0.99915370220315, 0.99971490181441,
  0.99974216625611, 0.99923531727051, 0.99871458948366, 0.99817074232315, 
    0.99761443879884, 0.9970407053136, 0.99645238873888, 0.99583440268011, 
    0.99523381044764, 0.99453316450399, 0.99389078823398, 0.99319022925108, 
    0.99248580984241, 0.9917365828139, 0.99095147531122, 0.99016473137999, 
    0.98932508252921, 0.98852024665376, 0.98758411380224, 0.98668292114839, 
    0.98573202241504, 0.9847955072277, 0.98370103479914, 0.98263772311779, 
    0.98155904085663, 0.98037425003285, 0.97922713718623, 0.97788617063476, 
    0.97666778099303, 0.97546949330564, 0.97395269572127, 0.97250422198259, 
    0.97114520692878, 0.96938385262249, 0.96776733657306, 0.96600746999039, 
    0.96435152473168, 0.96239735990684, 0.96041576859332, 0.95847668492905, 
    0.95644667405053, 0.95400878308521, 0.95178754212928, 0.94924247435284, 
    0.94683451756254, 0.94424740971438, 0.9410965648947, 0.938315956195, 
    0.93523880205842, 0.93210880785815, 0.92856819296449, 0.92459730953142, 
    0.92088298661883, 0.91708025646045, 0.91256501130046, 0.90856894847646, 
    0.90360597667364, 0.89834875084141, 0.89316308426066, 0.88727322861578, 
    0.88107989441388, 0.87473719928352, 0.86875761429464, 0.86094894874489, 
    0.85334832463982, 0.84463519863813, 0.83579665648983, 0.82612754086566, 
    0.81600449527093, 0.80564163323966, 0.79431754664012, 0.78136430235161, 
    0.76688103559802, 0.75322539150788, 0.73859017736142, 0.72102920328853, 
    0.7030552117294, 0.68359010130883, 0.66337850381609, 0.64018105269131, 
    0.6159405505236, 0.59001349827187, 0.56335147158681, 0.53158189255681, 
    0.50075282136098, 0.46497003568166, 0.43031750288383, 0.39195627764367, 
    0.35353197173248, 0.31105856132577, 0.27214983193249, 0.22809826149769, 
    0.18823188213557, 0.14767377704639, 0.11105214983583, 0.078366475023877, 
    0.047711581497996, 0.024677161063393, 0.0093486830850011, 
    0.0011836153103796, 0.00093680124817239, 0.0085327772229286, 
    0.02461066381764, 0.047458645970744, 0.076558052941852, 0.10878573544953, 
    0.14568273545796, 0.18680609440963, 0.22843352280143, 0.26756624799846, 
    0.31198638209064, 0.3513064688807, 0.39153598695651, 0.42898682541974, 
    0.4667295701282, 0.50049044565351, 0.53301574396231, 0.56177912873701, 
    0.59203462591823, 0.61684174247875, 0.6413662789757, 0.66405679932453, 
    0.68539343531605, 0.70457607461302, 0.72128232780807, 0.73917958429018, 
    0.75477420825215, 0.76998621990474, 0.78299862325651, 0.79520998843105, 
    0.80685754372158, 0.817830693427, 0.82798652547854, 0.83752285218666, 
    0.8457641430113, 0.85435245997312, 0.86276798897957, 0.86861006930269, 
    0.87620879048143, 0.88285038122607, 0.88871346061979, 0.89442557730117, 
    0.89952285420357, 0.90476949239499, 0.90899794356986, 0.91360477581686, 
    0.91790709284643, 0.92214511618945, 0.92581328765878, 0.92907791232901, 
    0.93268618123944, 0.93585625517925, 0.93871519493689, 0.94181284726634, 
    0.94463314833387, 0.94731761894341, 0.94964303719067, 0.95188326004527, 
    0.95431194820685, 0.9565172720171, 0.95860071493363, 0.96059104259049, 
    0.9625003433715, 0.96429486567337, 0.96607188619815, 0.96772278967958, 
    0.96925294885993, 0.97097247303441, 0.97231611969769, 0.97388070286602, 
    0.97520316853643, 0.97649727551881, 0.97777828628628, 0.97900920067829, 
    0.98018877606237, 0.98132073063612, 0.982435846566, 0.98349517928279, 
    0.98446512009489, 0.98552461647948, 0.98649676248062, 0.98734036482696, 
    0.98835815853205, 0.98910194865578, 0.98997248466391, 0.99082547090076, 
    0.99158856701641, 0.99233822812855, 0.99309282874553, 0.99379778182296, 
    0.99447026087354, 0.99515073071659, 0.99579273079583, 0.99641446274723, 
    0.99701438512839, 0.99759637515912, 0.99815924117954, 0.9987065609725, 
    0.99923248861109, 0.99974136848983,
  0.99974883359838, 0.9992537728586, 0.99873974775466, 0.99822015837811, 
    0.99767009923872, 0.99711148874292, 0.99654351723571, 0.99592846081254, 
    0.99533373770449, 0.99468595851056, 0.99402621749447, 0.99336342830235, 
    0.9926579754098, 0.99192012024112, 0.99116154017795, 0.99039354310225, 
    0.9896167160694, 0.98875887738515, 0.98785111045796, 0.98703356065746, 
    0.98608130705655, 0.98513090835481, 0.98414274965258, 0.98307704240276, 
    0.98194435989023, 0.98086591724137, 0.97972108779921, 0.97845143789233, 
    0.97723292522708, 0.97592445552499, 0.9745201991993, 0.97313968082301, 
    0.9716765844017, 0.97022704798529, 0.96851390477879, 0.96684702173259, 
    0.96514333484946, 0.96327057712223, 0.96133041051987, 0.9594184794978, 
    0.95727577156861, 0.95501620215107, 0.95300511919625, 0.95043351728872, 
    0.94800605813513, 0.94534478661997, 0.94262717652792, 0.93957947623308, 
    0.93674257804322, 0.9333797380989, 0.93001764417993, 0.92653496571909, 
    0.92306286821364, 0.91878422598184, 0.91455511192005, 0.91028464517762, 
    0.90547557373004, 0.90054431654078, 0.8954657725302, 0.8893898706366, 
    0.88403235594305, 0.87769133572321, 0.87096445100114, 0.86336642741651, 
    0.85594567819113, 0.84783696889805, 0.83921885315349, 0.83029132278923, 
    0.81942644555185, 0.80926574954158, 0.79772374063539, 0.78531838809649, 
    0.77132163876172, 0.75729790931278, 0.74242344043379, 0.7261801880777, 
    0.707817700407, 0.68810144262355, 0.66924052877231, 0.64428590865626, 
    0.62152592305048, 0.59657431504241, 0.56762441183089, 0.53745025619006, 
    0.50572628210719, 0.47207259449938, 0.43713743856525, 0.39770476876339, 
    0.35947905107168, 0.31750881350563, 0.27400257640089, 0.23380509691542, 
    0.19152969588626, 0.15211887985323, 0.11224677082718, 0.078850949099042, 
    0.047830358244159, 0.026063507829444, 0.0096228154630117, 
    0.0011787942695495, 0.00098387210393263, 0.008749814499432, 
    0.025236581540318, 0.047824563971794, 0.078704063828795, 
    0.11186938995683, 0.14779502497071, 0.18991402471717, 0.23299623092229, 
    0.27344925084194, 0.31728882817944, 0.35895796719972, 0.39671697330018, 
    0.43602834141191, 0.47247823645058, 0.50666967893999, 0.53882901643089, 
    0.56708341632869, 0.59677416702509, 0.62146665522954, 0.6465473058004, 
    0.66870448221164, 0.69056974379027, 0.70957525873561, 0.72706555132606, 
    0.74360923454207, 0.75919450598219, 0.7735203122787, 0.78663811526685, 
    0.79883204492584, 0.81069822929635, 0.82154065352963, 0.83128929587337, 
    0.84069399897527, 0.84913517590621, 0.85765985860512, 0.86526709895877, 
    0.87194754476904, 0.87874655921246, 0.88514996530674, 0.89100401585273, 
    0.8963744268697, 0.90172069369269, 0.90652840014772, 0.91124248487664, 
    0.91553312173042, 0.91980018598246, 0.92360087782221, 0.92733259021448, 
    0.9305803344776, 0.934244975327, 0.937087204596, 0.94013817378087, 
    0.94305940862646, 0.94576779400343, 0.94838349632973, 0.95070171764279, 
    0.9532707016228, 0.95530509045926, 0.95737557282101, 0.95956575729418, 
    0.96157879219502, 0.96331477744154, 0.96505014736914, 0.9668758926266, 
    0.96847558681034, 0.9699672919058, 0.97151832446219, 0.97313513221931, 
    0.97438178307043, 0.97571999086751, 0.97702233529187, 0.97831014968332, 
    0.97948645087937, 0.9806392133322, 0.98178711111852, 0.98281808174659, 
    0.98390296978061, 0.984914369963, 0.98583903899874, 0.98678771349705, 
    0.98767122178995, 0.98854420444656, 0.98944067885649, 0.99020718856075, 
    0.99101075084374, 0.99178652745481, 0.99253977450209, 0.99324481462635, 
    0.99395569222272, 0.99461164529979, 0.99525616244461, 0.99588727193165, 
    0.99649952364516, 0.99708628761842, 0.99765648902285, 0.99820517207034, 
    0.99873386812579, 0.99925154198096, 0.99974743776011,
  0.9997534646866, 0.99926961014293, 0.99877091532912, 0.99825548470533, 
    0.9977235635145, 0.99718163085466, 0.99660374014661, 0.99603931077835, 
    0.99543099213711, 0.99480569335371, 0.99417299490437, 0.99352899210962, 
    0.9928108652675, 0.99210740342489, 0.99140041096478, 0.99060665283775, 
    0.98981805486239, 0.98901191118424, 0.98818811006606, 0.98731108712346, 
    0.98640925329091, 0.98543251489257, 0.98450786106851, 0.98345110764819, 
    0.98243930393519, 0.98128284887961, 0.98019448095793, 0.97897037519407, 
    0.97772242503668, 0.97649221854835, 0.97518103868065, 0.97370385743309, 
    0.97233416179963, 0.97076049532802, 0.96931572406444, 0.96756825398155, 
    0.96588009650819, 0.96407813907102, 0.96232834322263, 0.96025240014655, 
    0.95820475581917, 0.95610016306759, 0.95388258032001, 0.95161946604437, 
    0.94909997522737, 0.94652421034558, 0.94377614840787, 0.94105893276463, 
    0.93790534785593, 0.93491027925856, 0.93160677113528, 0.92816028465348, 
    0.92427165416634, 0.92052848637568, 0.91670109557876, 0.91171131064516, 
    0.9073747955975, 0.90284639107006, 0.89754050804506, 0.89205072076177, 
    0.88579606637141, 0.87996816742047, 0.87361931631983, 0.8661648688098, 
    0.85919794882245, 0.85004252724625, 0.84235698053263, 0.83280647552997, 
    0.82309311721815, 0.81202543125171, 0.80158453893801, 0.78974755705626, 
    0.77541879072721, 0.76202740725546, 0.74676563239682, 0.7305863622959, 
    0.71160674657048, 0.69297010210833, 0.67343010079779, 0.65152419598741, 
    0.62720152385367, 0.60061168451328, 0.57311541980679, 0.54445073013479, 
    0.51058708948718, 0.47658333282346, 0.44147223876315, 0.40416677758253, 
    0.36293609292231, 0.32438966589552, 0.28028868509801, 0.23694465662414, 
    0.19501512554723, 0.15333060253939, 0.11547643905433, 0.080137952122812, 
    0.050172920210336, 0.02639229378429, 0.0098193094127902, 
    0.0011275192922408, 0.00098874638264249, 0.0087572741030965, 
    0.026271818771934, 0.049282092071127, 0.078698271974419, 
    0.11282701910047, 0.15248131042449, 0.19428802145538, 0.23519836539696, 
    0.27930895090834, 0.32104810707886, 0.36436559312027, 0.40475007021224, 
    0.44079362999862, 0.47803586970848, 0.51234905379303, 0.54353629637618, 
    0.57420406372253, 0.60130178468935, 0.62814089644551, 0.65236821482529, 
    0.67511514840501, 0.69463157180776, 0.71316452168099, 0.73217011096269, 
    0.74761350993323, 0.76359670636398, 0.77709979707666, 0.79118547440438, 
    0.80292421590614, 0.81391833216552, 0.8245355564463, 0.83466658227963, 
    0.84331795094377, 0.85206218434348, 0.8602990683839, 0.86773823639517, 
    0.8750897191299, 0.88130633094781, 0.88787310365246, 0.89308932979266, 
    0.89850411661698, 0.9034161892371, 0.90884135861804, 0.91319072715895, 
    0.91736489183897, 0.92128530661376, 0.92497644033119, 0.92884479799444, 
    0.93218093031752, 0.93555022170679, 0.93853849952635, 0.94158882786154, 
    0.94410574358744, 0.94687941571691, 0.94957533056343, 0.95192633387443, 
    0.9542511418781, 0.95628462194767, 0.95854844630995, 0.96026903001436, 
    0.96248793629705, 0.96417293571937, 0.96582522186298, 0.96763064034837, 
    0.96916111833473, 0.97067416073815, 0.97221413364267, 0.97361649490977, 
    0.97496760591496, 0.97629557431787, 0.97757296008665, 0.97880800134109, 
    0.97997378935319, 0.98109579879282, 0.98215562017865, 0.98323991856471, 
    0.98425205827174, 0.98524836984224, 0.98617128705384, 0.98712205356872, 
    0.98795322456524, 0.98881866681605, 0.9896723894711, 0.99044821990688, 
    0.99123874929388, 0.99198613083252, 0.99269182993449, 0.99340150047981, 
    0.99409726928421, 0.99472901314629, 0.99537828648909, 0.99598306545866, 
    0.99657859002545, 0.99716021704801, 0.99770459269561, 0.99824726219284, 
    0.99876501716148, 0.99926740218978, 0.99975262221121,
  0.99976347936473, 0.99930160573638, 0.99882227746305, 0.99833392663197, 
    0.99782196913991, 0.99730033058004, 0.99675816863603, 0.9961993053481, 
    0.99563088003974, 0.99504425140512, 0.99441369005225, 0.99379011592718, 
    0.99313372589009, 0.99246589952475, 0.9917727835765, 0.99101081241979, 
    0.99027494124779, 0.9895242881879, 0.98867355280538, 0.98785391465771, 
    0.98700486830027, 0.98613343691637, 0.98510520128815, 0.98411527214862, 
    0.98320782222607, 0.9821566598921, 0.98108459165987, 0.97992467332788, 
    0.9787498840467, 0.97748798054929, 0.9762197902326, 0.974909586339, 
    0.97339592187504, 0.97213172712459, 0.97050349879944, 0.96908146518063, 
    0.96729070953737, 0.96570757034753, 0.96388467733381, 0.96187433381787, 
    0.96008554781679, 0.95805591299438, 0.95583300656103, 0.95357661883533, 
    0.95124185907739, 0.94895068015068, 0.94627550859975, 0.94341440788694, 
    0.9407692426476, 0.93733812520901, 0.93438260298466, 0.9308004379668, 
    0.92764561343652, 0.9237851921464, 0.91988517276494, 0.91566402377613, 
    0.91087538610954, 0.90642653785616, 0.90151626725264, 0.89631140896374, 
    0.89060294458352, 0.88455584415516, 0.87829310569327, 0.87133263633593, 
    0.86365102446232, 0.85662252155937, 0.84865793651053, 0.83845272120012, 
    0.82913435742164, 0.81915520240408, 0.80714693414907, 0.79631674702914, 
    0.78367416651302, 0.76980637069865, 0.75467965145226, 0.73940843928058, 
    0.72170094971317, 0.70279379921411, 0.68270826073081, 0.65927616370809, 
    0.63602502151172, 0.61213320480324, 0.58388217189055, 0.55344041286628, 
    0.52269157585436, 0.49017983829144, 0.45248155818071, 0.41317899185777, 
    0.37288962122627, 0.33019757370753, 0.29042190635144, 0.24610379573324, 
    0.20237267296819, 0.15814932817245, 0.12040786690859, 0.083192711753062, 
    0.052401769682276, 0.027529248179231, 0.010609607306022, 
    0.0012125016865987, 0.0010356007889027, 0.0097718843771333, 
    0.026474993681497, 0.052203230298746, 0.081766176356332, 
    0.11705140602614, 0.15878506967828, 0.20207607555962, 0.24456489061522, 
    0.28678217219346, 0.33203691200751, 0.37310499694638, 0.41436971144161, 
    0.451923687499, 0.48928666562035, 0.52307120637413, 0.55458566431612, 
    0.58561131874038, 0.61391040649274, 0.6387358620243, 0.66311214488532, 
    0.68337029908993, 0.70352624148998, 0.7232188684294, 0.73933211840573, 
    0.75633568953946, 0.7714430072014, 0.78547614432185, 0.79758422663138, 
    0.80959403571385, 0.82049669285907, 0.83077127726573, 0.84167861465519, 
    0.84936296890096, 0.85799214577384, 0.86563066501643, 0.87261039928026, 
    0.87954503505704, 0.88582081629868, 0.89134950785556, 0.89711653192042, 
    0.90301997747512, 0.90773414377911, 0.91211209372244, 0.91626468963177, 
    0.92069788677689, 0.92453175027171, 0.92836108648162, 0.93178486825206, 
    0.93515125357857, 0.93832059805402, 0.94108934430451, 0.943980320859, 
    0.94655504388343, 0.94916845988099, 0.95153076217786, 0.95387709295335, 
    0.95601346661437, 0.95819434374877, 0.96008907615407, 0.96213413207282, 
    0.96389116380908, 0.96573910781485, 0.9673501471314, 0.96893142429818, 
    0.97051083681744, 0.97196983745482, 0.97332798801934, 0.97480369162947, 
    0.97610578008243, 0.9773499416506, 0.97851028936722, 0.97971938411585, 
    0.98084547266015, 0.98193506177802, 0.98294494679735, 0.98402850429421, 
    0.98497255209617, 0.98585732821927, 0.98678160730498, 0.98765271055444, 
    0.98851308586684, 0.98930465356441, 0.9901209177161, 0.99087820654831, 
    0.99162517192854, 0.99234920429212, 0.99304344934037, 0.99369311479319, 
    0.99434402524457, 0.99497630783801, 0.99558050410267, 0.99616016438718, 
    0.99672939579448, 0.99728107305665, 0.99781500558152, 0.99832145899824, 
    0.99882059527585, 0.99929828649063, 0.99976321213942,
  0.99978148981376, 0.99935543448604, 0.99891658583945, 0.99846367605554, 
    0.99800022124965, 0.99751110058465, 0.9970217738499, 0.99650377469683, 
    0.99598139258273, 0.99543935375106, 0.99487123874995, 0.99430668493449, 
    0.9936666062772, 0.99306223721288, 0.99239447701865, 0.99176697506467, 
    0.99109276003938, 0.99035955072014, 0.98958986295437, 0.98882104898754, 
    0.98802881184707, 0.98722226990249, 0.98634517341952, 0.98545381445099, 
    0.98460271284547, 0.98351495606787, 0.98259102878617, 0.9815696149963, 
    0.98037870183668, 0.97929510476445, 0.97811374990617, 0.976876436594, 
    0.97563679619742, 0.97426832740929, 0.97295888675709, 0.97132415535823, 
    0.97001712498802, 0.96834860720555, 0.96656456909489, 0.96501886129431, 
    0.96311545439489, 0.96136049294159, 0.9591876510344, 0.95721506434485, 
    0.95500796844222, 0.95279059090559, 0.95043266891918, 0.94770919661397, 
    0.94510060976552, 0.94241784487264, 0.93936056972373, 0.93613300542344, 
    0.93290874170144, 0.92951551732186, 0.92582841600829, 0.92181563556813, 
    0.9179617250323, 0.91295794425875, 0.90896656605697, 0.90336489561511, 
    0.89824870069398, 0.89273044750879, 0.88675091734827, 0.88030606184763, 
    0.87353048835989, 0.86626162373622, 0.85812895825486, 0.84970024716781, 
    0.84141908969765, 0.83096621353146, 0.82015949644935, 0.8090237480149, 
    0.79755515064215, 0.78380463977046, 0.76963462331877, 0.75398568405714, 
    0.73818444655135, 0.72059702516851, 0.6989859195142, 0.6791928791983, 
    0.65472186002797, 0.63174930636667, 0.60351373598342, 0.5738663367892, 
    0.54229715386342, 0.50944028203828, 0.47346943713838, 0.43466400993846, 
    0.39184508836552, 0.35110923702426, 0.30629026185446, 0.26068519826713, 
    0.21397632540156, 0.17149921614142, 0.12729641446638, 0.089810428545838, 
    0.056598179733238, 0.029910129306845, 0.011282953162232, 
    0.0012953315239348, 0.0010629380872959, 0.011158344863007, 
    0.028242003108943, 0.05618820177145, 0.089704258113067, 0.12635952521038, 
    0.17110324668561, 0.21359784199117, 0.25939572363947, 0.30627047153913, 
    0.35051436523833, 0.39359700950473, 0.43381182624105, 0.47282707658962, 
    0.51159365883411, 0.54298090790922, 0.57654327307881, 0.60522985063996, 
    0.6318843861562, 0.65756316852204, 0.68149265241673, 0.70130183983125, 
    0.72149119743781, 0.73977946647198, 0.75651276686259, 0.77140008872203, 
    0.78544874404331, 0.7987330221105, 0.81058354469416, 0.82194552616455, 
    0.83296408980934, 0.84282682436359, 0.85147373802854, 0.85980894207606, 
    0.86745188897007, 0.87466126440119, 0.88172433971915, 0.88820737251785, 
    0.89374788388879, 0.89976982720107, 0.90485960485925, 0.90973591278858, 
    0.91440515724331, 0.91856624531353, 0.9225177491621, 0.92662442912567, 
    0.93011311066342, 0.93365391627248, 0.93695805097444, 0.94000286241225, 
    0.9428329888852, 0.94557528189673, 0.94825454146438, 0.95057159339032, 
    0.95293663722408, 0.95530624296128, 0.95731793778742, 0.95956353502135, 
    0.96130515215373, 0.96331499920708, 0.96496113074225, 0.96667271019877, 
    0.96845320012705, 0.96992746462248, 0.97147175066396, 0.9727982713505, 
    0.97422584510371, 0.97549797253376, 0.97675101631163, 0.97802676236228, 
    0.97910662351542, 0.98023318297669, 0.98136021870068, 0.98246264897017, 
    0.98340439052794, 0.98434751952406, 0.98530665956359, 0.9861320552427, 
    0.9870436930097, 0.98786063019248, 0.98869017930853, 0.98945390049207, 
    0.99021348818825, 0.99092422497659, 0.99163808315059, 0.99231624390322, 
    0.99298129921577, 0.99360528051198, 0.99420093162821, 0.99481191388312, 
    0.9953725499277, 0.9959453845888, 0.99648106776327, 0.99699511740004, 
    0.99749682642218, 0.99798914363481, 0.99846045505642, 0.99891403692071, 
    0.99935577033135, 0.99978142141754,
  0.99979778344139, 0.99940611992618, 0.99899996165692, 0.99857133045752, 
    0.99814853804508, 0.99770590916041, 0.99725651889184, 0.99677950552035, 
    0.9962965377177, 0.99573365734292, 0.99523894386481, 0.99474454339588, 
    0.99414315723181, 0.99358040109227, 0.99293810297096, 0.99232849697893, 
    0.99171508950288, 0.99111425213036, 0.99037880702133, 0.98968233818842, 
    0.98883687687874, 0.98809838593129, 0.98739452152578, 0.98660239722557, 
    0.98579431289356, 0.98483378905171, 0.98377108104402, 0.98277080220374, 
    0.98187575138477, 0.98085969504396, 0.97980493231576, 0.97875751569579, 
    0.97734041491475, 0.97619869737853, 0.97510000012623, 0.97367452317009, 
    0.97215727931499, 0.97061297420454, 0.96908753903252, 0.96754212769465, 
    0.96573051627644, 0.96403707340879, 0.96213108784606, 0.95985857212283, 
    0.95809445760117, 0.95599180703572, 0.95391125409222, 0.95140195961987, 
    0.94908460003136, 0.94678100869554, 0.94358971444684, 0.94070452656873, 
    0.93765882726717, 0.93444525639905, 0.93098167429729, 0.92744157117485, 
    0.92377493548492, 0.91930456950798, 0.91429351725966, 0.90999479454967, 
    0.90548544672797, 0.89969489280121, 0.894560776011, 0.88919961072685, 
    0.88133999609159, 0.8743964261206, 0.86591617018775, 0.85939159498742, 
    0.85043279702591, 0.84191740583746, 0.83104334581472, 0.82041078431852, 
    0.80774887027591, 0.79654252298773, 0.78359736805847, 0.77006923174408, 
    0.75368374664188, 0.7352557578316, 0.71536553507616, 0.69315155333355, 
    0.6715943701673, 0.65080079152746, 0.62327188523518, 0.59423008316313, 
    0.5596008798758, 0.52693016529377, 0.49137456190756, 0.45201373942669, 
    0.41169960536842, 0.36562649075595, 0.32145840539423, 0.27196786595155, 
    0.22704393510794, 0.18311195830871, 0.14064163021309, 0.095223247396541, 
    0.060242561289561, 0.030711035366732, 0.011023454809568, 
    0.0015356497896226, 0.00097402099884918, 0.010283175390779, 
    0.029777153171709, 0.06059463699015, 0.096024073122303, 0.13551036798915, 
    0.18255306938446, 0.23008876880837, 0.27281250818438, 0.32207900400039, 
    0.36443702222455, 0.41185884927143, 0.45676289237438, 0.49307925938354, 
    0.5298653672634, 0.56539852658548, 0.59483161085507, 0.62298132110322, 
    0.64929393509525, 0.67542309602135, 0.69668709723969, 0.71830825686921, 
    0.73453136059621, 0.75358878488591, 0.77200941061925, 0.78621502477201, 
    0.79860789437782, 0.80904138025086, 0.82120185702988, 0.83278985007337, 
    0.84327802489913, 0.85318601201125, 0.86209688834125, 0.86873426895679, 
    0.87562823005542, 0.88234280520669, 0.88914528345902, 0.89579219014869, 
    0.90210551298797, 0.90647114508295, 0.91110051794038, 0.9156578141566, 
    0.92004000785012, 0.92407560519286, 0.92787526169167, 0.93167631699499, 
    0.9350164560889, 0.93827140977291, 0.941579798561, 0.94399887500048, 
    0.94691852297944, 0.94959189968627, 0.95151238932205, 0.9543756009783, 
    0.95672388305334, 0.95834006057666, 0.9602447989723, 0.96229696098297, 
    0.9644463045941, 0.9659929216505, 0.96760168372875, 0.96895227872347, 
    0.97055171187424, 0.97204545336052, 0.97351329873886, 0.9748278614226, 
    0.97616346239557, 0.97734359936639, 0.97847829904872, 0.97973999169766, 
    0.9806409879277, 0.98167668469523, 0.98276611959845, 0.98359994518774, 
    0.98470840795862, 0.98552593656841, 0.98641834860865, 0.98721045604908, 
    0.98799966404294, 0.98876077375637, 0.98953715519178, 0.99027270504553, 
    0.99095087768127, 0.99167535677673, 0.99234095336421, 0.99288631090091, 
    0.99347881967955, 0.99405531056019, 0.99469192575997, 0.99520113898243, 
    0.99573465711728, 0.99625822003047, 0.99673113376571, 0.99722018133532, 
    0.99770137611419, 0.99814345401965, 0.99856542440267, 0.9989910766949, 
    0.99940394987128, 0.99979823104967,
  0.99981105216474, 0.99944536330554, 0.999066648429, 0.99867845026012, 
    0.99827588846322, 0.99786295053878, 0.99743718498022, 0.99699683053934, 
    0.9965364992812, 0.99607449852978, 0.99559043351659, 0.99507639023151, 
    0.99456668704205, 0.99402959972065, 0.99348233054668, 0.99289619176256, 
    0.99230154805173, 0.99170415842651, 0.99103599244633, 0.99037181681877, 
    0.98970900103442, 0.98900405396754, 0.98822345600126, 0.98748093075023, 
    0.9866499602495, 0.9858319579026, 0.98499162798721, 0.98405553767269, 
    0.98313867851203, 0.98214262162779, 0.98113431250715, 0.98003133599135, 
    0.97900043145042, 0.97787643491356, 0.97655940435676, 0.97532377414895, 
    0.97402792315634, 0.97261803647322, 0.97122384052071, 0.96974894282952, 
    0.96814127958565, 0.96642616626225, 0.9648137523772, 0.96298100815724, 
    0.96098464108766, 0.95905455323035, 0.95703214666633, 0.95471518429388, 
    0.95236227497411, 0.94992406089361, 0.94734586300586, 0.94446373095166, 
    0.94179688618739, 0.9385986963261, 0.93528494400529, 0.93189939768391, 
    0.92811923310357, 0.92441943420329, 0.92015361597955, 0.915688948851, 
    0.9112214140892, 0.90625028931304, 0.9006299588865, 0.89496008536656, 
    0.88865101958825, 0.88242284254746, 0.87540211925303, 0.86801638714339, 
    0.85931605522387, 0.8506689040391, 0.84135714747375, 0.83064398861385, 
    0.81998137276424, 0.80726152754581, 0.79392694220957, 0.78061739582751, 
    0.76517124909661, 0.74846562845681, 0.73052143682496, 0.70958907177604, 
    0.68836015434184, 0.66403266465334, 0.63776910652253, 0.61029308136073, 
    0.57838575028834, 0.54555393568384, 0.50983868067049, 0.46976890864823, 
    0.42827014708581, 0.38568448845021, 0.33821449885269, 0.29118226643733, 
    0.24118809291034, 0.19273699458439, 0.14522267557303, 0.10216284730577, 
    0.0654470450535, 0.034063088122067, 0.012589763724512, 
    0.0016264004253476, 0.0013363783798251, 0.012562630348383, 
    0.033605190742324, 0.064153583423394, 0.10182480286432, 0.14377378812771, 
    0.19145958067355, 0.24079125977721, 0.29001234813848, 0.33782614562491, 
    0.38368693893453, 0.43004153544798, 0.47187120920719, 0.51113726946344, 
    0.54742860366802, 0.58067478263151, 0.61044996402185, 0.64083511858854, 
    0.6658317878512, 0.68974449799536, 0.71194909704324, 0.73164452960089, 
    0.75098557665944, 0.76730069928615, 0.78212001195434, 0.79674556472609, 
    0.80923314033673, 0.82157743969816, 0.83312775518648, 0.84276993838863, 
    0.8523394523393, 0.86153321325558, 0.86946522613941, 0.87685264401522, 
    0.8835627914768, 0.89020618112306, 0.89634924694087, 0.90214054885067, 
    0.9075070536575, 0.91210061471743, 0.9165541052991, 0.92120882098009, 
    0.92512332969154, 0.92909081298443, 0.93270127871053, 0.93604442597474, 
    0.93949324282846, 0.94238991297856, 0.94511357565413, 0.94784466955843, 
    0.95013373638648, 0.95293361636051, 0.95504807884407, 0.95735878644941, 
    0.95930535027152, 0.96118039231914, 0.9632589158742, 0.96504539981828, 
    0.96652382540148, 0.96832776103822, 0.96980741751693, 0.97132086853613, 
    0.97271769412352, 0.97400659960458, 0.97530706682769, 0.97661713218465, 
    0.97775024264086, 0.97890304927165, 0.97999459083882, 0.98106869899259, 
    0.98204878859398, 0.98303344165585, 0.98396161099865, 0.98479287833185, 
    0.98573701495478, 0.98656611559046, 0.98732965889024, 0.98812859559994, 
    0.98884645026196, 0.98957357758711, 0.99028245263179, 0.99095338885307, 
    0.99160569010181, 0.99220115899596, 0.99280743593912, 0.99339478039504, 
    0.99396038860326, 0.99450705239708, 0.99502112232945, 0.99554289891155, 
    0.99603677151352, 0.99650645928042, 0.99697481677424, 0.99741938076547, 
    0.99784781373342, 0.99827103685992, 0.99867401287937, 0.99906399477031, 
    0.99944417641202, 0.99981084564411,
  0.99982796410243, 0.99949655013457, 0.99915391873637, 0.99880376598456, 
    0.99844135337217, 0.99806659170544, 0.99767677919292, 0.99728811039772, 
    0.99686379082557, 0.9964428858673, 0.9960023852605, 0.99554737200602, 
    0.99509926896104, 0.99458976174077, 0.99409630775974, 0.99355253236735, 
    0.99304518510557, 0.9924732146761, 0.99189715366907, 0.99128858394701, 
    0.99068010106865, 0.99002018344099, 0.98934118256772, 0.98863033079011, 
    0.98793289596961, 0.98713573709572, 0.98636603144757, 0.98557962395812, 
    0.98469672792833, 0.98381735662778, 0.98288563111172, 0.98194327514607, 
    0.98089503204082, 0.97984829655933, 0.97874145450512, 0.97762537152161, 
    0.97643794001034, 0.97509831822878, 0.9738393960982, 0.97255178087805, 
    0.97107045541634, 0.96958082189919, 0.96790221496197, 0.9663730688694, 
    0.96445190183123, 0.96281566976894, 0.96083325435935, 0.95876451315773, 
    0.95647911067896, 0.9544423289279, 0.95200617001843, 0.94957004132093, 
    0.94679619419454, 0.9441520132303, 0.94095297845575, 0.93775249603767, 
    0.93444858350518, 0.93095799307114, 0.92713707886318, 0.92317671254283, 
    0.91882146375844, 0.91405698823337, 0.90936440362773, 0.90364997213795, 
    0.89831852952047, 0.89159473703648, 0.88583763304256, 0.87881623484329, 
    0.87056430811498, 0.86324436743786, 0.85430205440076, 0.84400448100176, 
    0.83402165131141, 0.82212732171837, 0.81012658687002, 0.79671105041153, 
    0.78251017496378, 0.76587095158713, 0.74841733224497, 0.72960942431689, 
    0.70911488505426, 0.68530797992955, 0.66084200966205, 0.63381251151494, 
    0.60292258536771, 0.56874405340933, 0.53441477655025, 0.4944345656981, 
    0.45234148913434, 0.4063590389123, 0.36069222630265, 0.31097997789308, 
    0.25948265634113, 0.20679396827843, 0.16057322082352, 0.11144036810061, 
    0.070375143442519, 0.037674266404307, 0.013944001958685, 
    0.0015798859822841, 0.0014847394297306, 0.013364182007257, 
    0.036327329284, 0.069923300057189, 0.11124891279911, 0.15795441989848, 
    0.20686826925635, 0.26013850969734, 0.31100104558304, 0.36084028835631, 
    0.40542790695634, 0.45477725181284, 0.49666563571962, 0.53448589158186, 
    0.57226937192164, 0.60319773775086, 0.63368404858753, 0.66289994328107, 
    0.68667485576169, 0.71010435227316, 0.73175996386915, 0.75099408734676, 
    0.76819595960532, 0.78438616241861, 0.79820516332347, 0.81243632158776, 
    0.82435950773131, 0.83539659765544, 0.8458562930391, 0.85537196571597, 
    0.8641480311318, 0.87261685974321, 0.88041960788869, 0.88706455013621, 
    0.8936927747234, 0.8993200743566, 0.90512388520085, 0.91051763802344, 
    0.91506250881353, 0.91988781255718, 0.92422754311361, 0.92816051041598, 
    0.93167421280552, 0.93531108024274, 0.93876874203097, 0.94173835435577, 
    0.94480759733435, 0.94728977843933, 0.94999163437538, 0.95240896023988, 
    0.95482080294578, 0.95706891781876, 0.95916371006606, 0.96111545661712, 
    0.96295599128091, 0.96496247804109, 0.96652465982791, 0.96817156231279, 
    0.96973420623086, 0.97115529019806, 0.97258197763854, 0.97392426787467, 
    0.97514361454081, 0.97647973457598, 0.97764507001208, 0.97873824337163, 
    0.97986878058411, 0.98091898070856, 0.98186610315807, 0.98278473933803, 
    0.98370954224973, 0.98462366190927, 0.98547897790016, 0.98630158571533, 
    0.98704070429363, 0.98783265215939, 0.98851500071536, 0.98927343762508, 
    0.9898963735303, 0.99058952361969, 0.99117190356345, 0.99177792616896, 
    0.99240248768682, 0.99295709270257, 0.99350776699655, 0.99401243343951, 
    0.9945200121842, 0.99503688052034, 0.99549334945456, 0.99597013189807, 
    0.99640595144254, 0.99684066623013, 0.99726240131863, 0.99766424844514, 
    0.99804995007394, 0.99843709687162, 0.99879780882351, 0.99915406059052, 
    0.99949571769234, 0.99982782443078,
  0.9998336662314, 0.99951352555144, 0.99917807904392, 0.99883645854011, 
    0.99848214894076, 0.99813036362413, 0.99774373617231, 0.99737370241596, 
    0.99696319629837, 0.99655681116692, 0.99611422525556, 0.99569704221991, 
    0.99522455285456, 0.99475000198315, 0.99429063953939, 0.99377568483378, 
    0.99323859462858, 0.9927041137451, 0.99214820598786, 0.99153662725175, 
    0.99091979117422, 0.99036124747381, 0.98972003122979, 0.98892018113621, 
    0.98823429999664, 0.98758839833033, 0.98677049462005, 0.98594761130906, 
    0.98519968528777, 0.98426555707547, 0.98340626403261, 0.98244457988706, 
    0.98146896190681, 0.98038867752832, 0.97942979809755, 0.97828334569119, 
    0.97710683624787, 0.97598421438535, 0.97470731931088, 0.97330936086428, 
    0.97175141452789, 0.97055671444872, 0.96883834678229, 0.96730355409185, 
    0.9656077126903, 0.96386776140564, 0.96197703834648, 0.95986771546181, 
    0.95802505323479, 0.95540774692313, 0.95337987384947, 0.95131316038108, 
    0.94839299174944, 0.94571246255752, 0.94262946489083, 0.93941647920472, 
    0.93652836378093, 0.93293302899503, 0.92910717576869, 0.92529625357158, 
    0.92076362876978, 0.91649929997177, 0.91173148966938, 0.90627079555981, 
    0.90107496290984, 0.89492212880079, 0.88871842047267, 0.88143698057456, 
    0.87487655052524, 0.86599140616773, 0.85765825501356, 0.84854180451466, 
    0.83762256320425, 0.82769858335729, 0.81500316969498, 0.80143102288867, 
    0.78762485218114, 0.7713651312425, 0.75450166013662, 0.73548946832824, 
    0.71585167363623, 0.69181514334144, 0.66601142067417, 0.64048850972306, 
    0.61059149737763, 0.57722658543421, 0.54162929255531, 0.50413735654395, 
    0.45925388696411, 0.41281201145991, 0.36832188727248, 0.31393955630377, 
    0.26453127073998, 0.21472731419663, 0.16381895288933, 0.11455252471166, 
    0.07245032951265, 0.038190333208101, 0.014635981082564, 
    0.0017818017693699, 0.0015831280184339, 0.014192073266231, 
    0.036842512693429, 0.071081675433533, 0.11424007205278, 0.16196194031896, 
    0.21412505839004, 0.26536182114265, 0.31543863801453, 0.36890160741901, 
    0.41211219827243, 0.46132267924411, 0.50242230255062, 0.54302145971699, 
    0.57828058541788, 0.60969418008456, 0.64213859604584, 0.66839642289854, 
    0.69329889624008, 0.71864237394291, 0.73766891067091, 0.75557161467596, 
    0.77337378889107, 0.78962944118793, 0.80422672991688, 0.81747323532895, 
    0.82929388709776, 0.83914576139915, 0.84923900702506, 0.85871672965357, 
    0.86766791928613, 0.87598437458946, 0.88392111417046, 0.89021773283729, 
    0.89595228974203, 0.90188520020258, 0.90736739793092, 0.91258100650251, 
    0.91776217868306, 0.92212765410499, 0.92653974252984, 0.92982000583484, 
    0.93399981158673, 0.93714563734115, 0.94017475116358, 0.94344011494901, 
    0.94639011292938, 0.9489930943677, 0.95155388185779, 0.95391678141917, 
    0.95599573673751, 0.95846505338534, 0.96045233969326, 0.9621064224274, 
    0.96416859542282, 0.96586457817601, 0.9674546238502, 0.96888028288198, 
    0.97067660638411, 0.97190652790924, 0.97344860927497, 0.97476840834432, 
    0.97596950089724, 0.97724108205202, 0.97835146155857, 0.97941209755324, 
    0.98046023977167, 0.98147389464064, 0.98245233195025, 0.98330414591099, 
    0.98423039340088, 0.98505408079061, 0.98591411636717, 0.98665902503132, 
    0.98747456792506, 0.98819201952596, 0.9888826780437, 0.98963471168402, 
    0.9901970313462, 0.99082967598552, 0.99147959300482, 0.99201227527863, 
    0.99263036798681, 0.99318736058979, 0.99370576748374, 0.99417776611401, 
    0.99468504096113, 0.99517513381339, 0.99565960824365, 0.99608682555463, 
    0.99651357015429, 0.99692741597049, 0.99734944466426, 0.99774192082485, 
    0.99810055802253, 0.99847838072461, 0.99883865168835, 0.9991784855018, 
    0.99951043769455, 0.99983318134124,
  0.99985044707244, 0.99956420916375, 0.99926796950124, 0.99896468281629, 
    0.9986505260337, 0.99832399409362, 0.99799878000731, 0.99764618688545, 
    0.99729223786498, 0.99692933217368, 0.99654785254923, 0.99614623314488, 
    0.9957459393022, 0.99534988658562, 0.99487590350298, 0.99443097748085, 
    0.99396702938781, 0.99348213154559, 0.99298766286397, 0.99249895983378, 
    0.99190429538255, 0.99135267537838, 0.99076784814212, 0.99016655388994, 
    0.98952150825151, 0.98889957817132, 0.98817927290516, 0.98750170725973, 
    0.98675305267748, 0.98592764578811, 0.98516719980771, 0.98428986295979, 
    0.98340842677485, 0.98256373866836, 0.98164402329019, 0.98051634372928, 
    0.97960435300266, 0.97845660018588, 0.97731988018182, 0.97605234046119, 
    0.97490785895049, 0.97351688613978, 0.97217461019705, 0.97078278443575, 
    0.96917026278773, 0.96758200383094, 0.96593028345276, 0.9641408100758, 
    0.96227599209903, 0.96021542336152, 0.95837720999809, 0.95589969254913, 
    0.95370097145578, 0.95120589861361, 0.94858937050653, 0.94587140918364, 
    0.94287867065591, 0.93976909828128, 0.93615905409052, 0.93303165586484, 
    0.92868925671459, 0.92502523445757, 0.92030278423059, 0.91563214135428, 
    0.91104173301607, 0.90519130798636, 0.8993596388595, 0.89324880660009, 
    0.88644153765961, 0.87918324919182, 0.87054400686093, 0.86265273708847, 
    0.85291780441961, 0.84286364569999, 0.83085442201208, 0.81974203604681, 
    0.80549983696667, 0.7914151317485, 0.7747015282628, 0.75679436522103, 
    0.73794226834933, 0.7161580724235, 0.69309176428182, 0.66580960318255, 
    0.63660639991036, 0.60492635754538, 0.56983732638079, 0.53102038155215, 
    0.48829077389476, 0.44334788748153, 0.39177798624527, 0.34316198114462, 
    0.28838373889333, 0.2330960928286, 0.1784033274016, 0.12655049133944, 
    0.080719353029007, 0.04274410788691, 0.01637678639787, 
    0.0020451390120542, 0.0016774388290988, 0.015553767322186, 
    0.042758605220392, 0.079671847514674, 0.12766210114558, 0.17864555338985, 
    0.2304243883969, 0.28783291496924, 0.3430930134508, 0.39503059893927, 
    0.4437136293449, 0.48868102342138, 0.53063825334346, 0.57113565718408, 
    0.60559595845034, 0.63812807163601, 0.66744928703969, 0.6941089509133, 
    0.71775743548762, 0.73910997759046, 0.75907247335487, 0.7764212970774, 
    0.79315084106034, 0.80759692536393, 0.82077823236551, 0.83243443421365, 
    0.84362876261975, 0.85483894951956, 0.86428094624009, 0.87214070413141, 
    0.88050385829715, 0.8874350243665, 0.89459679314737, 0.90074267088548, 
    0.90619451857392, 0.91143729968975, 0.916808206148, 0.92153885892645, 
    0.92568506125934, 0.92998987047892, 0.93333531850065, 0.9371454583601, 
    0.94053820862151, 0.9436111265075, 0.94628311627934, 0.94909755318472, 
    0.95172660518046, 0.95423230889642, 0.95657049321398, 0.95869548516509, 
    0.96060085802181, 0.96267962814816, 0.96447260827333, 0.96619438124319, 
    0.96775711253406, 0.96933276867816, 0.97087079572621, 0.97233630408843, 
    0.97379186555144, 0.97501906406161, 0.97626276157115, 0.9773997030362, 
    0.97849740146346, 0.97955288804782, 0.98057187206966, 0.98160230396364, 
    0.98249505403163, 0.98343601286521, 0.98429034446571, 0.98513703549742, 
    0.98592295413752, 0.98671268975622, 0.9874307495718, 0.98814163116323, 
    0.98879960884234, 0.98942369445571, 0.99009326058831, 0.99070492341129, 
    0.99126232051148, 0.99187613591607, 0.9924041209599, 0.99290792160883, 
    0.99340716888545, 0.99389535324786, 0.99440617566868, 0.9948330978942, 
    0.99527540484861, 0.99571120413962, 0.99611825498165, 0.9965147852922, 
    0.99690063619465, 0.9972743161271, 0.99763413983155, 0.99797275692766, 
    0.99832686278952, 0.99864261342473, 0.99896278909131, 0.99926667786079, 
    0.99956322216403, 0.99984994754695,
  0.99985730728261, 0.99958541068613, 0.99930508533053, 0.99901638893196, 
    0.99871738521081, 0.99841416058026, 0.99809575004422, 0.99776630959498, 
    0.99743422611417, 0.99708009609329, 0.99672144124135, 0.99635404775724, 
    0.99596273360687, 0.99556884661047, 0.99514598158365, 0.99471434250421, 
    0.99427297819918, 0.99383025267943, 0.9933374287136, 0.99282648515063, 
    0.99232533873687, 0.99180926822281, 0.99123595317037, 0.99064917349509, 
    0.99004974093099, 0.98943838118279, 0.98879034872066, 0.98810656172099, 
    0.98737539936788, 0.98665088945134, 0.98591807827426, 0.98513051268936, 
    0.98426578145881, 0.98337118405858, 0.98249629610887, 0.98157897844506, 
    0.98054867010112, 0.97953445694583, 0.9784687286095, 0.97727549571002, 
    0.97610744690431, 0.97484490652794, 0.97355683876454, 0.97206865776053, 
    0.97081207733607, 0.96918248302424, 0.96759116166988, 0.96590289886886, 
    0.96420335508067, 0.96217765410402, 0.96026613860673, 0.95826874535168, 
    0.95593772164621, 0.95349567142011, 0.95114520799143, 0.94856151090324, 
    0.94553303126487, 0.94261328847799, 0.93936060155289, 0.93584509358813, 
    0.93228892592635, 0.92861809638171, 0.92428403762339, 0.91950147079486, 
    0.91499454222615, 0.90978557588478, 0.90416691250778, 0.89807805383675, 
    0.89162618775817, 0.88472237317498, 0.87680782415363, 0.86854832757066, 
    0.85932225759845, 0.84924364695254, 0.83885087037711, 0.82699292472805, 
    0.81401281378647, 0.80015324106343, 0.78389544292823, 0.76682712659646, 
    0.74786954775588, 0.72636041488942, 0.70322122512053, 0.6780024810244, 
    0.64782803775108, 0.61812149218155, 0.58105136936378, 0.54530793691842, 
    0.50259070966742, 0.45607143795333, 0.40784710901645, 0.35379209544766, 
    0.2986762802123, 0.24150661023888, 0.18549752831401, 0.13392439816902, 
    0.084989925797726, 0.045003937984756, 0.016660175063776, 
    0.0020115790593614, 0.0017212881539766, 0.016567622445174, 
    0.045108333363228, 0.083771024405837, 0.13259736702836, 0.18508717998529, 
    0.24303473546172, 0.29883556892489, 0.3538222186663, 0.40598956340117, 
    0.45703230686783, 0.50277814577425, 0.54591968590632, 0.58243574294555, 
    0.61916046662368, 0.65109537850726, 0.67795714002913, 0.70457052494999, 
    0.72745732779335, 0.74973264915323, 0.76804607923319, 0.78559596040593, 
    0.80122934891955, 0.8155246019496, 0.82784285661606, 0.83998958413682, 
    0.85094219212241, 0.86100846557461, 0.86947040334682, 0.87816994836631, 
    0.88575987308714, 0.8925425545005, 0.89928382983327, 0.90506930124901, 
    0.9106767806867, 0.91584548770638, 0.92074083135618, 0.92509767775086, 
    0.92941465578758, 0.93289085300114, 0.93693311402938, 0.93989893215814, 
    0.94326347475105, 0.94632932042765, 0.94881543798257, 0.9515600088659, 
    0.95394940015847, 0.95644394880065, 0.95848624084817, 0.96068926911839, 
    0.96264576805788, 0.96437495596506, 0.96615629091646, 0.96792592309233, 
    0.96942399717131, 0.97099657847357, 0.97228897029767, 0.97373656637306, 
    0.97494718591317, 0.97624303012351, 0.97742136016781, 0.97849035134724, 
    0.97956840402615, 0.98059294476499, 0.98157751689882, 0.98251472364556, 
    0.98341527494367, 0.98429177626035, 0.9850777998007, 0.98587061728183, 
    0.9865924135056, 0.98738351358592, 0.98806713907603, 0.98873657095187, 
    0.98938304302894, 0.99000116451087, 0.99059463253303, 0.99119375060978, 
    0.99172960712541, 0.9922487814147, 0.99279454126815, 0.99329091797765, 
    0.99377163598978, 0.99422325588198, 0.99467093816616, 0.99510586261267, 
    0.99551978725839, 0.99592451059344, 0.99632349476083, 0.99670224848771, 
    0.99705533470115, 0.99741226399329, 0.99775990866554, 0.99808313328012, 
    0.99840491376207, 0.99871411845297, 0.99901351984316, 0.99930394065931, 
    0.9995850597017, 0.99985751116018,
  0.99986389336822, 0.99960506027409, 0.99933827803332, 0.99906393729815, 
    0.99877806157765, 0.99848737686751, 0.99818686935799, 0.99787714325282, 
    0.99755476738337, 0.99721958698395, 0.99687966570117, 0.99652419459206, 
    0.99615251030205, 0.99578074517674, 0.99538178555429, 0.99497825574351, 
    0.99456507465978, 0.99409887407786, 0.99363650787928, 0.99318659647234, 
    0.99268393479839, 0.99217237884121, 0.99166508828703, 0.99111776213718, 
    0.99051782856628, 0.98992464610519, 0.98933779270217, 0.98865668695209, 
    0.9879751860943, 0.98729480779257, 0.98656682782284, 0.98581486990774, 
    0.98501917845474, 0.98418052349998, 0.98338848381663, 0.98236343546856, 
    0.98149847244197, 0.98049902139236, 0.97948538236587, 0.97834658043053, 
    0.97725283310542, 0.97601076678793, 0.97487470446292, 0.97350613346281, 
    0.97203515993887, 0.97058138492031, 0.96911743480489, 0.9674802489436, 
    0.96596648026848, 0.96402165138461, 0.96212126654139, 0.96014523893636, 
    0.95790401232902, 0.95583748040127, 0.95332336152106, 0.95091362249888, 
    0.94801312219576, 0.94536412263632, 0.94214955726045, 0.93880516733325, 
    0.93540361406049, 0.93163326378552, 0.92765865499012, 0.92350238735297, 
    0.91899838115553, 0.91350807926405, 0.90832740784701, 0.90275239993745, 
    0.89631668052242, 0.88977677413063, 0.88205439762777, 0.87447360407313, 
    0.86538557034922, 0.85604574305949, 0.84516652352298, 0.83406949315883, 
    0.82156358783362, 0.80725847287955, 0.79190831550824, 0.77587925340766, 
    0.75726121313246, 0.73677335769645, 0.71337093377918, 0.68792611558896, 
    0.66053635552578, 0.62989291341383, 0.59526791707981, 0.55615505604866, 
    0.51300375516962, 0.46750373425003, 0.41901496383918, 0.36550647760291, 
    0.30932724697479, 0.25338521567769, 0.19332150456147, 0.13969234845701, 
    0.089126623343549, 0.046625467014727, 0.017341971071812, 
    0.0019795355619478, 0.0018436524348644, 0.017379884735009, 
    0.048148475618749, 0.08674766354063, 0.13822736405751, 0.19394360866289, 
    0.25089219063895, 0.30865839759069, 0.36496074372779, 0.42128518668856, 
    0.46875893445776, 0.51475274237258, 0.55761630880158, 0.59583796429484, 
    0.6292631232383, 0.66153311570512, 0.69055644205351, 0.71431599597819, 
    0.73861565952132, 0.75780446375421, 0.77634636136614, 0.79354326509776, 
    0.80877480574758, 0.82321385725779, 0.83476883534377, 0.8462021868464, 
    0.8567189397407, 0.86652032433974, 0.87514892246787, 0.88315722633053, 
    0.89052746939551, 0.89745512997388, 0.90313651424799, 0.90934948613474, 
    0.9148236695334, 0.91929916126215, 0.92421164707857, 0.92818656144267, 
    0.93239038357459, 0.93595186270458, 0.93954373711053, 0.94261975752295, 
    0.94583379464639, 0.94853835458267, 0.95133644721652, 0.95372267266905, 
    0.95621342420523, 0.95836238165065, 0.96047837454903, 0.96246102329957, 
    0.96428841558518, 0.9661144126809, 0.96782309902879, 0.96931774499853, 
    0.97092568579555, 0.97228399277585, 0.97359760175216, 0.97487560696452, 
    0.9761975572376, 0.97733455030679, 0.97845136063681, 0.97952846548659, 
    0.98055879159729, 0.98148414819286, 0.98251876698789, 0.9833913739669, 
    0.98415653845975, 0.98505962212187, 0.98582908674755, 0.98656936577849, 
    0.98727730983976, 0.9879716357362, 0.98861067931803, 0.98928480454533, 
    0.98990327366702, 0.99047781696278, 0.99107029983444, 0.99162540549415, 
    0.99213611772807, 0.99263656518967, 0.99313811482738, 0.99359751792786, 
    0.99406797130205, 0.99451187887254, 0.99493323179655, 0.99535426298413, 
    0.99573012309845, 0.99613539104422, 0.99649475312709, 0.9968677451825, 
    0.99720634343784, 0.99754256160936, 0.99786625345261, 0.99817755604935, 
    0.99848303429419, 0.99877410114046, 0.99906087414593, 0.99933732879679, 
    0.99960434084177, 0.99986351059882,
  0.99986664857751, 0.99961359234683, 0.99934870419362, 0.99908859221607, 
    0.99881834614205, 0.99851642019812, 0.99823887533218, 0.99791523123194, 
    0.99760763249265, 0.99731858435377, 0.99689196474451, 0.99663316838283, 
    0.99625889855342, 0.99589361380773, 0.99548165054844, 0.99508167004283, 
    0.99469694763677, 0.994244663208, 0.99380995335097, 0.99329107345698, 
    0.99292353428185, 0.99232201490496, 0.99194535612795, 0.99130534418226, 
    0.99063473839328, 0.99011234584377, 0.98961639500751, 0.98890095871812, 
    0.98834097879011, 0.98761142040688, 0.98682731877236, 0.98617340932427, 
    0.9853723224756, 0.98448251724981, 0.98372372864267, 0.98295565241654, 
    0.98193336419454, 0.98084558528604, 0.97988451913038, 0.97904188681207, 
    0.97772797989478, 0.97652185311712, 0.97541035692342, 0.97398535599317, 
    0.97269702061074, 0.97145444623832, 0.97011926792029, 0.96842273114351, 
    0.96671637221056, 0.96480269070799, 0.96269684009627, 0.96077118147837, 
    0.95887788383713, 0.95701193438552, 0.9548525855349, 0.95223066795875, 
    0.94913090945898, 0.94603009242633, 0.94310937295484, 0.94026636034559, 
    0.93685067734335, 0.93354533387129, 0.92962147992884, 0.92474788253431, 
    0.9201310269915, 0.91513291175856, 0.91003706011728, 0.90498026301766, 
    0.89927405106187, 0.89275759022287, 0.88558762141328, 0.87642175761091, 
    0.86722923826849, 0.85787061789724, 0.84754040782059, 0.8390655132324, 
    0.82640670918067, 0.8112726009048, 0.79655626832482, 0.77981202611086, 
    0.75993817637913, 0.7393630548729, 0.71963782831942, 0.69548920804513, 
    0.66624355918228, 0.63166353623369, 0.59970849013307, 0.56195602619801, 
    0.52134847990365, 0.47571981439, 0.42547985455987, 0.37184378376166, 
    0.31235433829521, 0.25549211515992, 0.1962205349047, 0.14373120436868, 
    0.092103573848417, 0.049932570163638, 0.016545472461787, 
    0.0023613875258121, 0.0022685154888188, 0.01745672510524, 
    0.046094844797691, 0.087968292942644, 0.14451564300782, 0.19674277037537, 
    0.25999954620124, 0.31884956710539, 0.37283094739499, 0.42305574879004, 
    0.4743562122055, 0.51689623443394, 0.56208142478857, 0.60015057901303, 
    0.63459034722802, 0.66763582130521, 0.6951769386282, 0.71885103023365, 
    0.74214292437687, 0.76166941692611, 0.78080423916151, 0.79750895932142, 
    0.81258597737652, 0.82563906931209, 0.83892673694328, 0.84990343303515, 
    0.86043993942273, 0.87004941448275, 0.87719436322631, 0.88490664471983, 
    0.8919311387184, 0.89950460761754, 0.90573699273546, 0.91233577079612, 
    0.91662485895273, 0.92093225881546, 0.92552735202931, 0.9302730957517, 
    0.93377295404506, 0.93747176123252, 0.94075258763136, 0.94374372070173, 
    0.9472531292172, 0.94974182464737, 0.95238327481726, 0.95489706664713, 
    0.95695527627584, 0.95959120212282, 0.96145297900115, 0.96297218110798, 
    0.96486781289515, 0.96670957333298, 0.96848438826327, 0.97020465578539, 
    0.97150591886002, 0.9730523865242, 0.97419995230693, 0.97562357172336, 
    0.97674561930268, 0.97783512439523, 0.97891448518582, 0.98002446060204, 
    0.98091359721388, 0.98188352673277, 0.98280479863589, 0.98367495741571, 
    0.9846263122936, 0.98537733487104, 0.98609758978988, 0.98680013975759, 
    0.98763618897219, 0.98830805924939, 0.98898378629489, 0.98949870592741, 
    0.99014239600125, 0.99065947717028, 0.99126104693442, 0.99184836100064, 
    0.99237932685105, 0.99288302126254, 0.99330199646558, 0.99373737576406, 
    0.99418179389229, 0.99462468221237, 0.99502683300104, 0.99545917350964, 
    0.99589597511686, 0.9962323710898, 0.99658523477056, 0.99691129580305, 
    0.99726619485002, 0.99759335546306, 0.99790805985129, 0.99824132106471, 
    0.99851574278731, 0.99880252109384, 0.99908524209808, 0.99935459037328, 
    0.99961605992702, 0.99986691653237,
  0.99987499334911, 0.99963846846195, 0.99939571280596, 0.99914486790764, 
    0.99888673830732, 0.9986195950523, 0.99834618743621, 0.99806171055933, 
    0.99776593131061, 0.99746578879909, 0.99715280228825, 0.9968246042042, 
    0.99649386180219, 0.99614436661921, 0.99577333743255, 0.99541637753459, 
    0.99501559764138, 0.99461399833667, 0.99419865114985, 0.99378346731375, 
    0.99331446005656, 0.9928403023589, 0.99238027892206, 0.99186322452916, 
    0.99133861229949, 0.99077170595156, 0.99026793749433, 0.98965218783775, 
    0.9890164867857, 0.98836266277255, 0.98772540169023, 0.98701459231202, 
    0.98627898410871, 0.9855816646287, 0.98469581484102, 0.98399128514305, 
    0.98308298065487, 0.98214796905381, 0.98123301708931, 0.98025353877508, 
    0.97920796338368, 0.97807646587114, 0.97698917468711, 0.97578849699097, 
    0.9744539757583, 0.97308603443102, 0.97179684452847, 0.97031578488767, 
    0.96868883569607, 0.96715750444202, 0.96534627569528, 0.96341718497845, 
    0.96166061984939, 0.95954116731974, 0.95726949666883, 0.95490660560852, 
    0.95256685518981, 0.95009849015828, 0.94688730119351, 0.94393098548632, 
    0.94089856954081, 0.93742643616056, 0.93386495286472, 0.92970930729263, 
    0.92561700337066, 0.9208038897449, 0.91589223768424, 0.91040893615589, 
    0.90487429039761, 0.89857015904963, 0.89158793613134, 0.88407806274011, 
    0.87595863593826, 0.86710072940741, 0.85753620202758, 0.84612902544173, 
    0.83484828362705, 0.82195416290687, 0.80754475323566, 0.79139545945778, 
    0.77344913827327, 0.75484803466651, 0.73207588391683, 0.70804210903897, 
    0.68033341866889, 0.65034353371277, 0.61678758720854, 0.57987443413702, 
    0.53757438064709, 0.49131590204023, 0.44188494508929, 0.38720945214926, 
    0.32977855716505, 0.26836410896391, 0.20877362384503, 0.15050706040989, 
    0.096602739009155, 0.05068307618488, 0.019234794924854, 
    0.0020336819415284, 0.0020924184706647, 0.019015298476881, 
    0.051963258850431, 0.095884468281232, 0.15004727827511, 0.20861514664429, 
    0.26875824992564, 0.32785211425073, 0.38878601518619, 0.44099538460018, 
    0.49225818932939, 0.53729108721812, 0.58098492913974, 0.61615488631955, 
    0.65190757949814, 0.68178252625197, 0.70836687560365, 0.73264438969539, 
    0.75584692037153, 0.77418609245725, 0.79252789311507, 0.80770876372875, 
    0.82226999102498, 0.83525171999886, 0.84711913620985, 0.85842638310697, 
    0.86714011027253, 0.87694343563436, 0.88491125690171, 0.89199996947992, 
    0.89898182000344, 0.9053367198331, 0.91098672388276, 0.91668063132529, 
    0.9212858064963, 0.92581560184939, 0.9301821979552, 0.93411858166334, 
    0.93774798721556, 0.94126624589857, 0.94444185885153, 0.94741395060049, 
    0.95014180416175, 0.95291450508091, 0.95526845963648, 0.95753383987422, 
    0.95966519999555, 0.96185876097069, 0.96367728301439, 0.96564538659229, 
    0.96722576952951, 0.96898178966576, 0.97049410017715, 0.97187710204553, 
    0.97328349975387, 0.97464572297584, 0.97587912863859, 0.97709584247056, 
    0.97820276345944, 0.97927897447577, 0.98026698423695, 0.98128478342401, 
    0.98220507066008, 0.98310006513144, 0.98400980940607, 0.98481790007826, 
    0.98554762024223, 0.98633841742762, 0.98701759261327, 0.98773453834832, 
    0.98839016164479, 0.98903614761938, 0.98963420002085, 0.99024120503372, 
    0.99076449072342, 0.99134731222853, 0.99184751524196, 0.99232739243625, 
    0.9928437285468, 0.99329258145061, 0.99376741619071, 0.99418012513891, 
    0.99459549624995, 0.9949974273777, 0.99538677389759, 0.99576246200294, 
    0.99613204098222, 0.9964644244853, 0.99680863220818, 0.99714250668946, 
    0.99745001884625, 0.99776042483299, 0.99805347954968, 0.99833994721075, 
    0.99861563562756, 0.99888225002277, 0.99914350809059, 0.99939402833514, 
    0.99963845083683, 0.99987493579829,
  0.99988000900631, 0.99965326424171, 0.99942142638871, 0.99917914542265, 
    0.99893450942111, 0.99867585023725, 0.99841396435804, 0.99814566262429, 
    0.99786100327707, 0.9975687845791, 0.99726972251602, 0.99696551743216, 
    0.99662544892814, 0.99631409440886, 0.99594578740596, 0.99559114751719, 
    0.99523932943805, 0.99485277797986, 0.99443387289029, 0.99401654144369, 
    0.99360430925972, 0.99315932922686, 0.9926950069871, 0.99218178551532, 
    0.9916951639215, 0.99118089285473, 0.99063893066627, 0.99006116287982, 
    0.98947680136591, 0.98888051975711, 0.98825245241509, 0.98755290924627, 
    0.98689764952689, 0.98612516721056, 0.98542678280856, 0.98457830997937, 
    0.98379306125312, 0.98288577283976, 0.98201476789183, 0.98105560772273, 
    0.98003676413756, 0.97904251145327, 0.97794281892431, 0.97674902636019, 
    0.97559562136896, 0.97420439350593, 0.97296348379814, 0.97154415718509, 
    0.97001376290215, 0.96832494667018, 0.96677587468842, 0.96511728879394, 
    0.96308702361021, 0.96120975728712, 0.95898973850765, 0.95691206425843, 
    0.95439295894024, 0.95196775626528, 0.94916335878207, 0.94616717669483, 
    0.94322798263007, 0.93976016341429, 0.93653275374858, 0.93275835795382, 
    0.9285580020795, 0.92397857845728, 0.91915523873462, 0.91380086163262, 
    0.90872094646678, 0.90219504449144, 0.89536556160145, 0.88871228508349, 
    0.88089953956116, 0.87218172403672, 0.86245475105954, 0.85206656347968, 
    0.84116033485338, 0.82809368866607, 0.81405872698217, 0.79845739887118, 
    0.78155460771148, 0.76193960183334, 0.74081902215425, 0.71745833607239, 
    0.6898112083102, 0.66030265689144, 0.62789255902721, 0.58911006459102, 
    0.54834617482061, 0.50204975584599, 0.45218476032695, 0.39797212797904, 
    0.33771014706612, 0.27712178607534, 0.21630406934315, 0.15585446792976, 
    0.10027198266505, 0.054257787702978, 0.020027106085268, 
    0.0022706619055483, 0.0023055525598021, 0.02047135554633, 
    0.054010641010668, 0.10030667626276, 0.15472798854949, 0.21467776450528, 
    0.27880580790871, 0.33871780990308, 0.39801232739722, 0.45065789386079, 
    0.50336140560139, 0.55056142750953, 0.58992251305353, 0.62689427167276, 
    0.65991686051084, 0.69071847729326, 0.71750750264014, 0.74196964068199, 
    0.76288403740518, 0.78210561696614, 0.79916045487872, 0.81476382364372, 
    0.82787238405201, 0.84102194071509, 0.85237268092288, 0.86321609329315, 
    0.87245713667724, 0.88118876621279, 0.88943492096037, 0.89620547507037, 
    0.90258255277613, 0.90837220286948, 0.91477483997188, 0.91949009345463, 
    0.92432998820464, 0.9288453604182, 0.93284480250049, 0.93671134528901, 
    0.94021387643471, 0.94351525288003, 0.94646625502588, 0.94951423098321, 
    0.95208905783338, 0.9546745015541, 0.95699254008659, 0.95937142545057, 
    0.96136794997929, 0.96338565456985, 0.9650708720035, 0.96694785766313, 
    0.96872091802128, 0.97013106751092, 0.97166604400259, 0.97304516824287, 
    0.97443785548165, 0.97560504582047, 0.97682785856801, 0.97801904464836, 
    0.97907472717686, 0.98011220144072, 0.98117685664665, 0.98204176630072, 
    0.98296696663961, 0.98378345215423, 0.98460166368206, 0.98541243963373, 
    0.98613488494945, 0.98692473886195, 0.9875672053756, 0.98827365980037, 
    0.98884169949106, 0.98950769690941, 0.99007369112059, 0.9906424367244, 
    0.99116301741772, 0.99171427522786, 0.99217175588709, 0.99267395859379, 
    0.99312938728787, 0.99358428450447, 0.9940255457688, 0.99442898937063, 
    0.9948156636477, 0.99521844582679, 0.99558499505734, 0.99593672376534, 
    0.99629602518289, 0.99662863735819, 0.99693887637352, 0.99725984590324, 
    0.99756474132028, 0.99785351596866, 0.99813240944749, 0.99840880562721, 
    0.9986743834879, 0.99892989469575, 0.99917845946532, 0.99941951956258, 
    0.99965297361008, 0.99987967564379,
  0.99989925045671, 0.99971212223545, 0.999520786658, 0.99932374489996, 
    0.99910817615074, 0.99891305922831, 0.9986711153494, 0.99846264588019, 
    0.99823668711651, 0.99797786736838, 0.9977282290304, 0.99749548755546, 
    0.99720909176679, 0.9969259723028, 0.99665766804554, 0.99633175528316, 
    0.99603307167498, 0.99572455113266, 0.99543135076718, 0.99502300660419, 
    0.99469885087306, 0.99431993756831, 0.99391434913973, 0.99352268805482, 
    0.99312011844412, 0.99270925705158, 0.99219025421681, 0.99175734136673, 
    0.9913000594904, 0.99080249942361, 0.99024269225613, 0.9896752974071, 
    0.98913965941931, 0.98850843147316, 0.98788358249913, 0.98723294589804, 
    0.98650866867849, 0.98584766196806, 0.98507012662708, 0.98434183376818, 
    0.98346229956477, 0.98256697717439, 0.98165827880701, 0.9808294245431, 
    0.97972166401726, 0.97868285033033, 0.97762342437134, 0.97638652920326, 
    0.97517214208202, 0.97383000016142, 0.97230253833705, 0.9708662084477, 
    0.96948062556655, 0.96776398547943, 0.9660824908281, 0.96415490478087, 
    0.96211457124883, 0.96011741529994, 0.95783273596878, 0.95537648339601, 
    0.95261254461523, 0.95018789695275, 0.94712876539827, 0.94387872175754, 
    0.94073306209386, 0.93654096635678, 0.9325198933068, 0.92793534135221, 
    0.92363932927313, 0.91842864578064, 0.9125128671265, 0.90629658990813, 
    0.89962837943315, 0.89225612225555, 0.88421625958423, 0.87459114464715, 
    0.86547127017165, 0.85384596295382, 0.84176239880573, 0.82779393603665, 
    0.81334264995182, 0.79550912270215, 0.77568533493156, 0.75557869766522, 
    0.73043737859907, 0.70224403032706, 0.6719010839506, 0.63641960055466, 
    0.59587399071679, 0.55010970545594, 0.49728467451084, 0.44432486421401, 
    0.3857013719635, 0.31491138575921, 0.25014352607412, 0.18252351116675, 
    0.11903178985595, 0.063065995787243, 0.02439052675473, 
    0.0031244165734346, 0.0029310419367534, 0.024186576013702, 
    0.064634844757667, 0.11936778642812, 0.18097723599439, 0.25360086015955, 
    0.31679073337285, 0.38216774786211, 0.44487554836644, 0.49937820587103, 
    0.54755099276099, 0.59661863634283, 0.63593389938954, 0.67101006413796, 
    0.70311013144611, 0.73076358506379, 0.75404462225768, 0.77697196967185, 
    0.79416401345629, 0.8127362568144, 0.82771035742817, 0.84094443811625, 
    0.85372913072859, 0.86472478256742, 0.87441032709771, 0.88378938385182, 
    0.89183328487283, 0.89915157371731, 0.9061956795051, 0.91218566344744, 
    0.91811416316047, 0.9232124103083, 0.92778128919587, 0.9324063660442, 
    0.93628143370615, 0.9399871671717, 0.9435546368874, 0.94672542232802, 
    0.94967945244639, 0.95288793985615, 0.95514872453544, 0.95742308127821, 
    0.95996038660863, 0.96206377440867, 0.96395824596599, 0.96589825541143, 
    0.96775429545796, 0.96936304541756, 0.97088243561958, 0.97243079537382, 
    0.97375667443966, 0.97506956968144, 0.97639844026275, 0.9775644705249, 
    0.97864151843531, 0.97963128891393, 0.9807418579092, 0.9817231230795, 
    0.98258507003846, 0.98347118759029, 0.98426367331863, 0.98505513753214, 
    0.98593521759348, 0.98654802310947, 0.98715697386579, 0.98789478358033, 
    0.98853950198356, 0.98913691824542, 0.98975176124534, 0.99020360709514, 
    0.99082552658551, 0.99127361435328, 0.99179582813037, 0.99230166046144, 
    0.99266821846239, 0.99316608939968, 0.99352797386633, 0.99395877360199, 
    0.99432491257909, 0.99465911299244, 0.99507581069741, 0.99543480274311, 
    0.99573621740198, 0.99602871709459, 0.99636112210444, 0.99666686398505, 
    0.99693978190227, 0.99720887263586, 0.99748709255059, 0.99773161047265, 
    0.99799858576831, 0.99822804085349, 0.99846046505649, 0.99868840978245, 
    0.99890439470827, 0.99911590383157, 0.99931843555225, 0.99952021594488, 
    0.99971223480063, 0.99989892196589,
  0.99991267991037, 0.99975261295193, 0.99958790351018, 0.99941853560338, 
    0.99924368732002, 0.9990610709144, 0.99887761839427, 0.99868200398862, 
    0.99848100334945, 0.99827898443045, 0.99806030652476, 0.99784314788754, 
    0.9976086571684, 0.9973763692976, 0.99712540429765, 0.99687559218445, 
    0.99660518384592, 0.99633658881402, 0.99604283436775, 0.99575769011206, 
    0.99544888058012, 0.99513167354405, 0.99479823655229, 0.99444853577194, 
    0.99409585908619, 0.99372762460336, 0.99333827401467, 0.99292225719798, 
    0.99252184437892, 0.99209349540627, 0.99162025448134, 0.99117626253191, 
    0.99065907383749, 0.99013260429569, 0.98964536043689, 0.98904526533284, 
    0.98844385686785, 0.98786904865814, 0.98721558431088, 0.98655776543719, 
    0.98581253487553, 0.98506570168008, 0.98429374646376, 0.98352797661488, 
    0.98264518025991, 0.98171388574688, 0.98073720082714, 0.97983992476691, 
    0.9787209054664, 0.97755929588366, 0.97640157102858, 0.97521611612731, 
    0.97373749778622, 0.97241007281812, 0.97089683418008, 0.96925557906503, 
    0.96764138024513, 0.96571512131216, 0.96378962514376, 0.96168513613646, 
    0.95954743353979, 0.95707405871529, 0.95460624508312, 0.95156225247545, 
    0.94878135127802, 0.94541885940592, 0.94203774114521, 0.93813977858822, 
    0.93397432696356, 0.9294982060525, 0.92466869509411, 0.91924333239553, 
    0.91338027105724, 0.90660016901789, 0.89964173240048, 0.89150589382675, 
    0.88277926456656, 0.8730000263667, 0.8617575063838, 0.84953675646483, 
    0.83583815094469, 0.82004977141407, 0.8030049789008, 0.78248346936509, 
    0.76036744462785, 0.73453089521226, 0.7047212672029, 0.67198873878012, 
    0.63358572841359, 0.58875284781791, 0.54058914844505, 0.48319533331859, 
    0.42134170280357, 0.35302274392073, 0.27921320279116, 0.20755379641557, 
    0.13631750656983, 0.07368693979733, 0.0281101278944, 0.0034376913960752, 
    0.0033520092943731, 0.028450018419281, 0.075660351862104, 
    0.1368506102785, 0.20785561234118, 0.28135104539545, 0.3529503360466, 
    0.42069457229688, 0.48406352168589, 0.53897650360815, 0.58727134747037, 
    0.6327151568246, 0.67096648930189, 0.70340772463412, 0.73376007468319, 
    0.75907245247494, 0.78179563583474, 0.80140874193435, 0.81952809717199, 
    0.83490246407527, 0.8483429056909, 0.86094360107724, 0.87169473920823, 
    0.88186302533753, 0.89069013264312, 0.89862776666629, 0.90599029503056, 
    0.9124140556173, 0.91829205386095, 0.9237984945075, 0.92889834855849, 
    0.93350549957659, 0.93747944296043, 0.94144773831951, 0.94485361209816, 
    0.94824654068339, 0.95126238323315, 0.9540359510016, 0.95664400182289, 
    0.95914337006329, 0.96135229924838, 0.96348814308798, 0.96549205355926, 
    0.96729941521615, 0.96906329310762, 0.97065819922624, 0.97212333779504, 
    0.97367413799577, 0.97508670046663, 0.97620071474486, 0.97742378958009, 
    0.97862248161204, 0.97970924234228, 0.98071778263022, 0.98172039933793, 
    0.98257219393435, 0.98348934857259, 0.98433433093021, 0.98506539781712, 
    0.98580770847134, 0.98655227016538, 0.98724336007516, 0.98786190514827, 
    0.98850392476079, 0.98908110040622, 0.98964798974541, 0.99019820270456, 
    0.99069196964944, 0.99123106959688, 0.99166972702086, 0.99213988718264, 
    0.99257435970329, 0.99298901781555, 0.99337766270749, 0.99378203420691, 
    0.99413737457759, 0.99450812447603, 0.99483514642719, 0.99516397752681, 
    0.99548340330372, 0.9957847852998, 0.99608473937791, 0.99635919223544, 
    0.99663848804518, 0.99688939316245, 0.99714935894357, 0.99738884877567, 
    0.997628430078, 0.99784903732901, 0.99807048020644, 0.99828310419729, 
    0.99848662370806, 0.99868530730604, 0.99887900458764, 0.99906441876038, 
    0.99924283034489, 0.99941843611974, 0.99958795015897, 0.9997523460111, 
    0.99991261923904,
  0.9999225443078, 0.99978262719187, 0.99963849844115, 0.9994902500636, 
    0.9993371322698, 0.99918028925658, 0.99901740871019, 0.99884766474312, 
    0.99867368171863, 0.99849293862972, 0.99830475674604, 0.99811398969468, 
    0.99791326987599, 0.997704040559, 0.99748789471273, 0.99727058387904, 
    0.9970306172408, 0.99679445710137, 0.99654326667901, 0.99628304422548, 
    0.99601659042652, 0.99574151460599, 0.99545756593952, 0.99513546623531, 
    0.99482138251042, 0.99453510839977, 0.99416082004718, 0.9938432086583, 
    0.99344971666869, 0.99307420568547, 0.99266140834724, 0.99226650786929, 
    0.99184891872648, 0.99139122969646, 0.99090637791691, 0.99039543078662, 
    0.98990803302735, 0.98938269303295, 0.98879487057763, 0.98825701082794, 
    0.98760006924802, 0.98695576397163, 0.98627746429266, 0.98555107953762, 
    0.98480321821106, 0.98401059536733, 0.98319709437323, 0.98232349746638, 
    0.98135664586885, 0.98041483035189, 0.97932612807953, 0.9782713492401, 
    0.97706252953539, 0.97579087036272, 0.97459077700466, 0.97310232488975, 
    0.97162301944234, 0.96996969945532, 0.96829646025686, 0.96647312821269, 
    0.96451998633191, 0.96239113267048, 0.96008301356667, 0.95759649983774, 
    0.95512108942906, 0.95204627835637, 0.94913119618695, 0.94566340152794, 
    0.94184067814452, 0.93796968546857, 0.93353856153875, 0.92892416905119, 
    0.92331507187013, 0.91758000888116, 0.91136742824554, 0.90419020583201, 
    0.89584608618919, 0.88761144499698, 0.87736330485556, 0.86620783300413, 
    0.8532996129688, 0.83941934313036, 0.8238604983601, 0.80529952371122, 
    0.78388019614724, 0.75982388343599, 0.73226112005322, 0.7008594872804, 
    0.66324924380237, 0.62209177115534, 0.57235886467255, 0.51728232817168, 
    0.45495413704991, 0.38392682139657, 0.30691046369111, 0.2292908643174, 
    0.15371658823226, 0.083878083718948, 0.031721486947958, 
    0.0033927413031519, 0.0035065528532715, 0.03207770996875, 
    0.085294906485776, 0.15281588571482, 0.22945781468108, 0.30778630817631, 
    0.38433551304621, 0.45254416802387, 0.51647372247134, 0.57194238195882, 
    0.61973023131853, 0.66274746183858, 0.69905883114656, 0.73121581329802, 
    0.75798297105377, 0.78237803663632, 0.8029255678459, 0.82180011407528, 
    0.83812889862068, 0.85187377898875, 0.86482281009285, 0.87593247596462, 
    0.88630795598839, 0.8944663656164, 0.90270756063191, 0.91001935767958, 
    0.91668955720528, 0.92219261965564, 0.92783108727493, 0.93256079252786, 
    0.93714849084379, 0.94102768627352, 0.94502119630261, 0.94817185526355, 
    0.9513867154928, 0.95444400181268, 0.95704487035899, 0.95961860052699, 
    0.96178005994252, 0.96419435786029, 0.96596182397655, 0.96787458633344, 
    0.96968881578987, 0.97121575259895, 0.97294677533988, 0.97419853431656, 
    0.97560402427366, 0.97687370443774, 0.97808268302408, 0.97924071069902, 
    0.98023371635948, 0.98129373469056, 0.98219733141172, 0.9831147961267, 
    0.9839803775476, 0.98476448396383, 0.98557338818922, 0.98627478558715, 
    0.98696628481526, 0.98762124853955, 0.98827360062902, 0.98883504342955, 
    0.98943319836103, 0.98996383724976, 0.99048121242664, 0.99097297837894, 
    0.99143742728451, 0.99187935970628, 0.99235469596603, 0.99273582855682, 
    0.99316326045585, 0.99350879428969, 0.99389252593715, 0.99423724938922, 
    0.99456279606603, 0.99489586176184, 0.99521177180163, 0.99550052135908, 
    0.99578612273219, 0.99605833005815, 0.99632686226247, 0.99658326358636, 
    0.99682788404253, 0.99705955144086, 0.99728917128175, 0.99750762938492, 
    0.99772029078997, 0.99792328290363, 0.99812575703171, 0.99831106238111, 
    0.99849629789384, 0.99867629098222, 0.99885136221102, 0.99901595113667, 
    0.99917925585345, 0.99933638993412, 0.9994897573556, 0.99963820348799, 
    0.99978228241163, 0.99992226876095,
  0.99993016012667, 0.99980665702355, 0.99967919733932, 0.99954527610918, 
    0.9994059352246, 0.99927136663076, 0.99912936933994, 0.99897539004039, 
    0.9988394116332, 0.99864274717407, 0.99849381564639, 0.99831403208588, 
    0.99816595153257, 0.99795026804737, 0.99779149818669, 0.99756344485035, 
    0.99734694086672, 0.99713441395468, 0.99694753370341, 0.99670822837286, 
    0.99645671959759, 0.99618062586766, 0.99594329018435, 0.9957048504304, 
    0.99550346604071, 0.99512326187234, 0.99484512300335, 0.9944647356606, 
    0.99414581376934, 0.9937834319546, 0.99355812631991, 0.99320207202652, 
    0.99274557631344, 0.99231673601987, 0.991855390459, 0.99148606030959, 
    0.99106088807452, 0.99062003241763, 0.98999923979173, 0.9895950933622, 
    0.98899057395314, 0.98842550060577, 0.98776407833363, 0.9871338228527, 
    0.98641579465316, 0.98568049532276, 0.98512078247392, 0.98439694615195, 
    0.98359166511314, 0.98242210368183, 0.98140733731502, 0.98053028742112, 
    0.97956048607535, 0.97881541023191, 0.97777409412689, 0.97601614774298, 
    0.97458209480607, 0.97298614726718, 0.9716026640998, 0.97046024058027, 
    0.96847737699537, 0.96650592286894, 0.96471613410032, 0.96226847579044, 
    0.95968962269252, 0.95714932074478, 0.95463591486036, 0.95144453229699, 
    0.94818095064323, 0.94457938626639, 0.94070436234657, 0.93601156790095, 
    0.93134997687419, 0.92605857862379, 0.91987712777245, 0.91402509273543, 
    0.90726806008898, 0.89846724170409, 0.88917747674806, 0.87980107292335, 
    0.86783646268962, 0.85423223798162, 0.83880817320503, 0.82306029986703, 
    0.80353445571152, 0.78124217288286, 0.75460919577636, 0.72450801145991, 
    0.68823961614694, 0.64742620506509, 0.6012573834425, 0.54964848617973, 
    0.48694843589671, 0.41442261667188, 0.33515614619954, 0.24716193528854, 
    0.16779802351098, 0.092256752563915, 0.035397671136877, 
    0.004012570050569, 0.0040996763047621, 0.036269515349152, 
    0.092186625190339, 0.16838547598462, 0.25284348068427, 0.336804920861, 
    0.41259642667422, 0.4780859200936, 0.54154999738539, 0.59941760685503, 
    0.6458655551883, 0.69037474368685, 0.72520483793784, 0.75146934999831, 
    0.77766128606983, 0.80124379023218, 0.82188649487062, 0.83860074236077, 
    0.85221423049393, 0.86741431403756, 0.87743724553472, 0.88753764071882, 
    0.89741503288349, 0.90577007921375, 0.91191134213783, 0.91882574607869, 
    0.92525422292393, 0.93066759160673, 0.93521448786831, 0.93946470895316, 
    0.94331334115045, 0.94737216431323, 0.95055342383536, 0.95380048422737, 
    0.95669012349801, 0.95915106219483, 0.96144116655454, 0.96420738247801, 
    0.96602597768258, 0.96778365093929, 0.96945752259479, 0.97140984673438, 
    0.97307799860048, 0.97464114741455, 0.97598093676807, 0.97712409336619, 
    0.97817181934209, 0.97902502832653, 0.98043770399305, 0.98160683486367, 
    0.98254975808182, 0.9833708317613, 0.98395651686481, 0.98482043394135, 
    0.98572777131236, 0.98660373786136, 0.98727142699303, 0.98773645875769, 
    0.9884208216228, 0.98892834020731, 0.98938126147443, 0.99007101192119, 
    0.99076055801876, 0.99116713749647, 0.99157108681238, 0.99192951565953, 
    0.99240652273728, 0.99277698221134, 0.99320158821218, 0.99358606847768, 
    0.99389916280029, 0.99424031746531, 0.99458179196175, 0.99490477276149, 
    0.99521967130767, 0.99547772834799, 0.99573022756059, 0.99598084004738, 
    0.99632284936365, 0.99653984186391, 0.99671751903242, 0.99694415837548, 
    0.99716122390651, 0.99738343503565, 0.99761386501404, 0.99779993204343, 
    0.9979813243673, 0.99814681630827, 0.99831557083546, 0.99850577310181, 
    0.9986720582496, 0.99880757025547, 0.99896656929575, 0.99912912594094, 
    0.99927574109212, 0.99941347396273, 0.99954556492817, 0.99967452508973, 
    0.99980260336384, 0.99992903883553,
  0.99993616794442, 0.99982416241219, 0.99970863572389, 0.99959063530027, 
    0.99946828549134, 0.9993424267662, 0.99921258799721, 0.99907753365828, 
    0.99893958855563, 0.99879431728542, 0.99864644354458, 0.99849156443466, 
    0.99833431674652, 0.99816638245592, 0.997995080226, 0.99781531537868, 
    0.99763614097847, 0.99744092241792, 0.99723822991539, 0.99704107137049, 
    0.99682353976249, 0.99659768543105, 0.99636716650127, 0.99613054881382, 
    0.99587676486721, 0.9956262004352, 0.99535056878272, 0.99506851093925, 
    0.994773406195, 0.99446911092087, 0.99417788721578, 0.99381621196864, 
    0.99348916631923, 0.99311465448863, 0.99275199974354, 0.99235966805813, 
    0.99194012240768, 0.99151720564045, 0.99106495503959, 0.99058841606272, 
    0.99009587646996, 0.98960031055434, 0.98903476520802, 0.98846422469976, 
    0.98781964136421, 0.98724736052263, 0.98657513802386, 0.98583399190061, 
    0.98509959761935, 0.98431038053814, 0.98345882474181, 0.98259009814546, 
    0.98165832295674, 0.98064033964847, 0.97961998063328, 0.97842500294461, 
    0.97722937289086, 0.97588395973101, 0.97456572282459, 0.97305525143303, 
    0.97152891023878, 0.96978786170222, 0.96791394709428, 0.96591861022307, 
    0.96373954331952, 0.96149386760364, 0.9589007012078, 0.95605195367172, 
    0.95329133738176, 0.94978148853016, 0.94620869285587, 0.9422039411448, 
    0.93793447441963, 0.93317049203755, 0.92783785427859, 0.92203553707268, 
    0.91519080109964, 0.9078480621319, 0.89967780089661, 0.89018213699863, 
    0.87944070973267, 0.86760393226753, 0.85379079406412, 0.83761979519443, 
    0.81990690675414, 0.79794161735642, 0.77421191090244, 0.74536200900562, 
    0.71129399012334, 0.67244767029575, 0.62619705736385, 0.57349884523771, 
    0.50932288956741, 0.43835026556203, 0.35776200987955, 0.27064317157705, 
    0.18487143421342, 0.10291025332355, 0.03913533439792, 0.0047755192643044, 
    0.0045620759314443, 0.040433030245144, 0.10139276841909, 
    0.18377472950177, 0.27097931623999, 0.35681632403716, 0.4361839132831, 
    0.50825637089003, 0.57151068603004, 0.62378900269835, 0.67087272679191, 
    0.7093483041676, 0.74245955852324, 0.77214722077072, 0.7961672132621, 
    0.81773852870337, 0.83517968155146, 0.85187646407407, 0.86539970689042, 
    0.87760945071221, 0.88857064760126, 0.89803176446362, 0.90632421878046, 
    0.91370382782736, 0.92058955959132, 0.9262903444513, 0.93189487351331, 
    0.93682364715797, 0.94132422942483, 0.94530545210795, 0.94881896723385, 
    0.9521728280102, 0.9553118605214, 0.95816844379372, 0.9606019367339, 
    0.96307708166235, 0.96532283309786, 0.96734601815519, 0.96926285265531, 
    0.97105958632046, 0.97256133154367, 0.97410803605982, 0.97561649532062, 
    0.97686805993507, 0.97815967907038, 0.97930871683066, 0.98039445056952, 
    0.98142866329534, 0.98243456533472, 0.98331257639261, 0.98419861631697, 
    0.98495909462929, 0.98577901597388, 0.98650112684112, 0.98716315736269, 
    0.98783309750262, 0.98844078781356, 0.98902241444038, 0.98961034827295, 
    0.9900978903248, 0.99061668650593, 0.99111079853795, 0.99154379820954, 
    0.99199564371096, 0.99241740494837, 0.99280802865826, 0.99318700461644, 
    0.99354124843992, 0.99389731181366, 0.9942290646434, 0.99453779134226, 
    0.99483933275459, 0.99512245044883, 0.99541494190483, 0.99567905462782, 
    0.99592875462804, 0.99619193761704, 0.99641089860863, 0.99664190641642, 
    0.99686316118038, 0.99707272610568, 0.99727851483158, 0.99746775695041, 
    0.99765877833896, 0.99783767014183, 0.99801172867442, 0.99818213205647, 
    0.99834307006036, 0.99850145593447, 0.9986516308661, 0.99880090889788, 
    0.99894092935893, 0.99908024209519, 0.999211150257, 0.9993428553106, 
    0.99946731170738, 0.99959004529889, 0.9997082650238, 0.99982365326197, 
    0.99993606661189 ;

 ens_sizes = 5, 6, 7, 8, 9, 10, 12, 14, 15, 16, 18, 20, 22, 24, 28, 30, 32, 
    36, 40, 44, 48, 49, 50, 52, 56, 60, 64, 70, 72, 80, 84, 88, 90, 96, 100, 
    120, 140, 160, 180, 200 ;
}
