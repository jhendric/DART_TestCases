netcdf pmo_input_member_0001 {
dimensions:
	domain_size = 40 ;
variables:
	double state(domain_size) ;
		state:units = "none" ;
	int dart_days ;
		dart_days:long_name = "days" ;
		dart_days:calendar = "no calendar" ;
		dart_days:units = "days since 0000-00-00 00:00:00" ;
	int dart_seconds ;
		dart_seconds:long_name = "seconds" ;
		dart_seconds:calendar = "no calendar" ;
		dart_seconds:units = "seconds since midnight" ;

// global attributes:
		:DART_file_information = "pmo_output member 0001" ;
		:DART_creation_date = "YYYY MM DD HH MM SS = 2016 11 18 11 16 27" ;
		:DART_source = "$URL: https://svn-dares-dart.cgd.ucar.edu/DART/branches/rma_fixed_filenames/io/direct_netcdf_mod.f90 $" ;
		:DART_revision = "$Revision: 10764 $" ;
		:DART_revdate = "$Date: 2016-11-18 09:03:39 -0700 (Fri, 18 Nov 2016) $" ;
data:

 state = -3.28383139922584, 2.98704435990934, 4.55877380586871, 
    6.15959210780279, -0.281343330323014, 1.78387200717577, 5.31530936897607, 
    6.18557938209699, -4.47093827823083, 5.08970322698255, 4.98419785217518, 
    3.00529335030821, 6.07878439203022, 4.0238500054969, 1.12271717800905, 
    3.89024750883235, 3.43764594930604, -1.95564593185033, 2.39194147665145, 
    3.41560530024931, 7.62619228013192, -2.55495233111732, -1.0108023620781, 
    1.59247191413994, 3.29985732255473, 4.19214385497745, 5.57756946998301, 
    -3.39854453293347, -0.435493083918519, -1.80144058187616, 
    8.64152948040963, 1.36741791127309, 1.39710986155821, 1.83257243925778, 
    3.6134909515423, 7.87047194181955, 0.90080119522991, 2.40795732830126, 
    5.75681171165689, 5.79527934521291 ;

 dart_days = 41 ;

 dart_seconds = 57600 ;
}
