netcdf Posterior_Diag {
dimensions:
	metadatalength = 64 ;
	locationrank = 1 ;
	copy = 24 ;
	time = UNLIMITED ; // (200 currently)
	NMLlinelen = 129 ;
	NMLnlines = 200 ;
	StateVariable = 1 ;
variables:
	int copy(copy) ;
		copy:long_name = "ensemble member or copy" ;
		copy:units = "nondimensional" ;
		copy:valid_range = 1, 24 ;
	char CopyMetaData(copy, metadatalength) ;
		CopyMetaData:long_name = "Metadata for each copy/member" ;
	char inputnml(NMLnlines, NMLlinelen) ;
		inputnml:long_name = "input.nml contents" ;
	double time(time) ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:cartesian_axis = "T" ;
		time:calendar = "no calendar" ;
		time:units = "days since 0000-00-00 00:00:00" ;
	double loc1d(StateVariable) ;
		loc1d:long_name = "location on unit circle" ;
		loc1d:dimension = 1 ;
		loc1d:units = "nondimensional" ;
		loc1d:valid_range = 0., 1. ;
	int StateVariable(StateVariable) ;
		StateVariable:long_name = "State Variable ID" ;
		StateVariable:units = "indexical" ;
		StateVariable:valid_range = 1, 1 ;
	double state(time, copy, StateVariable) ;
		state:long_name = "model state or fcopy" ;

// global attributes:
		:title = "posterior ensemble state" ;
		:assim_model_source = "$URL: https://proxy.subversion.ucar.edu/DAReS/DART/releases/Kodiak/assim_model/assim_model_mod.f90 $" ;
		:assim_model_revision = "$Revision: 4933 $" ;
		:assim_model_revdate = "$Date: 2011-06-01 11:55:44 -0600 (Wed, 01 Jun 2011) $" ;
		:creation_date = "YYYY MM DD HH MM SS = 2012 06 03 13 24 51" ;
		:model_source = "$URL: https://proxy.subversion.ucar.edu/DAReS/DART/releases/Kodiak/models/lorenz_63/model_mod.f90 $" ;
		:model_revision = "$Revision: 4933 $" ;
		:model_revdate = "$Date: 2011-06-01 11:55:44 -0600 (Wed, 01 Jun 2011) $" ;
		:model = "Lorenz_63" ;
		:model_r = 28. ;
		:model_b = 2.6666666666667 ;
		:model_sigma = 10. ;
		:model_deltat = 0.01 ;
data:

 copy = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24 ;

 CopyMetaData =
  "ensemble mean                                                   ",
  "ensemble spread                                                 ",
  "ensemble member      1                                          ",
  "ensemble member      2                                          ",
  "ensemble member      3                                          ",
  "ensemble member      4                                          ",
  "ensemble member      5                                          ",
  "ensemble member      6                                          ",
  "ensemble member      7                                          ",
  "ensemble member      8                                          ",
  "ensemble member      9                                          ",
  "ensemble member     10                                          ",
  "ensemble member     11                                          ",
  "ensemble member     12                                          ",
  "ensemble member     13                                          ",
  "ensemble member     14                                          ",
  "ensemble member     15                                          ",
  "ensemble member     16                                          ",
  "ensemble member     17                                          ",
  "ensemble member     18                                          ",
  "ensemble member     19                                          ",
  "ensemble member     20                                          ",
  "inflation mean                                                  ",
  "inflation sd                                                    " ;

 inputnml =
  "&perfect_model_obs_nml                                                                                                           ",
  "   start_from_restart    = .false.,                                                                                              ",
  "   output_restart        = .true.,                                                                                               ",
  "   async                 = 2,                                                                                                    ",
  "   init_time_days        = 0,                                                                                                    ",
  "   init_time_seconds     = 0,                                                                                                    ",
  "   first_obs_days        = -1,                                                                                                   ",
  "   first_obs_seconds     = -1,                                                                                                   ",
  "   last_obs_days         = -1,                                                                                                   ",
  "   last_obs_seconds      = -1,                                                                                                   ",
  "   output_interval       = 1,                                                                                                    ",
  "   restart_in_file_name  = \"perfect_ics\",                                                                                        ",
  "   restart_out_file_name = \"perfect_restart\",                                                                                    ",
  "   obs_seq_in_file_name  = \"obs_seq.in\",                                                                                         ",
  "   obs_seq_out_file_name = \"obs_seq.out\",                                                                                        ",
  "   adv_ens_command       = \"./advance_model.ksh\",                                                                                ",
  "   output_timestamps     = .false.,                                                                                              ",
  "   trace_execution       = .false.,                                                                                              ",
  "   output_forward_op_errors = .false.,                                                                                           ",
  "   print_every_nth_obs   = -1,                                                                                                   ",
  "   silence               = .false.,                                                                                              ",
  "  /                                                                                                                              ",
  "                                                                                                                                 ",
  "&filter_nml                                                                                                                      ",
  "   async                    = 2,                                                                                                 ",
  "   adv_ens_command          = \"./advance_model.ksh\",                                                                             ",
  "   ens_size                 = 20,                                                                                                ",
  "   start_from_restart       = .false.,                                                                                           ",
  "   output_restart           = .true.,                                                                                            ",
  "   obs_sequence_in_name     = \"obs_seq.out\",                                                                                     ",
  "   obs_sequence_out_name    = \"obs_seq.final\",                                                                                   ",
  "   restart_in_file_name     = \"perfect_ics\",                                                                                     ",
  "   restart_out_file_name    = \"filter_restart\",                                                                                  ",
  "   init_time_days           = 0,                                                                                                 ",
  "   init_time_seconds        = 0,                                                                                                 ",
  "   first_obs_days           = -1,                                                                                                ",
  "   first_obs_seconds        = -1,                                                                                                ",
  "   last_obs_days            = -1,                                                                                                ",
  "   last_obs_seconds         = -1,                                                                                                ",
  "   num_output_state_members = 20,                                                                                                ",
  "   num_output_obs_members   = 0,                                                                                                 ",
  "   output_interval          = 1,                                                                                                 ",
  "   num_groups               = 1,                                                                                                 ",
  "   input_qc_threshold       =  3.0,                                                                                              ",
  "   outlier_threshold        = -1.0,                                                                                              ",
  "   output_forward_op_errors = .false.,                                                                                           ",
  "   output_timestamps        = .false.,                                                                                           ",
  "   output_inflation         = .true.,                                                                                            ",
  "   trace_execution          = .false.,                                                                                           ",
  "   silence                  = .false.,                                                                                           ",
  "                                                                                                                                 ",
  "   inf_flavor                  = 0,                       0,                                                                     ",
  "   inf_initial_from_restart    = .false.,                 .false.,                                                               ",
  "   inf_sd_initial_from_restart = .false.,                 .false.,                                                               ",
  "   inf_output_restart          = .true.,                  .true.,                                                                ",
  "   inf_deterministic           = .true.,                  .true.,                                                                ",
  "   inf_in_file_name            = \'prior_inflate_ics\',     \'post_inflate_ics\',                                                    ",
  "   inf_out_file_name           = \'prior_inflate_restart\', \'post_inflate_restart\',                                                ",
  "   inf_diag_file_name          = \'prior_inflate_diag\',    \'post_inflate_diag\',                                                   ",
  "   inf_initial                 = 1.0,                     1.0,                                                                   ",
  "   inf_sd_initial              = 0.0,                     0.0,                                                                   ",
  "   inf_damping                 = 1.0,                     1.0,                                                                   ",
  "   inf_lower_bound             = 1.0,                     1.0,                                                                   ",
  "   inf_upper_bound             = 1000000.0,               1000000.0,                                                             ",
  "   inf_sd_lower_bound          = 0.0,                     0.0                                                                    ",
  "/                                                                                                                                ",
  "                                                                                                                                 ",
  "&smoother_nml                                                                                                                    ",
  "   num_lags              = 0,                                                                                                    ",
  "   start_from_restart    = .false.,                                                                                              ",
  "   output_restart        = .false.,                                                                                              ",
  "   restart_in_file_name  = \'smoother_ics\',                                                                                       ",
  "   restart_out_file_name = \'smoother_restart\'  /                                                                                 ",
  "                                                                                                                                 ",
  "&ensemble_manager_nml                                                                                                            ",
  "   single_restart_file_in  = .true.,                                                                                             ",
  "   single_restart_file_out = .true.,                                                                                             ",
  "   perturbation_amplitude  = 0.5  /                                                                                              ",
  "                                                                                                                                 ",
  "&assim_tools_nml                                                                                                                 ",
  "   filter_kind                     = 1,                                                                                          ",
  "   cutoff                          = 0.00001,                                                                                    ",
  "   sort_obs_inc                    = .true.,                                                                                     ",
  "   spread_restoration              = .false.,                                                                                    ",
  "   sampling_error_correction       = .false.,                                                                                    ",
  "   adaptive_localization_threshold = -1,                                                                                         ",
  "   output_localization_diagnostics = .false.,                                                                                    ",
  "   localization_diagnostics_file   = \'localization_diagnostics\',                                                                 ",
  "   print_every_nth_obs             = 0  /                                                                                        ",
  "                                                                                                                                 ",
  "&cov_cutoff_nml                                                                                                                  ",
  "   select_localization = 1  /                                                                                                    ",
  "                                                                                                                                 ",
  "&reg_factor_nml                                                                                                                  ",
  "   select_regression    = 1,                                                                                                     ",
  "   input_reg_file       = \"time_mean_reg\",                                                                                       ",
  "   save_reg_diagnostics = .false.,                                                                                               ",
  "   reg_diagnostics_file = \"reg_diagnostics\"  /                                                                                   ",
  "                                                                                                                                 ",
  "&obs_sequence_nml                                                                                                                ",
  "   write_binary_obs_sequence = .false.  /                                                                                        ",
  "                                                                                                                                 ",
  "&obs_kind_nml                                                                                                                    ",
  "   assimilate_these_obs_types = \'RAW_STATE_VARIABLE\'  /                                                                          ",
  "                                                                                                                                 ",
  "&assim_model_nml                                                                                                                 ",
  "   write_binary_restart_files = .false.,                                                                                         ",
  "   netCDF_large_file_support  = .false.                                                                                          ",
  "  /                                                                                                                              ",
  "                                                                                                                                 ",
  "&model_nml                                                                                                                       ",
  "   sigma  = 10.0,                                                                                                                ",
  "   r      = 28.0,                                                                                                                ",
  "   b      = 2.6666666666667,                                                                                                     ",
  "   deltat = 0.01,                                                                                                                ",
  "   time_step_days = 1,                                                                                                           ",
  "   time_step_seconds = 0  /                                                                                                      ",
  "                                                                                                                                 ",
  "&utilities_nml                                                                                                                   ",
  "   TERMLEVEL = 1,                                                                                                                ",
  "   module_details = .false.,                                                                                                     ",
  "   logfilename = \'dart_log.out\',                                                                                                 ",
  "   nmlfilename = \'dart_log.nml\',                                                                                                 ",
  "   write_nml   = \'terminal\'  /                                                                                                   ",
  "                                                                                                                                 ",
  "&preprocess_nml                                                                                                                  ",
  "    input_obs_def_mod_file = \'../../../obs_def/DEFAULT_obs_def_mod.F90\',                                                         ",
  "   output_obs_def_mod_file = \'../../../obs_def/obs_def_mod.f90\',                                                                 ",
  "   input_obs_kind_mod_file = \'../../../obs_kind/DEFAULT_obs_kind_mod.F90\',                                                       ",
  "  output_obs_kind_mod_file = \'../../../obs_kind/obs_kind_mod.f90\',                                                               ",
  "               input_files = \'../../../obs_def/obs_def_1d_state_mod.f90\'  /                                                      ",
  "                                                                                                                                 ",
  "                                                                                                                                 ",
  "&obs_sequence_tool_nml                                                                                                           ",
  "   num_input_files   = 2,                                                                                                        ",
  "   filename_seq      = \'obs_seq.one\', \'obs_seq.two\',                                                                             ",
  "   filename_out      = \'obs_seq.processed\',                                                                                      ",
  "   first_obs_days    = -1,                                                                                                       ",
  "   first_obs_seconds = -1,                                                                                                       ",
  "   last_obs_days     = -1,                                                                                                       ",
  "   last_obs_seconds  = -1,                                                                                                       ",
  "   print_only        = .false.,                                                                                                  ",
  "   gregorian_cal     = .false.                                                                                                   ",
  "   /                                                                                                                             ",
  "                                                                                                                                 ",
  "# other possible obs tool namelist items:                                                                                        ",
  "#                                                                                                                                ",
  "# keep only the U and V radiosonde winds:                                                                                        ",
  "#   obs_types          = \'RADIOSONDE_U_WIND_COMPONENT\',                                                                          ",
  "#                        \'RADIOSONDE_V_WIND_COMPONENT\',                                                                          ",
  "#   keep_types         = .true.,                                                                                                 ",
  "#                                                                                                                                ",
  "# remove the U and V radiosonde winds:                                                                                           ",
  "#   obs_types          = \'RADIOSONDE_U_WIND_COMPONENT\',                                                                          ",
  "#                        \'RADIOSONDE_V_WIND_COMPONENT\',                                                                          ",
  "#   keep_types         = .false.,                                                                                                ",
  "#                                                                                                                                ",
  "# keep only observations with a DART QC of 0:                                                                                    ",
  "#   qc_metadata        = \'Dart quality control\',                                                                                 ",
  "#   min_qc             = 0,                                                                                                      ",
  "#   max_qc             = 0,                                                                                                      ",
  "#                                                                                                                                ",
  "# keep only radiosonde temp obs between 250 and 300 K:                                                                           ",
  "#   copy_metadata      = \'NCEP BUFR observation\',                                                                                ",
  "#   copy_type          = \'RADIOSONDE_TEMPERATURE\',                                                                               ",
  "#   min_copy           = 250.0,                                                                                                  ",
  "#   max_copy           = 300.0,                                                                                                  ",
  "#                                                                                                                                ",
  "                                                                                                                                 ",
  "                                                                                                                                 ",
  "&restart_file_tool_nml                                                                                                           ",
  "   input_file_name              = \"filter_restart\",                                                                              ",
  "   output_file_name             = \"filter_updated_restart\",                                                                      ",
  "   ens_size                     = 1,                                                                                             ",
  "   single_restart_file_in       = .true.,                                                                                        ",
  "   single_restart_file_out      = .true.,                                                                                        ",
  "   write_binary_restart_files   = .true.,                                                                                        ",
  "   overwrite_data_time          = .false.,                                                                                       ",
  "   new_data_days                = -1,                                                                                            ",
  "   new_data_secs                = -1,                                                                                            ",
  "   input_is_model_advance_file  = .false.,                                                                                       ",
  "   output_is_model_advance_file = .false.,                                                                                       ",
  "   overwrite_advance_time       = .false.,                                                                                       ",
  "   new_advance_days             = -1,                                                                                            ",
  "   new_advance_secs             = -1,                                                                                            ",
  "   gregorian_cal                = .false.                                                                                        ",
  "/                                                                                                                                ",
  "                                                                                                                                 ",
  "&obs_diag_nml                                                                                                                    ",
  "   obs_sequence_name  = \'obs_seq.final\',                                                                                         ",
  "   iskip_days         = 0,                                                                                                       ",
  "   obs_select         = 1,                                                                                                       ",
  "   rat_cri            = 4.0,                                                                                                     ",
  "   input_qc_threshold = 3.0,                                                                                                     ",
  "   bin_width_seconds = 0,                                                                                                        ",
  "   lonlim1   = 0.0, 0.0, 0.5, -1.0,                                                                                              ",
  "   lonlim2   = 1.0, 0.5, 1.5, -1.0,                                                                                              ",
  "   reg_names = \'whole\', \'yin\', \'yang\', \'bogus\',                                                                                  ",
  "   verbose   = .false.  /                                                                                                        ",
  "                                                                                                                                 " ;

 time = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 107, 
    108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 121, 
    122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 
    136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 149, 
    150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 
    164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 177, 
    178, 179, 180, 181, 182, 183, 184, 185, 186, 187, 188, 189, 190, 191, 
    192, 193, 194, 195, 196, 197, 198, 199, 200 ;

 loc1d = 0 ;

 StateVariable = 1 ;

 state =
  -77.4417879203855,
  0.289858816773224,
  -77.3719792673194,
  -77.066952930688,
  -77.3848416764962,
  -77.0638814066748,
  -77.490827457118,
  -78.041477025344,
  -77.2747855499996,
  -77.7592746634996,
  -77.7363916977634,
  -77.9278868162742,
  -77.2728340368974,
  -77.8293313423879,
  -77.2640117988257,
  -77.2325394853575,
  -77.5563304121142,
  -77.0658982245246,
  -77.5078661955036,
  -77.4926044146548,
  -77.2316813783518,
  -77.2643626279141,
  1,
  0,
  -77.3435068222765,
  0.276932963622954,
  -76.752488168745,
  -77.4076650491113,
  -77.3585873586531,
  -77.2212576065384,
  -77.3964542305478,
  -77.77989340311,
  -76.8319211828801,
  -77.5123798762732,
  -77.5872527195869,
  -77.319373358156,
  -76.9653779837115,
  -77.344376186094,
  -77.0997894549077,
  -77.5868174180175,
  -77.6483490023437,
  -77.3061295197595,
  -77.4251570118043,
  -77.6980357727656,
  -77.1483909074553,
  -77.4804402350691,
  1,
  0,
  -77.3188878920056,
  0.267589588827667,
  -76.8143596533116,
  -77.2278154334656,
  -77.3885898383173,
  -77.0351025037252,
  -77.0395001173535,
  -77.6524950449936,
  -77.5161947951363,
  -77.5507031124298,
  -77.5306912475655,
  -77.3363337255612,
  -77.2425702559209,
  -76.93670104881,
  -76.9529561071794,
  -77.2556849025569,
  -77.6102244839014,
  -77.1302136426932,
  -77.6564400856109,
  -77.549013501654,
  -77.3050986684366,
  -77.6470696714888,
  1,
  0,
  -77.4420358803461,
  0.251342685380029,
  -77.3326561543242,
  -77.5838791195958,
  -77.4402076503423,
  -76.8381513188308,
  -77.527136424921,
  -77.385447099469,
  -77.4505587768335,
  -77.5156795693324,
  -77.584705687237,
  -77.4256129888194,
  -77.3035970066318,
  -77.5156089058421,
  -77.010913573085,
  -77.4354908928257,
  -77.560434061439,
  -77.2418622123523,
  -78.0675045362038,
  -77.3434251037797,
  -77.7482896016703,
  -77.5295569233873,
  1,
  0,
  -78.0167712226106,
  0.284800168748313,
  -78.3409244644376,
  -77.9750693808697,
  -78.0751829347868,
  -77.680498939484,
  -77.9398851094283,
  -77.8494716852766,
  -78.2166999777074,
  -78.1816522291233,
  -77.9680988373805,
  -78.2219528173011,
  -77.3928789855697,
  -78.3395935238813,
  -77.4720640564996,
  -78.0669068404407,
  -78.2072036626488,
  -78.0860439920125,
  -78.0250605231901,
  -77.6958729761527,
  -78.493642298422,
  -78.1067212175993,
  1,
  0,
  -78.7600432625476,
  0.312264446525049,
  -78.988751932379,
  -78.4877661863549,
  -79.1850190232496,
  -78.5717177458594,
  -78.2374815843187,
  -78.5976213109195,
  -79.1750118678688,
  -78.7241965208683,
  -78.6916312468296,
  -78.8112350500633,
  -78.3389909597162,
  -79.3737682167103,
  -78.4700881157672,
  -78.5710253318184,
  -79.0350965197294,
  -78.7349026691725,
  -78.9075371535219,
  -78.4470167657105,
  -79.1552040824785,
  -78.6968029676157,
  1,
  0,
  -79.5569321671627,
  0.304627405702061,
  -79.4390505672494,
  -79.23979038414,
  -79.9575900097053,
  -78.9248782816824,
  -79.3781180039325,
  -79.4850813288607,
  -79.8361598001698,
  -79.7211225631142,
  -79.8368636597013,
  -79.8267856863564,
  -79.2527977314505,
  -79.6127645399361,
  -79.0814441257294,
  -79.488876169426,
  -80.156763760342,
  -79.4046424267438,
  -79.8430476173759,
  -79.4989369070707,
  -79.5826906143887,
  -79.5712391658788,
  1,
  0,
  -80.2626332921205,
  0.311477817703548,
  -80.0137260582428,
  -79.9963206246364,
  -80.0594003598037,
  -79.6597488327838,
  -80.4067588720868,
  -79.9057197505171,
  -80.7870633490283,
  -80.5238007236066,
  -80.4398570541022,
  -80.1720280697883,
  -80.1484763126414,
  -80.7170283936533,
  -80.3283007391754,
  -80.6944032021483,
  -80.5091165490073,
  -79.818155533328,
  -80.449881662584,
  -80.4096396052835,
  -80.126312475497,
  -80.0869276744961,
  1,
  0,
  -81.285876903475,
  0.331136721089038,
  -80.8947366765723,
  -81.2067440358726,
  -81.0846914153933,
  -80.8012071919675,
  -81.7535258778295,
  -80.8404684651537,
  -81.2851062385271,
  -81.8095513960717,
  -81.484380734681,
  -81.3176791000887,
  -81.2664204779543,
  -82.0189913055963,
  -81.4634659301884,
  -81.1804668906529,
  -81.6292699647001,
  -81.0532819413066,
  -81.1421036495681,
  -81.4150560067073,
  -81.0081122098815,
  -81.0622785607876,
  1,
  0,
  -82.2653042012421,
  0.316820127999305,
  -81.782011599861,
  -82.453616734364,
  -82.0272292889626,
  -81.7966351532789,
  -82.8885302824536,
  -82.3328815914734,
  -81.8820975163379,
  -82.4261186375151,
  -81.7825693994343,
  -82.2105048427819,
  -82.4946956247259,
  -82.8925919592994,
  -82.1395397154673,
  -82.2729721311817,
  -82.2912293380381,
  -82.1191510974544,
  -82.4248413883515,
  -82.4838048925945,
  -82.3077338907433,
  -82.2973289405242,
  1,
  0,
  -83.1786365438853,
  0.284657537879281,
  -82.9957865298759,
  -83.3687095513826,
  -83.0926777088326,
  -82.7596126532667,
  -83.9057884527846,
  -83.3609359967169,
  -82.9286788975589,
  -83.0229239729661,
  -83.0860657065153,
  -83.0041698725847,
  -83.3819664926879,
  -83.1556237891951,
  -83.1329339840571,
  -82.877073786366,
  -83.3658411739745,
  -82.8211950979763,
  -83.160186874638,
  -83.6663391158677,
  -83.0771273106669,
  -83.4090939097925,
  1,
  0,
  -84.0351513244424,
  0.330744355423971,
  -83.5786030221388,
  -83.9876045525517,
  -84.3283215466103,
  -83.8675404167309,
  -84.4885310970688,
  -84.6015575854808,
  -83.8661334119188,
  -83.9098077382962,
  -84.1206897802809,
  -83.5637468416529,
  -84.2928908278388,
  -83.6395916940705,
  -83.7896649552773,
  -83.7510452716335,
  -84.3909899970126,
  -83.6271686733814,
  -84.3686371349584,
  -84.4283708719462,
  -84.1740093034921,
  -83.9281217665077,
  1,
  0,
  -85.3093990395676,
  0.359600058263196,
  -84.6672271222524,
  -85.5664478482093,
  -85.8821880744157,
  -85.586201186148,
  -85.4533779099907,
  -85.3317853624729,
  -84.9454459331769,
  -84.9452444894088,
  -85.7351456497268,
  -85.271303376414,
  -85.663046424567,
  -85.0825379667749,
  -85.2368276180773,
  -85.1341866865446,
  -85.6844354212224,
  -84.5835323658149,
  -85.525729417367,
  -85.4625772724691,
  -84.9538602604156,
  -85.476880405883,
  1,
  0,
  -87.0680468642142,
  0.405136737620315,
  -86.8482244365158,
  -87.2440149051447,
  -87.7559853791898,
  -87.4296696763306,
  -87.215474198599,
  -86.7747358943827,
  -87.0456869145269,
  -86.8761516142855,
  -87.4354319277728,
  -87.0139874673693,
  -87.6340032833319,
  -86.3141885198576,
  -86.2856146655117,
  -87.2199265921332,
  -87.2855884529632,
  -86.4307898663085,
  -86.8035504466584,
  -87.3130785797201,
  -87.2040169948096,
  -87.2308174688725,
  1,
  0,
  -88.2192121829823,
  0.370846027287119,
  -87.3928669637747,
  -88.3571085858898,
  -88.2689618472559,
  -88.069653554419,
  -88.3417637951933,
  -88.1442855319669,
  -88.2045158711266,
  -88.5924552342399,
  -88.3143256437822,
  -88.2501365234556,
  -88.5494187498733,
  -87.5126161536469,
  -87.6862681712433,
  -88.7356337134302,
  -88.3179392252283,
  -88.1045920239257,
  -88.34454522707,
  -88.8485920902464,
  -88.4175491873028,
  -87.9310155665743,
  1,
  0,
  -88.7308440849555,
  0.323546710364468,
  -88.0985528185793,
  -88.7809451796063,
  -88.8218589574816,
  -88.1480829868936,
  -88.9925935135749,
  -88.7263394739696,
  -89.3357366932097,
  -89.3317861498367,
  -88.8419269024702,
  -88.6991556665608,
  -88.4909224428427,
  -88.6491967846254,
  -88.5423611799116,
  -88.9442017034154,
  -88.7940635552957,
  -88.4730733495731,
  -88.7560773729481,
  -88.7616098428047,
  -89.0397838745666,
  -88.3886132509447,
  1,
  0,
  -89.8890759406767,
  0.43334634947856,
  -89.6991387480609,
  -89.8640129143272,
  -89.9807096897793,
  -89.4476834627067,
  -90.0475317084991,
  -89.4648667633931,
  -90.614910370983,
  -90.8218003773635,
  -90.1128674172685,
  -89.9550293302764,
  -89.087228915025,
  -90.2400494599224,
  -89.2426881923943,
  -89.9455752629111,
  -89.8874208671623,
  -89.2697302850656,
  -89.9328363472264,
  -89.9566738358549,
  -90.127240465545,
  -90.0835243997689,
  1,
  0,
  -91.1486434203632,
  0.499487655341717,
  -90.8298378758942,
  -90.8964974611005,
  -91.4655620071978,
  -91.1771730461293,
  -91.0552496966859,
  -90.9862276983147,
  -91.985018902938,
  -91.8283228437488,
  -91.2123368879879,
  -91.3947065540919,
  -90.7267610388265,
  -91.8281460479081,
  -90.8736377499695,
  -90.6970697563177,
  -90.2142244069112,
  -90.130293166145,
  -91.3335411268827,
  -91.3639103360391,
  -91.2955457574798,
  -91.6788060466953,
  1,
  0,
  -92.0320730786009,
  0.476032491539692,
  -91.6477061794846,
  -91.8466246832122,
  -91.8835767540283,
  -92.0251095378768,
  -91.816769285495,
  -92.3117758494972,
  -93.0041296318018,
  -92.618367638955,
  -92.3103053302054,
  -91.990202990241,
  -91.3437552162073,
  -92.6571698367945,
  -92.0169218462546,
  -91.7732680071552,
  -90.997485941293,
  -91.4346569447112,
  -92.1272747252377,
  -92.4716208136465,
  -92.2174023365108,
  -92.1473380234109,
  1,
  0,
  -92.4087070066804,
  0.401167444574236,
  -92.1192853392045,
  -92.7122226070306,
  -92.7511571709,
  -92.5486600945438,
  -92.0496492945725,
  -92.6296310203099,
  -93.2035623628315,
  -92.6340591940597,
  -92.2637146920914,
  -92.0031015239257,
  -91.9277209323876,
  -93.3296201477299,
  -91.8505346828269,
  -92.1375339675783,
  -92.6803077031282,
  -92.0953007081841,
  -92.3710776688527,
  -92.2656651231597,
  -92.2072700950097,
  -92.3940658052803,
  1,
  0,
  -92.8103609366166,
  0.506722874780497,
  -92.9704903731832,
  -92.7693756005773,
  -93.0541643002851,
  -93.0555780810025,
  -92.7085984731262,
  -93.4083664148309,
  -93.5917822361414,
  -93.0977866804822,
  -91.5850866337701,
  -92.2233096040659,
  -92.7655799076428,
  -93.7855942959906,
  -92.8566164974368,
  -92.6399604226301,
  -92.7728074237549,
  -92.9532183271519,
  -92.5372493253797,
  -91.987087198951,
  -92.5632071920619,
  -92.881359743867,
  1,
  0,
  -93.0474542420966,
  0.519399919306764,
  -93.5037729454825,
  -92.4999255013532,
  -93.3196429970632,
  -93.3035988831933,
  -92.8865158120926,
  -93.7795431324912,
  -93.7062013172876,
  -93.4985362844753,
  -92.7040762130618,
  -92.6778059624185,
  -92.4799974005758,
  -94.2440827867768,
  -93.1316392953769,
  -92.5604578997891,
  -92.989695277921,
  -92.7908985613087,
  -92.5737333618879,
  -92.5825424860358,
  -92.3866728678573,
  -93.3297458554835,
  1,
  0,
  -92.9879120416694,
  0.568816147402591,
  -93.5883729611989,
  -92.8032356634133,
  -93.2968305579092,
  -93.2230059848153,
  -93.1881116993049,
  -93.3218420658196,
  -94.324404408981,
  -93.2469802248339,
  -92.721714973199,
  -92.6184609741111,
  -92.0403284299632,
  -93.9181646426736,
  -92.4758456018418,
  -92.3248834638363,
  -93.160439737973,
  -92.9037953788042,
  -92.4480890791823,
  -92.672692158817,
  -92.3076634827802,
  -93.1733793439292,
  1,
  0,
  -93.3213997939107,
  0.52451325330789,
  -94.0908479486529,
  -92.9925593482625,
  -93.5320790248078,
  -93.6540768946587,
  -93.3565929916402,
  -93.1147419691521,
  -94.1456437035687,
  -93.112865101497,
  -93.4008686415707,
  -93.2191889743517,
  -92.3060471009449,
  -93.6703486056093,
  -93.0908802089568,
  -92.6401846531282,
  -94.338353896025,
  -93.1370336431993,
  -92.424524783302,
  -93.5327564000797,
  -93.3132352085286,
  -93.3551667802772,
  1,
  0,
  -93.6329604513416,
  0.511448135484627,
  -94.4554034541069,
  -93.0081276867926,
  -93.7168975541398,
  -93.8637732215848,
  -93.9619599430962,
  -93.1797800694742,
  -93.9390260339061,
  -93.3068888627054,
  -93.6673409571999,
  -93.3958273059486,
  -92.4845514808615,
  -93.8061942069596,
  -93.5105916132763,
  -93.205189982423,
  -94.6092442571328,
  -93.5170454777991,
  -93.4726745841206,
  -94.237183726253,
  -94.0886133302811,
  -93.2328952787699,
  1,
  0,
  -93.5828869226736,
  0.53874109170709,
  -94.6364839893105,
  -93.2405832455627,
  -93.7317164337519,
  -93.9646901886466,
  -93.5653678083387,
  -92.9123207190501,
  -94.5148957936042,
  -93.1170053907083,
  -93.5740703298038,
  -93.2482246014944,
  -93.3772182975022,
  -93.9395166140558,
  -92.8561163449865,
  -93.0955483596312,
  -93.8730051244155,
  -93.7681005566545,
  -93.7212366607237,
  -94.206134913081,
  -93.7273987375721,
  -92.5881043445791,
  1,
  0,
  -92.9849365431669,
  0.680329625316594,
  -93.8088543348182,
  -92.675185328246,
  -93.1041878300504,
  -93.846366316323,
  -92.9511361702633,
  -91.7306712467414,
  -93.8924273468848,
  -93.0425526796034,
  -92.9047736688693,
  -92.0508886105797,
  -93.1462452811894,
  -93.3170590169817,
  -92.9008984021834,
  -92.678968396584,
  -93.3064723081054,
  -93.8784099084759,
  -93.2669808732109,
  -93.009492936881,
  -92.8601070512074,
  -91.3270531561399,
  1,
  0,
  -92.5170650238064,
  0.786534600609623,
  -93.6849860452238,
  -92.2781109674604,
  -92.9230410710991,
  -93.5789862211306,
  -92.3778928315213,
  -91.0109197439227,
  -93.4798296089368,
  -91.9030128626957,
  -92.8123475797746,
  -91.8066453859867,
  -93.1759878575699,
  -93.0006775167483,
  -91.848045448081,
  -92.2390008111668,
  -92.4823535258971,
  -93.3851810170118,
  -92.4832168161755,
  -92.9575866401409,
  -91.9390126023958,
  -90.9744659231895,
  1,
  0,
  -92.0598371637222,
  0.802414363473412,
  -93.4384143922775,
  -91.9313469655798,
  -92.4212561303176,
  -93.0423636013151,
  -91.7432107800116,
  -90.9648143381099,
  -92.807782690003,
  -91.3917361005275,
  -92.96061830282,
  -91.5946110425403,
  -92.6319859595285,
  -91.5288474452153,
  -91.7201322343324,
  -92.1571255190403,
  -91.952834412824,
  -93.2766221488961,
  -91.053462478535,
  -92.2864408868353,
  -91.8281658474057,
  -90.4649719983286,
  1,
  0,
  -91.720147897021,
  0.959680171547131,
  -93.7201784465194,
  -92.1350903019647,
  -91.5378332976697,
  -92.7929837859012,
  -91.9911921971193,
  -91.2197826837405,
  -93.2536846001295,
  -91.408305488817,
  -91.5770991978616,
  -90.4126037112332,
  -91.7593409333265,
  -90.7670636059327,
  -92.0721384482733,
  -91.9959154871557,
  -91.5906066208998,
  -92.4021371573675,
  -90.7058578533974,
  -92.1170067784772,
  -91.4063727499083,
  -89.5377645947254,
  1,
  0,
  -91.6533574203075,
  0.836340535279564,
  -93.4400075181097,
  -92.0603411406963,
  -91.8142579334988,
  -92.0581079243705,
  -91.5661105247345,
  -92.308317014158,
  -92.4953807037784,
  -91.1484143348606,
  -91.0662728108524,
  -90.7671207424355,
  -91.5660444939576,
  -90.711692674178,
  -92.3891699239472,
  -91.4732664206356,
  -91.159625761352,
  -92.5109009097906,
  -90.9197268770953,
  -92.2053133030217,
  -91.7324212303297,
  -89.674656164348,
  1,
  0,
  -91.244724004021,
  0.945757161455055,
  -93.5999584550325,
  -92.084014905668,
  -91.3775120083979,
  -91.1787355014396,
  -91.1532960370755,
  -91.7145376218606,
  -91.7423740323831,
  -90.9924179810204,
  -90.5721356570609,
  -89.9537524677517,
  -91.0655412690945,
  -90.3824220340555,
  -91.5721145948355,
  -91.1942500596595,
  -90.9339636573045,
  -92.4958651086549,
  -90.1636237171655,
  -91.7462034284353,
  -91.6988305947418,
  -89.2729309487819,
  1,
  0,
  -91.1571213284126,
  1.03122395072777,
  -93.2737120271085,
  -91.7102027873135,
  -92.0547037711005,
  -91.2847938810089,
  -91.645944066812,
  -91.4097620718532,
  -91.5443309994272,
  -91.3814060800533,
  -90.6374335769658,
  -89.7539950468292,
  -90.4156347948377,
  -90.2241124668913,
  -90.8349792516131,
  -90.9043533181291,
  -90.9863643585791,
  -92.9637374129248,
  -90.627588633685,
  -91.7805661375051,
  -91.0608734279121,
  -88.647932457702,
  1,
  0,
  -91.1828498149771,
  1.20389661890764,
  -93.5229263342552,
  -91.7950110695484,
  -92.0040930452176,
  -91.1997801891093,
  -91.5109087356953,
  -91.5743708094384,
  -91.8133891270309,
  -91.2219685619959,
  -90.2474495838444,
  -88.8871808358422,
  -90.4224801054899,
  -90.3674666020474,
  -91.1529389257137,
  -90.8930920013813,
  -91.1938813479404,
  -93.1541328777448,
  -90.6926234646143,
  -91.9687326991533,
  -91.6632642410032,
  -88.3713057424764,
  1,
  0,
  -91.2477271317524,
  1.17780813768825,
  -93.4851906881043,
  -92.1609748965511,
  -92.1553493024725,
  -91.7811798053003,
  -91.4838189208934,
  -91.4708054016878,
  -91.2616695304971,
  -91.1469601075097,
  -89.9389911190607,
  -89.4036015549424,
  -90.5095862184757,
  -89.7438505546396,
  -90.8857600014714,
  -90.9638472304611,
  -91.6159279977834,
  -93.2628454602708,
  -90.6538388329001,
  -92.6774840045518,
  -91.2424308701869,
  -89.1104301372882,
  1,
  0,
  -91.5453718792286,
  1.28737570197909,
  -93.9995531700574,
  -91.8861771925324,
  -92.2502720369056,
  -91.7573810846028,
  -91.6417490756,
  -91.8577416897247,
  -92.1438572740997,
  -91.5591934952254,
  -90.361300790055,
  -89.2509570789981,
  -90.8497898014997,
  -90.3941657284019,
  -91.5216590090172,
  -90.9317566009723,
  -92.282690489199,
  -93.9400950861272,
  -90.617024492693,
  -92.969835195173,
  -91.6585454916067,
  -89.0336928020818,
  1,
  0,
  -90.9169603328278,
  1.31586333114255,
  -93.5958599119325,
  -92.0813980159602,
  -91.6412272159465,
  -90.2737565666174,
  -90.8904423880182,
  -92.1520119398532,
  -91.8947744107689,
  -90.8682832193686,
  -89.7787634285611,
  -89.6089501280404,
  -90.1473530540434,
  -88.9688352803959,
  -89.9770638047855,
  -90.8816615415761,
  -91.2803740894993,
  -93.2348870485095,
  -89.2833406102724,
  -91.7387207599383,
  -91.0718068415108,
  -88.9696964009571,
  1,
  0,
  -90.6016776949236,
  1.20116819565082,
  -93.5128299980851,
  -91.5762775700208,
  -91.2840574180449,
  -90.008744481035,
  -89.8921295039104,
  -91.2148420390812,
  -90.8890932886633,
  -91.017928001145,
  -90.0354777872319,
  -90.4961982195158,
  -90.1701469114528,
  -88.6641744217534,
  -89.3725035026952,
  -91.2748346971841,
  -90.4678583795049,
  -92.1394632168762,
  -89.0428827068196,
  -91.8987180963398,
  -90.2592632773953,
  -88.8161303817164,
  1,
  0,
  -90.4172363296271,
  1.14832566562483,
  -92.6824996960516,
  -91.099102271597,
  -91.1448658852002,
  -90.5492060197924,
  -88.9582480272211,
  -91.3012957963284,
  -91.1097068996961,
  -90.9591123835906,
  -89.1022279352261,
  -90.4169332479233,
  -90.2648355812163,
  -88.5095075246684,
  -89.9868440549568,
  -91.0708031404228,
  -89.8745006019685,
  -91.9121796239466,
  -88.8512596401136,
  -91.7575103837789,
  -89.8236011612077,
  -88.9704867176358,
  1,
  0,
  -90.1790498237717,
  1.04751879637327,
  -92.5541518713374,
  -90.7184090211609,
  -91.6049972290131,
  -89.7573831246987,
  -89.149022543567,
  -90.8152488788761,
  -90.2561500822966,
  -90.6999121642203,
  -88.7177443774389,
  -89.6221852992881,
  -90.2568181043341,
  -88.3804842154644,
  -89.9209447344788,
  -90.2985254060087,
  -89.9173909709831,
  -91.5872719695317,
  -89.4676754767893,
  -91.1224876184124,
  -89.8302451650479,
  -88.9039482224873,
  1,
  0,
  -89.5304637029681,
  0.939217589481229,
  -91.0937121305277,
  -89.556856715185,
  -90.838665323313,
  -88.5650684162206,
  -88.6083060293906,
  -89.9763858572493,
  -89.5160703187888,
  -90.5885637771675,
  -88.6066489211567,
  -89.2118855655908,
  -89.4547086122383,
  -88.1411772906887,
  -89.2530671828553,
  -89.2942088465901,
  -90.1109555722297,
  -91.4577730247931,
  -89.3842144698722,
  -89.9073349823611,
  -88.8613328214073,
  -88.1823382017355,
  1,
  0,
  -88.1674849578179,
  0.804409671056297,
  -89.4326853026922,
  -87.669719359822,
  -89.7429256434035,
  -87.6706105170859,
  -87.0300962201781,
  -88.649929525975,
  -88.0502021763585,
  -89.1366502436692,
  -88.1407569642982,
  -87.9938085796914,
  -87.604081796834,
  -87.5487548487899,
  -87.5988181840129,
  -88.1537814509062,
  -88.0178200339576,
  -89.6752597648926,
  -87.5820799985727,
  -88.7460693854642,
  -87.7595500162395,
  -87.146099143515,
  1,
  0,
  -87.2156060204776,
  0.720295318376311,
  -87.9015362584322,
  -87.1654130301594,
  -89.0713681040618,
  -87.3584075022323,
  -85.9023286054169,
  -87.6618427791139,
  -87.7135532201327,
  -87.4841415960983,
  -87.3679979475759,
  -86.6259323854283,
  -86.656320240622,
  -86.9042418088326,
  -86.2089012785152,
  -86.702035574912,
  -86.8429608050282,
  -88.1677430365619,
  -87.0095130450876,
  -87.7808377600292,
  -86.8501194101055,
  -86.9369260212066,
  1,
  0,
  -86.8216535419466,
  0.738209111377905,
  -86.9362141371183,
  -86.4835205534204,
  -88.609189820612,
  -86.5081346324693,
  -85.2150962050075,
  -86.8736222875301,
  -86.8690271379073,
  -86.4265385082835,
  -87.5197995215863,
  -86.3717609576265,
  -86.1216557862253,
  -86.6237384175398,
  -86.5162469936979,
  -86.659405647551,
  -86.2239334126723,
  -87.9587286340567,
  -86.5966135125109,
  -87.7906916828495,
  -87.2819351387713,
  -86.8472178514955,
  1,
  0,
  -85.0563586254005,
  0.649409294434984,
  -84.9032495005187,
  -84.7011783383513,
  -86.202262433689,
  -84.952463422679,
  -83.5284314314189,
  -85.3488465601337,
  -85.1520547143403,
  -84.4556374565112,
  -85.3925901078732,
  -84.7303676788353,
  -84.3032428073557,
  -85.1313327830299,
  -84.6051770828642,
  -84.6754714198703,
  -84.66688255142,
  -86.118399121532,
  -85.1587128634412,
  -85.9110145184979,
  -85.6576983822197,
  -85.532159333428,
  1,
  0,
  -83.472886332724,
  0.61909207981525,
  -83.543708162897,
  -83.1631718706932,
  -84.9801210629077,
  -83.2227322101816,
  -82.2750314484814,
  -83.4676444540973,
  -83.5924874206867,
  -83.603377446262,
  -83.6063123768191,
  -83.1730318755509,
  -82.5042515985731,
  -82.8583883591931,
  -83.5317103832341,
  -83.3749110370499,
  -82.7089273549334,
  -83.8345261165462,
  -83.8750398309458,
  -84.221641825214,
  -84.08698296044,
  -83.8337288597731,
  1,
  0,
  -82.9298146021312,
  0.534870902038586,
  -83.1586434036563,
  -82.5250745856322,
  -84.0857043873054,
  -82.8196213151525,
  -82.1120030107105,
  -83.1333846137833,
  -83.2325961230684,
  -83.1074886832127,
  -82.7826399599654,
  -82.4375497309637,
  -82.2194928290074,
  -82.4305345166729,
  -82.4240236137797,
  -83.0218409954702,
  -82.2853330949908,
  -83.208188536398,
  -83.432260302455,
  -83.8841697278236,
  -83.1949947362916,
  -83.1007478762848,
  1,
  0,
  -82.4804596108752,
  0.541954705635225,
  -82.1091005743637,
  -81.8922071778654,
  -83.4722446285837,
  -82.9803720273307,
  -81.6053708434872,
  -82.7119159622424,
  -82.7123095039162,
  -82.6525097446467,
  -82.5640794017646,
  -82.0163846086268,
  -81.9298030681713,
  -81.8961010257664,
  -81.8490349253024,
  -82.5235528379723,
  -81.9779770903969,
  -82.7894313496913,
  -82.7490804708465,
  -83.4614512449656,
  -82.9700233698127,
  -82.7462423617517,
  1,
  0,
  -82.3837120790225,
  0.51894397704842,
  -82.2527225605404,
  -81.9439495531622,
  -82.893741223573,
  -82.5607136860487,
  -81.9102057909624,
  -82.5301326062835,
  -82.7230777323879,
  -82.3105164484187,
  -82.3628295631687,
  -81.8942299824198,
  -81.5480914883704,
  -81.7060752094565,
  -81.5871403332705,
  -82.8263896320054,
  -82.1155104304229,
  -82.878973828548,
  -82.7630207049298,
  -83.5634455932233,
  -82.7614225398358,
  -82.5420526734213,
  1,
  0,
  -82.7009914508249,
  0.478522750302106,
  -82.0655513889751,
  -82.2389299530822,
  -83.258055870439,
  -82.8815320243287,
  -81.9450932293884,
  -83.0237450284898,
  -83.075384466196,
  -82.4247779565547,
  -83.2002782437266,
  -82.4034955884107,
  -81.9258749588941,
  -82.2997457943595,
  -82.1503104103599,
  -83.4155538539972,
  -82.9763142336052,
  -82.6477805926849,
  -82.8351755427132,
  -83.2469526008122,
  -82.9380590962676,
  -83.0672181832123,
  1,
  0,
  -82.4207302979028,
  0.424270658766876,
  -81.9330504311246,
  -81.8233044508154,
  -82.8620258322653,
  -82.2389805072986,
  -81.6563262765157,
  -82.5221771300126,
  -82.5724283654475,
  -82.4514937735681,
  -83.106049139213,
  -82.6224618845659,
  -81.9171677873088,
  -82.161045699379,
  -81.7265916273052,
  -82.5579094708038,
  -82.785689520883,
  -82.5621556849926,
  -82.5025713041227,
  -82.6904482930881,
  -82.9754787310888,
  -82.7472500482581,
  1,
  0,
  -83.2098210361415,
  0.441108842209545,
  -82.6974699529354,
  -82.6202217123319,
  -83.505284215384,
  -82.9934094757403,
  -82.2746624960731,
  -83.2339201792762,
  -83.0754457880496,
  -83.2396167173873,
  -83.9323444601018,
  -83.2980453599921,
  -83.2051078391608,
  -82.9072280417929,
  -82.6120908756718,
  -83.569211356805,
  -83.7952017309971,
  -83.2089160937074,
  -83.4249723766544,
  -83.4224571728424,
  -83.253558610697,
  -83.92725626723,
  1,
  0,
  -83.8818640599643,
  0.438150044293079,
  -83.2378870975253,
  -83.4229397244709,
  -84.7738222436006,
  -83.6736060809219,
  -83.2784207902352,
  -83.7475789802126,
  -84.0360663699116,
  -84.1681495169304,
  -84.3801648188904,
  -84.1224507138305,
  -83.7342736916872,
  -84.2823016842682,
  -83.1722021388454,
  -83.2439702681155,
  -84.2998437737439,
  -83.9154154506125,
  -84.0113117572543,
  -84.0394076394494,
  -83.9405837034435,
  -84.1568847553379,
  1,
  0,
  -85.3151912511418,
  0.454398065106879,
  -84.9945403858473,
  -84.840392655847,
  -85.9125696034824,
  -85.1664832960841,
  -85.0049523282758,
  -84.860630782834,
  -85.2010082602832,
  -86.1794766579287,
  -85.4202366134526,
  -85.5250425219364,
  -84.6826785872501,
  -86.1861186265871,
  -84.8337419658179,
  -84.7239942749267,
  -85.7791126995117,
  -85.3646964083043,
  -85.2705356966893,
  -85.2422552729997,
  -85.6454111430632,
  -85.4699472417154,
  1,
  0,
  -86.9204292708872,
  0.405891756433377,
  -86.8433268152784,
  -86.0204623050971,
  -87.3114675289413,
  -86.6977142148949,
  -86.5146068625873,
  -86.9741412326673,
  -87.2419826391873,
  -87.4566602516288,
  -87.203288161241,
  -87.5354788388899,
  -86.2342969790927,
  -87.1673813555805,
  -86.8502520976113,
  -86.8167270691037,
  -86.5314710767427,
  -87.254582155942,
  -86.577369794157,
  -86.8746365353163,
  -87.3219006649616,
  -86.9808388388236,
  1,
  0,
  -88.523758803711,
  0.344675885721162,
  -88.1526089219836,
  -87.5291907138775,
  -88.5603031525875,
  -88.2351576604904,
  -88.4429164544456,
  -88.8839375894497,
  -88.5088801983509,
  -88.7283198261123,
  -88.654626829439,
  -88.9017704257145,
  -88.1241471838679,
  -88.6127814895192,
  -88.4654502262134,
  -88.6596709647964,
  -88.2454442699935,
  -88.9040810052632,
  -88.5664765062815,
  -88.5659993325686,
  -89.0353894932679,
  -88.6980238299989,
  1,
  0,
  -90.097411713196,
  0.392459042028477,
  -90.3114837993205,
  -89.4783549763737,
  -90.5266677924685,
  -90.183889531227,
  -90.0983148307998,
  -90.5063315582677,
  -90.5108544702964,
  -90.1970836493891,
  -90.321222105767,
  -90.791561975677,
  -89.7465599815655,
  -89.7493342704767,
  -89.7681435267992,
  -89.651870792608,
  -89.2450565785927,
  -90.1353117004213,
  -90.1755448597815,
  -90.1984493084536,
  -89.9333878990876,
  -90.4188106565468,
  1,
  0,
  -92.4524969909906,
  0.355262065317156,
  -92.8163013723775,
  -92.2497054731438,
  -92.45325290092,
  -92.448482025102,
  -92.1990242700173,
  -92.2218097035043,
  -92.8653491268725,
  -92.8563356391066,
  -92.6269230129861,
  -93.050527614721,
  -92.3238331182093,
  -92.1020818722258,
  -91.7804769626958,
  -93.0507514508844,
  -92.0717094514665,
  -92.2487900840821,
  -92.361940826816,
  -92.7338572559172,
  -92.0569734824354,
  -92.5318141763288,
  1,
  0,
  -94.3523473227332,
  0.335829242127448,
  -94.4215791226735,
  -94.2950239441135,
  -94.8548785569373,
  -94.6368380912245,
  -94.082605227543,
  -94.1778458768419,
  -94.4126522396419,
  -94.3139552857594,
  -94.7194999918933,
  -94.8503602573334,
  -94.4181846264348,
  -94.0196732373314,
  -93.6935149848331,
  -94.8514008743898,
  -93.8404664722036,
  -94.2596068566935,
  -94.4023686313176,
  -94.560545754139,
  -94.3249725566582,
  -93.9109738667009,
  1,
  0,
  -96.1190933853008,
  0.324265004046224,
  -96.4048506848058,
  -96.0308125046334,
  -96.4324944592273,
  -96.0513874050748,
  -96.1521643393394,
  -95.5667407699311,
  -95.954100882826,
  -95.7435010122343,
  -96.1525376150656,
  -96.7775657741018,
  -96.270680754277,
  -96.1273712902536,
  -95.5438053863514,
  -96.5574624561594,
  -96.3317750640539,
  -96.2388943547155,
  -96.0382453021073,
  -96.3379842700789,
  -96.0276933913182,
  -95.6417999894614,
  1,
  0,
  -97.4322166048734,
  0.329599666618754,
  -96.6828539838396,
  -97.0840794075614,
  -97.323137191532,
  -97.3701805551982,
  -97.5251796967722,
  -97.1588700599588,
  -97.2159666284421,
  -96.9828997809089,
  -97.688576544258,
  -97.8970605072657,
  -97.4991378257927,
  -97.4638849056849,
  -97.4142230425775,
  -98.0225996108896,
  -97.5882540451034,
  -97.2614766881099,
  -97.8544536346649,
  -97.5606812547094,
  -97.7820872969712,
  -97.2687294372276,
  1,
  0,
  -97.1894203950696,
  0.340902641919001,
  -96.5957243512481,
  -97.2229897795426,
  -96.9641482172729,
  -97.2957605841427,
  -97.4603665591966,
  -97.3164632710581,
  -96.983918372068,
  -96.6291133208293,
  -97.1591768701203,
  -97.2632502392911,
  -96.7227108411434,
  -97.0467849060054,
  -97.7739513127516,
  -97.3189379405701,
  -97.3849319762864,
  -97.3133654702917,
  -97.9103485092124,
  -97.0020202656376,
  -97.4712886937347,
  -96.9531564209896,
  1,
  0,
  -97.0169171502849,
  0.321918919451295,
  -97.4286245251382,
  -97.3460733269769,
  -97.0964656118491,
  -96.8190785973073,
  -97.2240108638783,
  -97.4260871751469,
  -96.7841827467175,
  -96.7337630065449,
  -96.7557543972456,
  -96.8237257660992,
  -96.5860728574509,
  -97.3375484966013,
  -97.2757803763348,
  -96.968165424309,
  -97.0360831959101,
  -96.5878357391787,
  -97.6231165066004,
  -96.6775989882493,
  -97.1736168651885,
  -96.6347585389712,
  1,
  0,
  -96.6373389009419,
  0.301274614790868,
  -96.6378146393876,
  -96.8284055633152,
  -96.8445760770961,
  -96.5437701172246,
  -96.8345905965989,
  -96.8227188779158,
  -97.0119344295782,
  -96.4900420879756,
  -96.8645466121046,
  -96.8201983962868,
  -96.3612951555799,
  -96.8164094387777,
  -95.9043138097768,
  -96.3901224718468,
  -96.7458664197375,
  -96.1322958108625,
  -96.9175375423351,
  -96.1820602889863,
  -96.8454834921562,
  -96.7527961912957,
  1,
  0,
  -95.8866782628249,
  0.296215931833846,
  -96.0224462840065,
  -95.9633715633911,
  -95.8127804447678,
  -96.1731967284824,
  -95.5840585623202,
  -95.948400260173,
  -96.3229678990792,
  -95.7692069977877,
  -95.5516980499004,
  -95.9746215506394,
  -95.5264585084258,
  -96.1961879130209,
  -95.714307428963,
  -96.0493257295594,
  -96.3881218333814,
  -95.4563026027589,
  -96.3227751927441,
  -95.8362402230896,
  -95.4832563269551,
  -95.6378411570513,
  1,
  0,
  -94.9618804207444,
  0.291944192390313,
  -94.6360183348702,
  -94.7763531084202,
  -94.7506719924283,
  -95.0789811293296,
  -94.7953800509502,
  -95.1970480847904,
  -95.029856492829,
  -94.5868426681928,
  -94.5381843956076,
  -95.4760281532839,
  -95.2074796403099,
  -95.0104945936371,
  -94.9105804640306,
  -95.4488019429681,
  -95.3174489233831,
  -94.5377053416433,
  -94.8738857641054,
  -95.2140785922219,
  -94.7447713594159,
  -95.1069973824706,
  1,
  0,
  -93.1641398696602,
  0.29739306832261,
  -93.0495966754165,
  -93.0471509096744,
  -92.9668307427688,
  -92.7492028046664,
  -93.4510445852723,
  -93.4545314240149,
  -93.2576814712063,
  -92.6342451969001,
  -92.9380631941406,
  -93.1383570365822,
  -92.9336815752405,
  -93.3215358015774,
  -93.0309309729435,
  -93.7438164888459,
  -93.5412705739625,
  -92.694519942357,
  -93.2879400101272,
  -93.2931699638948,
  -93.2757555520219,
  -93.4734724715913,
  1,
  0,
  -90.6971768780282,
  0.28316915297929,
  -90.7586442909236,
  -90.7808660917546,
  -90.6731112031227,
  -90.7394398846495,
  -90.7846206566457,
  -90.7415241394724,
  -90.2445946776057,
  -90.2456810395861,
  -90.6240723899108,
  -90.7815870593853,
  -90.3840681577275,
  -90.5146702426874,
  -90.7741075499302,
  -91.4299946711583,
  -90.946600818919,
  -90.3021195744981,
  -90.9445116513032,
  -90.5078726658568,
  -90.985598971684,
  -90.7798518237433,
  1,
  0,
  -89.1687031861055,
  0.287996192226422,
  -88.9463339617363,
  -89.227250305283,
  -89.2787707951445,
  -89.1567144079718,
  -89.2421028431825,
  -89.0912796235791,
  -88.8727975484309,
  -88.8578147547743,
  -89.1037366824014,
  -88.9772606148,
  -89.1398559869901,
  -88.7856810129925,
  -89.176482098187,
  -89.7778312148134,
  -89.7943509995025,
  -88.6766204632483,
  -89.3324510884249,
  -89.1714415176434,
  -89.425753977081,
  -89.3395338259237,
  1,
  0,
  -87.6622971625669,
  0.248269561456589,
  -87.5919183280103,
  -87.6877998179171,
  -87.777788582421,
  -87.7042787687109,
  -87.3738203427332,
  -87.6755131539647,
  -87.8524605925683,
  -87.1176131100515,
  -87.5914221519017,
  -87.7662668676559,
  -87.7443231789132,
  -87.5428569312218,
  -87.6754008844324,
  -88.2750188499769,
  -87.7951763764286,
  -87.3391576104746,
  -88.0414820805571,
  -87.5372429619704,
  -87.6924603527086,
  -87.4639423087203,
  1,
  0,
  -85.8788388663509,
  0.24383167039075,
  -85.7910208847417,
  -85.9649426890899,
  -85.968466019404,
  -86.0361461378875,
  -85.6560817256332,
  -85.8608176078901,
  -85.9304464689294,
  -85.4563037682217,
  -85.7293813137351,
  -85.8007365077907,
  -85.8706132521762,
  -85.9621299635389,
  -85.8847647719686,
  -86.5105249269405,
  -85.8999031332173,
  -86.0308583679117,
  -86.2006484734814,
  -85.3692952394901,
  -85.9361954089175,
  -85.7175006660537,
  1,
  0,
  -84.196108975426,
  0.268409768308546,
  -84.253005657178,
  -84.1857421534307,
  -84.4284353466992,
  -84.3175670563272,
  -83.9613827496638,
  -84.479709513224,
  -84.2483924321807,
  -83.9356031179245,
  -84.3023182877938,
  -83.9553840874735,
  -84.2097081656752,
  -84.1219584078443,
  -84.0533983592992,
  -84.9124410771809,
  -84.1354369547541,
  -83.9263649269,
  -84.4203290318448,
  -83.6217632864166,
  -84.1175897065972,
  -84.3356491901114,
  1,
  0,
  -83.6092792359255,
  0.268380888243813,
  -83.7647862314648,
  -83.5143738274388,
  -83.7892175925431,
  -83.7644927657742,
  -83.6296723722388,
  -83.6179911946648,
  -83.6787638522286,
  -83.3504382695001,
  -83.6577035269836,
  -83.7751565536585,
  -83.6730359592169,
  -83.336697116521,
  -83.4611578963328,
  -84.2745906624455,
  -83.3347903407194,
  -83.43178890738,
  -83.9675475836617,
  -83.0442902906815,
  -83.3666814383435,
  -83.7524083367132,
  1,
  0,
  -83.4564455766042,
  0.24912656562502,
  -83.4419946045906,
  -83.3367460988332,
  -83.8029837712756,
  -83.1973109292452,
  -83.5346178180314,
  -83.368942225861,
  -83.3506019114308,
  -83.5306150241072,
  -83.2253914729106,
  -83.4056607456793,
  -83.721250581725,
  -83.2066060543572,
  -83.4482382980419,
  -84.0460946303824,
  -83.4074669622608,
  -83.2523569360695,
  -83.9339572245053,
  -83.0920554458105,
  -83.4453142116004,
  -83.3807065853669,
  1,
  0,
  -83.6467692433561,
  0.216936925695796,
  -83.3788672433483,
  -83.7598037534093,
  -83.5491973501292,
  -83.7866776592792,
  -83.655189565509,
  -83.3924614444266,
  -83.3771776914633,
  -83.8167747476689,
  -83.4777054744489,
  -83.819364608521,
  -83.6848206947151,
  -83.9017288288647,
  -83.7265564686547,
  -83.8450524384678,
  -83.5638041090354,
  -83.404878456172,
  -83.9147878164058,
  -83.1970885180665,
  -83.722893930493,
  -83.9605540680436,
  1,
  0,
  -83.8844922841222,
  0.231234789382933,
  -83.7978362479765,
  -83.6664189772959,
  -83.726036902809,
  -83.8127939078411,
  -84.0263246996577,
  -83.9776078939512,
  -83.3408684459374,
  -84.096748495693,
  -83.9371029262369,
  -84.3256772319372,
  -84.0865059633155,
  -84.255003694772,
  -83.7222907874533,
  -83.9911688419221,
  -83.7581246699611,
  -84.0452011910239,
  -83.998166184074,
  -83.7042353284594,
  -83.7274322752532,
  -83.6943010168739,
  1,
  0,
  -84.97020088464,
  0.237531886424767,
  -84.9588051768405,
  -84.4438550568261,
  -84.5474198483333,
  -85.009165896773,
  -85.1675283906311,
  -85.2580160045711,
  -84.9858500330253,
  -85.2952171084039,
  -84.7063631599055,
  -85.1521080178083,
  -84.9279018523594,
  -85.3706521517422,
  -85.0971069353717,
  -84.8406091478518,
  -85.0797357725724,
  -84.8444707980729,
  -85.0954026088424,
  -84.943730211579,
  -84.9145463204266,
  -84.7655332008633,
  1,
  0,
  -86.8291188109372,
  0.244356500845551,
  -86.7803413059947,
  -86.6546227373313,
  -86.0518531497893,
  -86.7801155318195,
  -86.7760991680601,
  -86.8001090342747,
  -87.0978679305978,
  -86.9961319276701,
  -86.9488862638177,
  -86.7897829375874,
  -87.0066067733469,
  -87.0483130178221,
  -87.0380909567306,
  -86.8305176160579,
  -87.198500058452,
  -86.9576468834658,
  -86.8687991303837,
  -86.661583796421,
  -86.6941279078107,
  -86.6023800913106,
  1,
  0,
  -89.0627731000847,
  0.237061555562201,
  -88.853109290277,
  -88.9289248613694,
  -88.8526488492218,
  -88.993555981288,
  -88.5662052199051,
  -88.8799071987377,
  -89.2902283915673,
  -89.1217621001902,
  -89.417199723509,
  -89.1081452606575,
  -89.0557953663958,
  -89.360737638626,
  -89.140074469298,
  -88.8424327899314,
  -89.5216044696928,
  -89.223063097498,
  -89.0321026920347,
  -88.766344522965,
  -89.2220430889951,
  -89.079576989535,
  1,
  0,
  -91.2979928017293,
  0.234309309595772,
  -91.1554556171531,
  -91.2171611460445,
  -91.1065018775447,
  -91.2578696567178,
  -90.9503953523777,
  -91.3307258949204,
  -91.4715508614909,
  -91.0361306692641,
  -91.2909124938289,
  -91.1743752389519,
  -91.5833574222881,
  -91.8043669628828,
  -91.6054484381126,
  -91.2139980940252,
  -91.6053672540919,
  -90.967183430113,
  -91.2248855211042,
  -91.1663357312692,
  -91.2320782694792,
  -91.5657561029263,
  1,
  0,
  -93.8109909779091,
  0.227536751804149,
  -93.4234554345328,
  -93.7153449745764,
  -93.8997635107042,
  -93.7997810885931,
  -93.3017587168511,
  -93.9426026561852,
  -94.0112855620006,
  -93.5529362750827,
  -94.0002602543075,
  -93.9305709351027,
  -93.9137871870899,
  -94.2134949281267,
  -94.0129740995789,
  -93.8031619772324,
  -93.8548308013139,
  -93.7074053556294,
  -93.8505930834817,
  -93.9192241909046,
  -93.4478221023974,
  -93.9187664244902,
  1,
  0,
  -96.0687682468217,
  0.229094928585299,
  -96.0076665417397,
  -95.662340082032,
  -95.7479913144598,
  -96.2528312159364,
  -95.7536707821784,
  -96.3438330512428,
  -95.9508199184594,
  -96.1790729185446,
  -96.1111175836631,
  -95.9479784510923,
  -96.246372632476,
  -96.3349235387722,
  -96.2932917545161,
  -95.8166325579731,
  -95.9991831569747,
  -96.018444934426,
  -96.3128495793062,
  -96.2710149709404,
  -95.7889792987733,
  -96.3363506529283,
  1,
  0,
  -98.4799317692609,
  0.227086537334192,
  -98.6221518190254,
  -98.4638266059714,
  -98.6083106398133,
  -98.5233787442742,
  -98.851502237923,
  -98.5328226858039,
  -98.2592555548487,
  -97.9452970219946,
  -98.3510907969245,
  -98.2018158802167,
  -98.6861927284754,
  -98.6295906638737,
  -98.4039087215098,
  -98.2133994900328,
  -98.3913095183715,
  -98.7035190810345,
  -98.8403968958015,
  -98.5147948181299,
  -98.2948860926655,
  -98.5611853885286,
  1,
  0,
  -100.68996093524,
  0.220556951129674,
  -100.727544495107,
  -100.691302833283,
  -100.659996597331,
  -100.525360448566,
  -100.607767869672,
  -100.952762613231,
  -100.860838067182,
  -100.391177069927,
  -100.712778718145,
  -100.459063896031,
  -101.28267910713,
  -100.903114702929,
  -100.696683528624,
  -100.407067530245,
  -100.494770887232,
  -100.714168297829,
  -100.928076014555,
  -100.42823730063,
  -100.731461145266,
  -100.624367581889,
  1,
  0,
  -101.78424530943,
  0.200238251851125,
  -101.70246870199,
  -101.772778174473,
  -101.461755283862,
  -101.815775415885,
  -102.078098560989,
  -101.777186500182,
  -101.526352932221,
  -101.405307827158,
  -102.038740744356,
  -101.956524057028,
  -101.970129229099,
  -101.833785762233,
  -102.022524343585,
  -101.864309305241,
  -101.503406030114,
  -101.777234770106,
  -101.678209656096,
  -101.64002471954,
  -101.981710148356,
  -101.878584026089,
  1,
  0,
  -102.831037884016,
  0.209495621810426,
  -102.978441840436,
  -102.50827862218,
  -103.022779113647,
  -103.134576452812,
  -102.917241260357,
  -102.630227259543,
  -102.539196699984,
  -102.925355558164,
  -103.209470657209,
  -102.816038342233,
  -102.734805274903,
  -102.809630353907,
  -102.988428043776,
  -102.904539076647,
  -102.570219715162,
  -102.930167360537,
  -102.563913083019,
  -102.580925818125,
  -103.036095322837,
  -102.820427824838,
  1,
  0,
  -103.009785225607,
  0.199913952297935,
  -102.646659961013,
  -103.072574211588,
  -102.849790192732,
  -103.410528104806,
  -103.107989223823,
  -102.72934422935,
  -103.173040582781,
  -103.079799633609,
  -103.33046312907,
  -102.95446071064,
  -103.145458954451,
  -102.699467084463,
  -102.829405351516,
  -102.887944027102,
  -103.085226453669,
  -103.055452348871,
  -103.099538396336,
  -102.866393346346,
  -103.058824747498,
  -103.113343822473,
  1,
  0,
  -102.485412069723,
  0.201329331862665,
  -102.142764747995,
  -102.61839278656,
  -102.854096212234,
  -102.816925907448,
  -102.343559609954,
  -102.405992940518,
  -102.400011556072,
  -102.568259072667,
  -102.815024042058,
  -102.448803815059,
  -102.56542314586,
  -102.237298535042,
  -102.413183398876,
  -102.256639238596,
  -102.627254778376,
  -102.620189088363,
  -102.291272341376,
  -102.440741190265,
  -102.305199804917,
  -102.53720918222,
  1,
  0,
  -101.437842497425,
  0.192575694770429,
  -101.426874957461,
  -101.672971216973,
  -101.715466914892,
  -101.348388278114,
  -101.551660008996,
  -101.677756610241,
  -101.308936414434,
  -101.27486605411,
  -101.520697469415,
  -101.042482536984,
  -101.399627360529,
  -101.051174736862,
  -101.270535650353,
  -101.318601366821,
  -101.636853928951,
  -101.642506492857,
  -101.507369709037,
  -101.522000469705,
  -101.415972812292,
  -101.452106959473,
  1,
  0,
  -100.5978481555,
  0.202065790420492,
  -100.628669127414,
  -100.74680714174,
  -100.552308227895,
  -100.576145171736,
  -100.520838707721,
  -100.944014171134,
  -100.752134615348,
  -100.609204289009,
  -100.514161647923,
  -100.065085883032,
  -100.711320536909,
  -100.496699404435,
  -100.550157502418,
  -100.643270000483,
  -100.782970828662,
  -100.240585900877,
  -100.490228297645,
  -100.720366414667,
  -100.518611553426,
  -100.893383687518,
  1,
  0,
  -99.5791694423702,
  0.193937801723771,
  -99.3869666386721,
  -99.4558336330423,
  -99.2119827006966,
  -99.5236814509195,
  -99.6272513534104,
  -99.888503565056,
  -99.295037922037,
  -99.7251372470048,
  -99.543466071728,
  -99.4753834106953,
  -99.4945770244807,
  -99.5180468967669,
  -99.7912382632238,
  -99.6633766177942,
  -99.6624777194248,
  -99.5409877028536,
  -99.6892801109576,
  -99.4572964884642,
  -99.5910818398017,
  -100.041782190374,
  1,
  0,
  -97.9408450407093,
  0.195918857138366,
  -97.6656382916394,
  -97.9234601946299,
  -97.676976636545,
  -98.2070061565105,
  -98.0065623086287,
  -97.8836251788643,
  -97.8223013507335,
  -98.2554340098505,
  -97.8583182999307,
  -98.0353403913564,
  -97.9801427919165,
  -98.100647752356,
  -97.9933258447922,
  -98.0790723745986,
  -97.5234765413662,
  -97.7705613509671,
  -98.1966579525811,
  -97.8144043235094,
  -98.1399534743436,
  -97.8839955890655,
  1,
  0,
  -96.8260180836903,
  0.185405658672094,
  -96.7439566663654,
  -97.046656873154,
  -96.8263660230512,
  -96.6150909022476,
  -96.9828864897787,
  -96.5859279505601,
  -97.0406779793945,
  -96.735180854591,
  -96.8235414274241,
  -97.1184585447063,
  -96.9572089735326,
  -96.7414906794756,
  -96.6658822507158,
  -96.5398651705401,
  -96.7215058208607,
  -96.9368444145681,
  -96.9117245794102,
  -96.5413283698525,
  -96.8665019724659,
  -97.1192657311118,
  1,
  0,
  -96.1107855491031,
  0.173099097544714,
  -95.8366699683876,
  -96.2193805734034,
  -95.9344023120621,
  -96.1273530204404,
  -96.4976744745129,
  -96.0938292181918,
  -96.1053827604348,
  -95.7634579731056,
  -96.2652379163813,
  -96.1744719573174,
  -96.0771164973087,
  -95.9932567786039,
  -96.2302628559833,
  -96.0384449412611,
  -96.0010962944346,
  -96.2873306848573,
  -96.3696105507905,
  -96.1034183279518,
  -96.0516652063918,
  -96.0456486702422,
  1,
  0,
  -95.928371942138,
  0.189114285919834,
  -95.6850190094509,
  -96.2819271042471,
  -95.7164114824714,
  -95.8358411248943,
  -96.1246226889172,
  -95.9550121882427,
  -96.2142632965487,
  -95.8892766569905,
  -95.6409032025679,
  -95.9563447778368,
  -95.7499438627955,
  -95.7451934269829,
  -95.8273613530956,
  -95.7911887335577,
  -95.9943181304697,
  -95.9819928117595,
  -96.0084917839141,
  -95.9607010512485,
  -95.9241888264543,
  -96.2844373303154,
  1,
  0,
  -96.0944343493361,
  0.184355705513357,
  -96.0539311815023,
  -96.2706439026973,
  -95.9083317349131,
  -95.7932624626523,
  -95.937551817299,
  -95.9647602930507,
  -96.3751666744306,
  -95.7676864244858,
  -96.0652709695692,
  -96.1887134453721,
  -95.9879786556488,
  -95.9668163878771,
  -95.9314300497323,
  -96.2955570426325,
  -96.2459166792021,
  -96.2810752747411,
  -96.1296971126728,
  -96.1914879409453,
  -96.3861712640146,
  -96.1472376732829,
  1,
  0,
  -96.8864917724335,
  0.182529067919128,
  -96.8736959285165,
  -96.8569780461966,
  -96.9514883648993,
  -97.0907458976168,
  -96.8521995402554,
  -96.6051904425668,
  -97.2670285264902,
  -96.7416210791072,
  -96.7896985034233,
  -96.9223052668186,
  -96.6530575749518,
  -96.7055779771726,
  -96.688631092369,
  -96.8562491523227,
  -97.0122647794704,
  -97.0713810080199,
  -96.752375126012,
  -97.2424323832055,
  -96.9577556170853,
  -96.8391591421698,
  1,
  0,
  -98.2936564674569,
  0.186492474074395,
  -98.4692399471261,
  -98.1812210569527,
  -98.3632920308674,
  -98.2502656538626,
  -98.2778929692819,
  -98.1750379229312,
  -98.8012804519458,
  -98.3439406060715,
  -98.221264247178,
  -98.075417780256,
  -97.992325973462,
  -98.1676046390162,
  -98.2683243609729,
  -98.512815385182,
  -98.171447027365,
  -98.6038860131004,
  -98.2708209345254,
  -98.2730771485636,
  -98.1685298785824,
  -98.285445321895,
  1,
  0,
  -100.873400723019,
  0.182438961506971,
  -101.112019983635,
  -100.652575462089,
  -100.959331378496,
  -100.722854332491,
  -100.990906474801,
  -100.711875608144,
  -101.148731087608,
  -100.860046144066,
  -100.995896620033,
  -100.85312867698,
  -100.858885500964,
  -100.978486916009,
  -100.888973799652,
  -100.848843450714,
  -100.849963265459,
  -101.107345704283,
  -100.751276997594,
  -100.558817080981,
  -100.512547601067,
  -101.105508375313,
  1,
  0,
  -103.709816685835,
  0.17971445523767,
  -103.916593040598,
  -103.636273948803,
  -103.460978004895,
  -103.942098679313,
  -103.672259480385,
  -103.473809246588,
  -103.837852298597,
  -103.838621051267,
  -104.032792835764,
  -103.571883906487,
  -103.656025780122,
  -103.696482038202,
  -103.665089277292,
  -103.853428599026,
  -103.637282153601,
  -103.761223311946,
  -103.940725673587,
  -103.492587448404,
  -103.390493803226,
  -103.719833138603,
  1,
  0,
  -106.143305749834,
  0.1742167482904,
  -106.069908773984,
  -106.116718486233,
  -105.901745610271,
  -106.318294353641,
  -106.08141564778,
  -106.498395992007,
  -106.232338946081,
  -106.085526070795,
  -106.231073141664,
  -105.854319780279,
  -106.331502790552,
  -106.385374253168,
  -105.899934355597,
  -106.222530466107,
  -106.270555978497,
  -106.182100844221,
  -106.087886291622,
  -105.887061398607,
  -106.092865676667,
  -106.116566138913,
  1,
  0,
  -108.296461516184,
  0.171916207223368,
  -108.353423513106,
  -108.29029522405,
  -108.188796788555,
  -108.405017316026,
  -108.205347643756,
  -108.426935963393,
  -108.148309730678,
  -108.351211364852,
  -108.306425385322,
  -108.073708836364,
  -108.448831385277,
  -108.751478658784,
  -107.992007052961,
  -108.34361989522,
  -108.377603711034,
  -108.353637875496,
  -108.111168327658,
  -108.064953239207,
  -108.339574256745,
  -108.396884155187,
  1,
  0,
  -110.365312291917,
  0.167306439158501,
  -110.483867209713,
  -110.660291517032,
  -110.232437402238,
  -110.340648470076,
  -110.385837638674,
  -110.134152973341,
  -110.271787987782,
  -110.173650757913,
  -110.365466600558,
  -110.24908319274,
  -110.240723620717,
  -110.657014921366,
  -110.402191693827,
  -110.087524494762,
  -110.414972932475,
  -110.388887529353,
  -110.439085377193,
  -110.504397423828,
  -110.640090954768,
  -110.234133139975,
  1,
  0,
  -112.537936918867,
  0.168375653829276,
  -112.686276778788,
  -112.675749040584,
  -112.448776585704,
  -112.442534329816,
  -112.586100075659,
  -112.500235163147,
  -112.455672632107,
  -112.341824273224,
  -112.666871012419,
  -112.479106423978,
  -112.097308238032,
  -112.412743833002,
  -112.796463938113,
  -112.364406740857,
  -112.56971080697,
  -112.744477178578,
  -112.73085600113,
  -112.665573709495,
  -112.486048204502,
  -112.608003411228,
  1,
  0,
  -114.492473535697,
  0.168777654323576,
  -114.59090246713,
  -114.401573575666,
  -114.470845441419,
  -114.504354207257,
  -114.756228862331,
  -114.427332717462,
  -114.286739115554,
  -114.342451971161,
  -114.457541163074,
  -114.503700973973,
  -114.328876495489,
  -114.590707317263,
  -114.774409542694,
  -114.341746353627,
  -114.587114818844,
  -114.512775694992,
  -114.103764933625,
  -114.488867203939,
  -114.636222376114,
  -114.743315482325,
  1,
  0,
  -115.753125729916,
  0.166466608633098,
  -115.987257766635,
  -115.802358992459,
  -115.974861429526,
  -115.740997427958,
  -116.04964962759,
  -115.710251147287,
  -115.548901628458,
  -115.63090569604,
  -115.63701477971,
  -115.701082641599,
  -115.577223449623,
  -115.670914446934,
  -115.726479997599,
  -115.628287389628,
  -115.952143639833,
  -116.051500682865,
  -115.501024466449,
  -115.755962697488,
  -115.648426034014,
  -115.767270656622,
  1,
  0,
  -116.620024057778,
  0.157288922075805,
  -116.955931785558,
  -116.670440779927,
  -116.676627408646,
  -116.73991502193,
  -116.52852024244,
  -116.451769341413,
  -116.614526271951,
  -116.794715384048,
  -116.434212323248,
  -116.393940872692,
  -116.738142068661,
  -116.700243855208,
  -116.544200417807,
  -116.556871103869,
  -116.572036941104,
  -116.573954031663,
  -116.344552646359,
  -116.63414532034,
  -116.889236790559,
  -116.586498548134,
  1,
  0,
  -117.210258304486,
  0.160399253040755,
  -117.417249274055,
  -117.207011535442,
  -117.459479764322,
  -117.312011748858,
  -117.060539523156,
  -117.116651176116,
  -117.293317113114,
  -117.048028948866,
  -117.191470722887,
  -117.184287930922,
  -117.314196104054,
  -116.932330774479,
  -117.333558949611,
  -117.304070702244,
  -117.501713407833,
  -117.114454601701,
  -117.197696080741,
  -117.230615671149,
  -117.053018814979,
  -116.933463245195,
  1,
  0,
  -117.327513104029,
  0.156424057370802,
  -117.658634663119,
  -117.445679361519,
  -117.256810056381,
  -117.043103744832,
  -117.294784720299,
  -117.314632847154,
  -117.215955481961,
  -117.248672972159,
  -117.256509897078,
  -117.279313202837,
  -117.412468219255,
  -117.107605975239,
  -117.442629428351,
  -117.255724753637,
  -117.27768793926,
  -117.3262386754,
  -117.342636400152,
  -117.371869576715,
  -117.71204367773,
  -117.287260487505,
  1,
  0,
  -117.233279834446,
  0.15206681498394,
  -117.377657933239,
  -117.496298303096,
  -117.183625686854,
  -117.384427216917,
  -117.499441905306,
  -117.309324299182,
  -117.099466558828,
  -117.105795963938,
  -117.213584197691,
  -117.289436512466,
  -117.172474111974,
  -117.140163645152,
  -117.162226104835,
  -117.237441860434,
  -117.022456143703,
  -116.959870088652,
  -117.299613635981,
  -117.163765768518,
  -117.100370521163,
  -117.448156230994,
  1,
  0,
  -116.31109720274,
  0.151438088212701,
  -116.450164286734,
  -116.463085610806,
  -116.305709248301,
  -116.399906492091,
  -116.153635099806,
  -116.519215112221,
  -115.958023636966,
  -116.318136883844,
  -116.154414195193,
  -116.335318064733,
  -116.346933538295,
  -116.290635764793,
  -116.39842625863,
  -116.522433238643,
  -116.03017815485,
  -116.302526199184,
  -116.225529122313,
  -116.421005107871,
  -116.226635600237,
  -116.400032439292,
  1,
  0,
  -115.334792073625,
  0.149121805439478,
  -115.23580706102,
  -115.53424842127,
  -115.239850837248,
  -115.372797658472,
  -115.412973740555,
  -115.417083606967,
  -115.206704997734,
  -115.670707704142,
  -115.432507151259,
  -115.151018671633,
  -115.258702544904,
  -115.265358351264,
  -115.2445930412,
  -115.230677555945,
  -115.157232467232,
  -115.312313041536,
  -115.158096917861,
  -115.580132174353,
  -115.489398661612,
  -115.325636866291,
  1,
  0,
  -114.145805295618,
  0.146663522028958,
  -114.015323310953,
  -114.002249049927,
  -114.055714050817,
  -114.312821221594,
  -114.013259537524,
  -114.160442172569,
  -114.345905406257,
  -114.234732384307,
  -114.35451797679,
  -114.046126100036,
  -114.315008986187,
  -114.310565304178,
  -114.11551026851,
  -114.20707773724,
  -114.054478401573,
  -113.868547492652,
  -114.174328879077,
  -114.317412364614,
  -113.985657084838,
  -114.02642818272,
  1,
  0,
  -113.208476421283,
  0.146256000986171,
  -113.310396122001,
  -113.05997574463,
  -113.107675905263,
  -113.246731046399,
  -113.106768605296,
  -113.25476374566,
  -113.147151051001,
  -112.953563950664,
  -113.351788531062,
  -112.972753010877,
  -113.426134834966,
  -113.197236657634,
  -113.113642667947,
  -113.120207062452,
  -113.323065527521,
  -113.421915908877,
  -113.484265210857,
  -113.219344410998,
  -113.132609525997,
  -113.219538905552,
  1,
  0,
  -112.815573754344,
  0.140599022770319,
  -112.930345631951,
  -112.981987337209,
  -112.688385695069,
  -112.93187986387,
  -112.79440665416,
  -112.790826512421,
  -112.645689769375,
  -112.672462340792,
  -112.817530152668,
  -112.764673543202,
  -113.01082830151,
  -112.556023504127,
  -112.762667558364,
  -112.94578882244,
  -112.750787643755,
  -112.982359441467,
  -112.615515345274,
  -113.041936650862,
  -112.771880858393,
  -112.855499459964,
  1,
  0,
  -112.812201233,
  0.141358628497562,
  -112.92401952672,
  -112.936413479982,
  -112.802621739071,
  -112.738397262505,
  -112.819769916966,
  -112.827823723133,
  -112.439595690536,
  -112.698225872562,
  -112.618180198605,
  -112.834938250769,
  -112.87297284366,
  -112.886047837785,
  -112.699789418181,
  -112.92439547692,
  -112.972951769383,
  -112.790861100729,
  -112.838007883346,
  -112.944708858057,
  -112.642513164678,
  -113.03179064641,
  1,
  0,
  -113.239582381771,
  0.139712604258642,
  -113.359845291168,
  -113.331968754697,
  -113.416185295652,
  -113.073649965643,
  -113.247018339255,
  -113.369482769838,
  -113.095896951206,
  -113.003376174884,
  -113.108751940405,
  -113.364591888132,
  -113.241405361832,
  -113.231885847732,
  -113.405738191079,
  -113.015743745546,
  -113.14016698224,
  -113.316199767647,
  -113.164801905873,
  -113.316930441257,
  -113.132737405877,
  -113.455270615452,
  1,
  0,
  -114.254496033416,
  0.138249647210013,
  -114.25642408335,
  -114.18574605927,
  -114.186198540885,
  -114.195005088441,
  -113.968543891544,
  -114.45858980082,
  -114.16926842467,
  -114.40607793949,
  -114.091317290158,
  -114.428754850343,
  -114.241810320123,
  -114.177446668747,
  -114.255058217007,
  -114.292923291105,
  -114.377924045909,
  -114.284993366662,
  -114.025265458618,
  -114.233262656072,
  -114.46540664028,
  -114.389904034829,
  1,
  0,
  -115.640889463305,
  0.135602367814316,
  -115.879883341223,
  -115.771150464535,
  -115.499123591424,
  -115.450486293578,
  -115.734163208173,
  -115.711539539201,
  -115.518610397973,
  -115.582693039793,
  -115.679644025354,
  -115.47248596943,
  -115.587316034772,
  -115.474881306465,
  -115.749602493127,
  -115.627423185626,
  -115.447585734862,
  -115.619377156145,
  -115.784611576509,
  -115.740348592891,
  -115.85569758332,
  -115.631165731705,
  1,
  0,
  -117.430700841611,
  0.135077475226752,
  -117.680109571471,
  -117.428826927364,
  -117.323942244745,
  -117.341020791624,
  -117.517010928366,
  -117.463180123809,
  -117.2606218211,
  -117.58999511522,
  -117.422171582282,
  -117.412284503029,
  -117.242804280999,
  -117.559730535019,
  -117.480161037882,
  -117.441499481166,
  -117.365809694293,
  -117.525397570768,
  -117.44687439438,
  -117.162797218067,
  -117.304342738558,
  -117.645436272087,
  1,
  0,
  -119.71586642095,
  0.131386097893287,
  -119.653349084701,
  -119.696963430409,
  -119.779716870039,
  -119.835000160316,
  -119.435588085473,
  -119.773235747954,
  -119.681731289687,
  -119.854075945716,
  -119.626707571421,
  -119.608391908288,
  -119.667713112084,
  -119.663942194519,
  -119.805882204926,
  -119.779313551343,
  -119.77253078456,
  -119.735353542929,
  -119.700662855746,
  -119.552977222123,
  -119.621382549825,
  -120.072810306932,
  1,
  0,
  -121.774890358041,
  0.131623235157372,
  -121.727167811276,
  -121.706778600485,
  -121.571373969745,
  -121.677668526061,
  -121.856399018207,
  -121.895203154202,
  -121.740662851097,
  -121.84716711187,
  -121.518512106136,
  -121.623377277439,
  -121.683041553864,
  -121.943060385371,
  -121.7808366531,
  -121.979841527891,
  -121.848960929907,
  -121.922539733304,
  -121.767563480803,
  -121.843492613071,
  -121.633296425159,
  -121.930863431841,
  1,
  0,
  -123.797627677646,
  0.129562010325352,
  -123.839207526181,
  -123.959761547755,
  -123.861104688705,
  -123.649496412488,
  -123.871291977336,
  -123.874234615832,
  -123.893573571737,
  -123.95835148389,
  -123.597025974415,
  -123.887695602856,
  -123.656635781414,
  -123.794925463954,
  -123.976106726194,
  -123.869209891308,
  -123.576963723877,
  -123.838578849749,
  -123.710435482353,
  -123.62716914185,
  -123.862174638171,
  -123.648610452863,
  1,
  0,
  -125.79132911035,
  0.12826987710339,
  -125.745282928634,
  -125.892562699141,
  -125.850140140798,
  -125.701562955844,
  -125.802991124052,
  -125.646035584042,
  -125.716744732875,
  -125.897710738125,
  -125.871932367346,
  -126.064671234893,
  -125.850720598282,
  -125.966517867251,
  -125.871004997796,
  -125.71950337977,
  -125.789919459472,
  -125.516419471731,
  -125.747680111296,
  -125.577894630687,
  -125.814714347742,
  -125.782572837218,
  1,
  0,
  -127.566356421656,
  0.127017364845391,
  -127.797907493013,
  -127.671426089585,
  -127.626962539304,
  -127.554522671291,
  -127.554716002146,
  -127.397252175815,
  -127.561605479097,
  -127.471876460733,
  -127.615008780671,
  -127.483663721424,
  -127.725065453726,
  -127.399668498554,
  -127.605215850956,
  -127.663653564317,
  -127.793978754548,
  -127.497703441709,
  -127.639243528745,
  -127.375504825664,
  -127.450169013615,
  -127.441984088218,
  1,
  0,
  -129.27743856,
  0.124040249614604,
  -129.305619261179,
  -129.199730326837,
  -129.424944912587,
  -129.497353355585,
  -129.171692326841,
  -129.188611690391,
  -129.182644460176,
  -129.245717440239,
  -129.312226855028,
  -129.215977142069,
  -129.397798522175,
  -129.019536603496,
  -129.115980334266,
  -129.343825983488,
  -129.465000615265,
  -129.360491017223,
  -129.349371459512,
  -129.288491004651,
  -129.327604813986,
  -129.136153075012,
  1,
  0,
  -129.850794753193,
  0.123065602716752,
  -129.815173441519,
  -129.673171253433,
  -129.963863045,
  -129.897211252456,
  -129.664007598739,
  -129.912301384035,
  -129.861452042858,
  -129.716410198733,
  -129.907434211492,
  -129.975833628347,
  -129.884018914507,
  -129.763865710349,
  -130.030799308568,
  -129.749191066742,
  -130.097097434821,
  -129.718460090386,
  -129.74688094879,
  -129.907825385467,
  -129.764779427415,
  -129.966118720205,
  1,
  0,
  -129.816455860793,
  0.122018126691159,
  -129.849304255382,
  -129.7248041846,
  -129.789913527123,
  -129.74331644204,
  -129.81612672677,
  -129.75607521076,
  -129.810986096101,
  -129.854471996928,
  -130.082668443925,
  -129.902342476587,
  -129.931120128685,
  -129.883060105633,
  -129.802282724957,
  -129.492814116051,
  -129.964422699076,
  -129.871435972974,
  -129.824641104383,
  -129.760448972417,
  -129.634746771721,
  -129.834135259748,
  1,
  0,
  -129.519763695754,
  0.119254412894993,
  -129.429738721715,
  -129.36783286255,
  -129.532364347069,
  -129.496366062168,
  -129.504815315675,
  -129.380848880297,
  -129.409560509205,
  -129.569803437186,
  -129.582709435434,
  -129.459901700133,
  -129.421990133629,
  -129.911298843715,
  -129.507071643698,
  -129.499734864103,
  -129.583582952022,
  -129.54503281462,
  -129.647880856151,
  -129.518796240636,
  -129.435636645345,
  -129.590307649733,
  1,
  0,
  -128.737357796315,
  0.11989201940735,
  -128.803127241237,
  -128.479072774425,
  -128.53716246088,
  -128.814428819479,
  -128.710940921899,
  -128.837639805841,
  -128.716231834312,
  -128.941794168219,
  -128.834206228589,
  -128.815677723677,
  -128.744944200663,
  -128.913930479002,
  -128.653900002213,
  -128.798124265895,
  -128.704927079559,
  -128.624035848882,
  -128.754841914126,
  -128.575197692916,
  -128.693083422025,
  -128.793889042454,
  1,
  0,
  -127.600156832383,
  0.117309304445995,
  -127.628762764729,
  -127.613276686435,
  -127.630525639132,
  -127.764938193937,
  -127.651878312975,
  -127.845937841648,
  -127.456314688741,
  -127.75717955459,
  -127.479156355155,
  -127.594875393774,
  -127.518910314906,
  -127.574674288943,
  -127.444685430555,
  -127.74703094877,
  -127.483727628088,
  -127.572647283116,
  -127.538742196886,
  -127.718898301974,
  -127.496443876776,
  -127.484530946542,
  1,
  0,
  -126.47671555415,
  0.11708703960286,
  -126.4288420428,
  -126.404450805288,
  -126.438406969894,
  -126.481445664017,
  -126.428621276505,
  -126.315074848614,
  -126.397170608916,
  -126.555961598599,
  -126.619008957272,
  -126.406752408953,
  -126.482080095475,
  -126.352323053391,
  -126.480548163682,
  -126.573940796901,
  -126.745943953829,
  -126.3129327353,
  -126.40286750649,
  -126.469018569445,
  -126.705310065704,
  -126.533610961928,
  1,
  0,
  -124.915450479066,
  0.115397487818306,
  -124.962013827643,
  -124.984575636508,
  -125.017149573249,
  -124.839388328753,
  -124.940476488024,
  -125.056176904759,
  -124.739974329965,
  -124.685916811319,
  -124.936516665866,
  -125.057234847222,
  -125.017728352885,
  -125.055953223549,
  -124.892123458448,
  -125.00447038308,
  -124.927916843635,
  -124.852342086901,
  -124.914562269609,
  -124.672614011575,
  -124.858840591764,
  -124.893034946569,
  1,
  0,
  -123.585048490081,
  0.114744556898546,
  -123.723617454858,
  -123.66470846113,
  -123.771431644951,
  -123.666209708275,
  -123.382619992978,
  -123.735137616895,
  -123.525785439094,
  -123.579842860598,
  -123.396143722582,
  -123.687949653944,
  -123.480447743976,
  -123.408873905095,
  -123.536544503187,
  -123.60330716523,
  -123.603304512655,
  -123.52921992025,
  -123.627822190642,
  -123.642963209148,
  -123.65712201521,
  -123.477918080924,
  1,
  0,
  -122.680751403305,
  0.113609443003947,
  -122.770382174651,
  -122.824073186363,
  -122.701426200803,
  -122.558268005311,
  -122.549877302079,
  -122.589704864459,
  -122.79624783684,
  -122.757565594361,
  -122.428799275471,
  -122.762059348876,
  -122.614190647286,
  -122.654270914701,
  -122.864602806621,
  -122.755391835872,
  -122.621992812878,
  -122.745461905861,
  -122.530283949755,
  -122.782112569813,
  -122.651997129675,
  -122.656319704419,
  1,
  0,
  -121.990602460068,
  0.114061763789315,
  -121.993099930485,
  -121.89178351446,
  -121.918597542557,
  -122.069930628698,
  -121.89531561789,
  -121.998737120158,
  -122.117169206463,
  -122.068639730115,
  -121.899257777259,
  -122.0561446883,
  -122.173115423555,
  -121.85794008107,
  -121.935886829554,
  -122.155965219573,
  -122.163420639817,
  -121.74772515074,
  -121.967406627458,
  -121.895237915453,
  -121.971818440672,
  -122.034857117089,
  1,
  0,
  -121.482514576214,
  0.112494442135766,
  -121.450063045165,
  -121.479741568575,
  -121.486544734362,
  -121.411713875624,
  -121.266360237916,
  -121.413680620091,
  -121.625206722817,
  -121.604531566394,
  -121.53639181756,
  -121.536118228378,
  -121.317535310344,
  -121.479518003354,
  -121.541775229214,
  -121.549734528683,
  -121.649037232236,
  -121.629583715207,
  -121.256133526986,
  -121.53377115587,
  -121.441743244169,
  -121.441107161336,
  1,
  0,
  -121.497988298516,
  0.112165562574285,
  -121.534595460269,
  -121.334490132717,
  -121.530363069613,
  -121.346920023399,
  -121.462318163903,
  -121.612749844844,
  -121.480446359988,
  -121.709308503497,
  -121.352290889501,
  -121.419354353186,
  -121.357501541182,
  -121.489087950391,
  -121.464144433116,
  -121.712534467529,
  -121.38850144388,
  -121.61645807362,
  -121.566186696579,
  -121.528138029102,
  -121.528442257098,
  -121.525934276906,
  1,
  0,
  -122.085311317559,
  0.112478556902754,
  -122.174536917196,
  -121.790188445563,
  -122.030283392383,
  -122.125323690102,
  -122.055836892363,
  -122.135154227305,
  -122.112103962673,
  -122.093869219058,
  -122.063537308771,
  -122.141531885054,
  -122.13421633819,
  -122.215256472628,
  -122.011480283235,
  -122.155639433649,
  -121.948048155119,
  -122.277543241402,
  -122.213523833994,
  -121.918065733521,
  -122.079535190534,
  -122.030551728433,
  1,
  0,
  -123.010355863338,
  0.111863081243618,
  -122.928358621406,
  -122.882281878683,
  -122.896987881127,
  -123.04491200639,
  -122.927166961905,
  -123.088584328449,
  -122.913417747286,
  -123.042196068754,
  -122.970007639077,
  -123.11786626585,
  -122.998633163101,
  -123.067211557355,
  -123.036850658665,
  -122.982969940292,
  -123.276157191564,
  -122.961425587702,
  -122.774049876075,
  -123.108666568092,
  -123.151024958292,
  -123.038348366697,
  1,
  0,
  -124.09955480294,
  0.110123328894475,
  -124.159312996584,
  -124.091046575733,
  -124.076734790989,
  -123.985775130939,
  -123.964707822181,
  -124.059540689047,
  -124.171049458628,
  -124.037611171811,
  -123.897094726872,
  -124.231780322384,
  -123.994186248166,
  -123.90805470769,
  -124.116159617124,
  -124.088783121284,
  -124.207665586152,
  -124.267435470812,
  -124.124270589923,
  -124.228287702105,
  -124.144831789694,
  -124.236767540691,
  1,
  0,
  -125.375466026254,
  0.110858088569851,
  -125.576332818786,
  -125.32027429978,
  -125.566750757647,
  -125.392826814298,
  -125.305932786006,
  -125.343668467841,
  -125.320256998557,
  -125.27558248392,
  -125.194449250571,
  -125.311851875693,
  -125.269904523459,
  -125.423662249245,
  -125.327510526339,
  -125.310044796049,
  -125.428035944953,
  -125.255001213056,
  -125.345907367259,
  -125.488175027766,
  -125.548538519864,
  -125.504613803986,
  1,
  0,
  -127.036355010938,
  0.109970303419101,
  -127.035880931601,
  -126.976586027712,
  -126.934408382377,
  -127.106878231735,
  -127.075231220682,
  -126.889723924861,
  -126.983861479607,
  -127.006999325591,
  -126.988690052759,
  -127.191707479024,
  -126.997154860981,
  -126.940051601881,
  -126.903134025777,
  -127.088149748458,
  -127.078827298747,
  -126.842267873093,
  -127.100465316629,
  -127.215118757419,
  -127.241851191089,
  -127.130112488731,
  1,
  0,
  -128.311120020032,
  0.11016823523549,
  -128.498820187212,
  -128.252539992025,
  -128.205190086388,
  -128.165289273259,
  -128.437075570848,
  -128.235112012244,
  -128.370303053512,
  -128.227939134098,
  -128.359250412837,
  -128.420325583865,
  -128.200929293988,
  -128.176114956789,
  -128.170197362131,
  -128.470677225606,
  -128.263342205281,
  -128.304791464588,
  -128.398233086357,
  -128.341922964605,
  -128.258762133509,
  -128.465584401499,
  1,
  0,
  -129.214403186641,
  0.109834010016199,
  -129.283077773845,
  -129.278632476138,
  -129.248468524502,
  -129.147182104149,
  -129.310857108594,
  -129.206035150101,
  -129.141377189591,
  -129.243132063964,
  -129.102399738661,
  -129.491972428147,
  -129.220600766428,
  -129.158303132229,
  -129.339342875782,
  -128.955319641695,
  -129.205591843317,
  -129.183139775266,
  -129.187266128584,
  -129.097278261495,
  -129.187570575497,
  -129.300516174835,
  1,
  0,
  -129.465657252361,
  0.109930917197491,
  -129.56021362632,
  -129.5094350695,
  -129.43112586847,
  -129.293254252541,
  -129.347629818156,
  -129.45171318755,
  -129.380315539006,
  -129.579439055796,
  -129.340479809385,
  -129.500649933351,
  -129.627611343195,
  -129.507073554732,
  -129.523243263643,
  -129.544716817147,
  -129.490152716754,
  -129.41744233803,
  -129.620804453979,
  -129.210886493912,
  -129.543860579977,
  -129.43309732577,
  1,
  0,
  -129.37123935153,
  0.10885368672056,
  -129.238136674859,
  -129.348933769058,
  -129.28577719782,
  -129.332146743723,
  -129.416053053212,
  -129.252158410112,
  -129.310110589211,
  -129.439907371027,
  -129.209413465892,
  -129.576683668621,
  -129.56092835843,
  -129.395102553163,
  -129.511470345802,
  -129.334025922816,
  -129.301276384937,
  -129.300292382202,
  -129.300417213127,
  -129.519805535306,
  -129.463902711537,
  -129.328244679744,
  1,
  0,
  -128.687426834448,
  0.108208332137921,
  -128.626898125092,
  -128.842132232519,
  -128.662777688472,
  -128.572988319531,
  -128.806316760955,
  -128.683630930169,
  -128.617034633607,
  -128.748359373991,
  -128.551275617183,
  -128.681038361175,
  -128.641280584908,
  -128.561082622981,
  -128.687798257148,
  -128.718701888604,
  -128.849359727908,
  -128.899969171486,
  -128.700075761946,
  -128.710286550147,
  -128.718426219531,
  -128.469103861617,
  1,
  0,
  -127.562596541183,
  0.109772578002375,
  -127.732550980207,
  -127.573473013004,
  -127.529262580014,
  -127.418976270496,
  -127.542542074842,
  -127.49859869127,
  -127.461855135393,
  -127.747463202101,
  -127.568172261033,
  -127.459112948437,
  -127.58267810885,
  -127.609826518419,
  -127.688948374298,
  -127.497158434549,
  -127.435726470221,
  -127.624705123724,
  -127.385282220949,
  -127.491021278426,
  -127.691758175376,
  -127.712818962049,
  1,
  0,
  -126.437445200564,
  0.108386077432882,
  -126.463806980469,
  -126.630116679699,
  -126.395065370992,
  -126.498507613553,
  -126.566616700969,
  -126.350585861912,
  -126.315110208605,
  -126.397796915018,
  -126.282613687567,
  -126.445494456099,
  -126.461224483999,
  -126.29829140399,
  -126.494610975319,
  -126.59762618247,
  -126.396833546469,
  -126.370005636994,
  -126.315117958825,
  -126.555663437751,
  -126.580006547169,
  -126.333809363417,
  1,
  0,
  -125.036231027223,
  0.108912221462493,
  -125.075393154829,
  -125.044518126392,
  -124.879890329263,
  -124.940355020211,
  -125.120469056323,
  -125.078230024528,
  -124.867741721458,
  -125.045782630241,
  -124.963131820679,
  -124.960064470598,
  -125.218011072106,
  -125.06982331924,
  -125.129131648171,
  -125.250037078568,
  -125.085171893181,
  -125.048120987911,
  -124.950159672099,
  -124.860772930781,
  -125.140573666927,
  -124.997241920951,
  1,
  0,
  -123.326325075874,
  0.109961116623221,
  -123.212505963053,
  -123.388606177214,
  -123.220778544843,
  -123.400653520104,
  -123.428080318414,
  -123.29609433361,
  -123.106974699487,
  -123.372431500548,
  -123.442975646899,
  -123.423516107737,
  -123.44308600009,
  -123.543017459154,
  -123.391531613921,
  -123.219412894837,
  -123.306091877526,
  -123.336211605,
  -123.159935494866,
  -123.271657526408,
  -123.271439931839,
  -123.291500301938,
  1,
  0,
  -121.587752049352,
  0.110205803017996,
  -121.634780866149,
  -121.747473961636,
  -121.532426092544,
  -121.674650759789,
  -121.530837646574,
  -121.496946591386,
  -121.598064036549,
  -121.514164850637,
  -121.670877616245,
  -121.656553396692,
  -121.546443805835,
  -121.520368452439,
  -121.67015285929,
  -121.541640938652,
  -121.273215287718,
  -121.772327520128,
  -121.554436993749,
  -121.605084411353,
  -121.6892647009,
  -121.525330198782,
  1,
  0,
  -119.982872444266,
  0.111401674164126,
  -120.107188730622,
  -119.94343098465,
  -119.919232334543,
  -120.088032212507,
  -120.030304739654,
  -119.983483378422,
  -119.985471751349,
  -119.962898482707,
  -119.885595145524,
  -120.052673359244,
  -119.854693149786,
  -119.819214150209,
  -120.030080152835,
  -120.014105690297,
  -119.733145686042,
  -120.126073187695,
  -120.137288705912,
  -120.103345955139,
  -119.852658956705,
  -120.028532131472,
  1,
  0,
  -118.565730067168,
  0.111209473052979,
  -118.671813722401,
  -118.682152793416,
  -118.581674278656,
  -118.459846808731,
  -118.640169577004,
  -118.575783106835,
  -118.568863550798,
  -118.730507143584,
  -118.644148009174,
  -118.385013822221,
  -118.582291649712,
  -118.438102843007,
  -118.484015062003,
  -118.572750668283,
  -118.789785514595,
  -118.505243661788,
  -118.609931018098,
  -118.521667322716,
  -118.357661060709,
  -118.513179729624,
  1,
  0,
  -117.582375422738,
  0.112146221833062,
  -117.595581186456,
  -117.618417540814,
  -117.593839540335,
  -117.442498596078,
  -117.574020005449,
  -117.70000009591,
  -117.615272212907,
  -117.434747486021,
  -117.713925302184,
  -117.72265219879,
  -117.57925976649,
  -117.627117290073,
  -117.389072483014,
  -117.421323410739,
  -117.732205779175,
  -117.625180683487,
  -117.58527152961,
  -117.504778836239,
  -117.741685317078,
  -117.430659193905,
  1,
  0,
  -116.970325019137,
  0.112779568289311,
  -116.979614551504,
  -117.088471226705,
  -117.144604991121,
  -116.874847804136,
  -117.091055761797,
  -117.048016370776,
  -117.004018954031,
  -116.795040105658,
  -117.065505402012,
  -116.992471204909,
  -116.941667928387,
  -116.853822885921,
  -116.892817304005,
  -117.069957509238,
  -117.023470953088,
  -116.829242435821,
  -116.980713109804,
  -116.79418719258,
  -117.113251671662,
  -116.823723019583,
  1,
  0,
  -116.566501014218,
  0.113033580880398,
  -116.651039065649,
  -116.504632480778,
  -116.440128187532,
  -116.420110421109,
  -116.711833728169,
  -116.546871139148,
  -116.43205375466,
  -116.402038773862,
  -116.708148365728,
  -116.726995701306,
  -116.557658379866,
  -116.625819782396,
  -116.491154528662,
  -116.581265124194,
  -116.573247689394,
  -116.499623187003,
  -116.602012289542,
  -116.771269568828,
  -116.43359014396,
  -116.650527972567,
  1,
  0,
  -116.40366114386,
  0.112867286936339,
  -116.391247011808,
  -116.250393157057,
  -116.514683030863,
  -116.447511894606,
  -116.499823076978,
  -116.587742595554,
  -116.442410175114,
  -116.463150919764,
  -116.395316475851,
  -116.379079703195,
  -116.530846612036,
  -116.263058191584,
  -116.443649191456,
  -116.35806198083,
  -116.494191468099,
  -116.404048863125,
  -116.321276819468,
  -116.486064250511,
  -116.125437280913,
  -116.275230178396,
  1,
  0,
  -116.49184742991,
  0.114596029342939,
  -116.446536139986,
  -116.629730967816,
  -116.308127848162,
  -116.476350978538,
  -116.328849248727,
  -116.598663638186,
  -116.527283116437,
  -116.603093431956,
  -116.516116585114,
  -116.477818101529,
  -116.662953223255,
  -116.353452048725,
  -116.457440166707,
  -116.478479361599,
  -116.473356212812,
  -116.552180213211,
  -116.36778854881,
  -116.721285903,
  -116.350356752835,
  -116.5070861108,
  1,
  0,
  -116.733928258506,
  0.116612967296125,
  -116.758091270307,
  -116.955277065312,
  -116.604701204074,
  -116.524246679917,
  -116.535128552502,
  -116.836168300507,
  -116.552875606261,
  -116.865435574238,
  -116.688062067534,
  -116.818063272139,
  -116.836851544051,
  -116.711509177998,
  -116.773863915913,
  -116.865522054969,
  -116.769731423543,
  -116.661389668934,
  -116.736037650135,
  -116.692515593214,
  -116.758951105043,
  -116.73414344354,
  1,
  0,
  -117.417638798094,
  0.114595807163695,
  -117.346349536886,
  -117.454486957168,
  -117.232195757268,
  -117.17223017835,
  -117.449073598228,
  -117.56629732455,
  -117.451421552514,
  -117.517818062159,
  -117.508601697013,
  -117.243570125396,
  -117.420071371381,
  -117.357241597717,
  -117.507129572215,
  -117.475283577384,
  -117.472754415418,
  -117.512542165185,
  -117.229511865214,
  -117.470238206915,
  -117.513733813896,
  -117.452224587016,
  1,
  0,
  -117.946389176125,
  0.116729800030019,
  -117.95181033307,
  -118.010642851823,
  -117.958181661233,
  -118.011758819212,
  -117.848627484821,
  -117.957197467828,
  -117.949706994463,
  -117.989644082262,
  -117.973535940479,
  -118.003044845643,
  -117.832689122524,
  -118.062953865846,
  -118.022688660393,
  -117.849330619052,
  -117.689975051706,
  -118.095103898176,
  -117.986793368956,
  -118.16523456333,
  -117.744365996716,
  -117.824497894961,
  1,
  0,
  -118.156094581169,
  0.117410337271347,
  -118.089762262859,
  -118.027909836477,
  -118.115142117401,
  -118.134423488431,
  -118.151913131673,
  -118.376087494233,
  -118.295752737168,
  -118.141228099419,
  -118.07937908421,
  -118.245166873383,
  -118.126428907934,
  -118.048482507553,
  -118.072874379502,
  -118.473224337704,
  -118.094524395026,
  -118.117891732148,
  -118.16706840829,
  -118.179637464301,
  -117.985235814745,
  -118.199758550922,
  1,
  0,
  -118.418347084454,
  0.119485831103467,
  -118.337182427608,
  -118.384499675294,
  -118.569314920023,
  -118.266749371277,
  -118.524832047044,
  -118.473869963454,
  -118.242073091587,
  -118.539715911169,
  -118.232431269607,
  -118.516405573226,
  -118.329390449467,
  -118.317829678422,
  -118.218958676487,
  -118.526618256057,
  -118.555837238945,
  -118.49712600478,
  -118.498135212284,
  -118.439325644315,
  -118.519529013898,
  -118.377117264144,
  1,
  0,
  -118.621529025432,
  0.121442008396594,
  -118.566107118106,
  -118.682180732597,
  -118.476593220725,
  -118.676368535248,
  -118.765978910305,
  -118.437903596367,
  -118.557642999456,
  -118.750740622609,
  -118.705201286988,
  -118.766034079493,
  -118.666425625393,
  -118.504213380144,
  -118.632586413627,
  -118.810997150618,
  -118.512167975048,
  -118.57536798288,
  -118.538003842273,
  -118.811430308784,
  -118.440653162723,
  -118.553983565246,
  1,
  0,
  -118.357409104694,
  0.121968274339996,
  -118.492981171003,
  -118.394856042233,
  -118.295009816089,
  -118.400588559805,
  -118.606473612449,
  -118.252014483294,
  -118.259888076188,
  -118.386132997962,
  -118.37679687722,
  -118.489168551604,
  -118.454978547822,
  -118.319011625487,
  -118.091502262557,
  -118.543338340429,
  -118.398055973985,
  -118.288028910736,
  -118.2762384829,
  -118.244692426259,
  -118.336985251581,
  -118.241440084284,
  1,
  0,
  -118.299100611063,
  0.1227618568219,
  -118.318229369913,
  -118.420400765244,
  -118.348291765543,
  -118.554629754175,
  -118.132499368399,
  -118.336255556747,
  -118.060550367242,
  -118.233844162987,
  -118.242509807151,
  -118.386194424738,
  -118.502390764688,
  -118.248440781462,
  -118.305757012069,
  -118.378299157307,
  -118.184054477675,
  -118.341116606695,
  -118.191763241856,
  -118.243651088596,
  -118.172564397158,
  -118.380569351624,
  1,
  0,
  -117.320547066733,
  0.125972853036038,
  -117.335618007104,
  -117.412659473269,
  -117.051207770227,
  -117.499259923999,
  -117.314563314257,
  -117.126569556747,
  -117.094617186145,
  -117.450688623761,
  -117.336867925438,
  -117.466941056923,
  -117.415739132379,
  -117.39343109192,
  -117.375508771117,
  -117.371137016613,
  -117.364599675752,
  -117.155155940138,
  -117.39380439657,
  -117.275488357451,
  -117.254746252177,
  -117.322337862663,
  1,
  0,
  -116.468434109565,
  0.127164463692187,
  -116.397627974011,
  -116.620127476614,
  -116.495390843266,
  -116.546018444993,
  -116.302234121582,
  -116.383700335612,
  -116.368102592179,
  -116.549062938126,
  -116.371522100925,
  -116.454948141752,
  -116.83063676704,
  -116.293569699518,
  -116.368497014352,
  -116.45459550709,
  -116.475681217223,
  -116.530925425449,
  -116.339836805083,
  -116.497640558551,
  -116.602291988676,
  -116.486272239262,
  1,
  0,
  -115.231186845938,
  0.124243490340841,
  -115.202688826585,
  -115.409201189114,
  -115.169874583217,
  -115.182875053584,
  -115.144518689211,
  -115.227247902998,
  -115.396734383033,
  -115.070789797088,
  -115.027570519504,
  -115.031200378854,
  -115.377337901263,
  -115.280579294342,
  -115.198082702053,
  -115.348730259362,
  -115.309765054698,
  -115.205596570965,
  -115.077751513714,
  -115.261672347047,
  -115.267168732469,
  -115.434351219657,
  1,
  0,
  -113.542378083378,
  0.129917769514696,
  -113.630582189572,
  -113.595525984522,
  -113.472271802675,
  -113.524847933085,
  -113.357144717707,
  -113.511242764053,
  -113.790016166,
  -113.463078094639,
  -113.352994343762,
  -113.379453063236,
  -113.512127632909,
  -113.506483162983,
  -113.418313709829,
  -113.573063025953,
  -113.784256088624,
  -113.73089958609,
  -113.628868169555,
  -113.454501999088,
  -113.514604362859,
  -113.647286870428,
  1,
  0,
  -112.073370665034,
  0.12895103690614,
  -112.129692439567,
  -112.272389360364,
  -112.317363438138,
  -112.122101670215,
  -112.063439352035,
  -112.031908621052,
  -112.252969269495,
  -112.004173301994,
  -111.970592715403,
  -112.037806326279,
  -111.968073991522,
  -112.028411006409,
  -111.863569691978,
  -112.169437835447,
  -112.017225325297,
  -112.196943390897,
  -111.977010991473,
  -112.089167589681,
  -112.132316667722,
  -111.822820315716,
  1,
  0,
  -110.589107196882,
  0.132016940349619,
  -110.528962278795,
  -110.730807746273,
  -110.306292433343,
  -110.632384093922,
  -110.570447517609,
  -110.625235421402,
  -110.579608203336,
  -110.777513240552,
  -110.542968064298,
  -110.5725635942,
  -110.498488618664,
  -110.616837996052,
  -110.672118005375,
  -110.81742265156,
  -110.599253226045,
  -110.439529482531,
  -110.415135189061,
  -110.418446020272,
  -110.685161296628,
  -110.752968857728,
  1,
  0,
  -109.241161917594,
  0.131768574913325,
  -109.155148601038,
  -109.334342225446,
  -109.219497460033,
  -109.341316617301,
  -109.190826997217,
  -109.161919037667,
  -109.10489129435,
  -109.480650870499,
  -109.286189110554,
  -109.403165684731,
  -109.089036990801,
  -109.301485725222,
  -109.336896719712,
  -109.278632695019,
  -109.195814968555,
  -109.354679577894,
  -109.093405501977,
  -109.069026124649,
  -109.007024378249,
  -109.419287770971,
  1,
  0,
  -107.978896088346,
  0.136203094519617,
  -107.72060313008,
  -108.073680190789,
  -108.057380220448,
  -108.042668557136,
  -108.080524458934,
  -108.10770949901,
  -107.87672239732,
  -107.835030503412,
  -108.191106774667,
  -107.94798113767,
  -107.971822590539,
  -108.16244430587,
  -107.885117598383,
  -107.807966571223,
  -107.896004065362,
  -108.123928334196,
  -108.090803827731,
  -107.83104664343,
  -107.825739644628,
  -108.049641316089,
  1,
  0,
  -106.750934961131,
  0.139630341290287,
  -106.60801431385,
  -106.878177274089,
  -106.751399425817,
  -107.085820717804,
  -106.635740303236,
  -106.749258313595,
  -106.786823295456,
  -106.669598497066,
  -106.613420382887,
  -106.859091362244,
  -106.666080504262,
  -106.936586846683,
  -106.764218071939,
  -106.891326856401,
  -106.529996562331,
  -106.913650672126,
  -106.649999407852,
  -106.687980809298,
  -106.72568848184,
  -106.615827123851,
  1,
  0,
  -105.826660514651,
  0.140007364656364,
  -105.598143194886,
  -105.882617698802,
  -105.71714874633,
  -105.734287893661,
  -105.920528935133,
  -105.79541070349,
  -106.011000363316,
  -105.833460039022,
  -105.758340712246,
  -105.95115851039,
  -105.831815428451,
  -105.752233927322,
  -105.699583701352,
  -105.939337603334,
  -105.597258371819,
  -105.961159185903,
  -105.839556613284,
  -105.643190065258,
  -106.097010609602,
  -105.969967989421,
  1,
  0,
  -105.534990346254,
  0.139270831190724,
  -105.512727706325,
  -105.610408902782,
  -105.403558850898,
  -105.409274471279,
  -105.518666570934,
  -105.675320731105,
  -105.753807743472,
  -105.572827235104,
  -105.414180617683,
  -105.601861323954,
  -105.368408763256,
  -105.391847170187,
  -105.329039724434,
  -105.601386886981,
  -105.54137259462,
  -105.498712695307,
  -105.408471983469,
  -105.673305718441,
  -105.865397655127,
  -105.549229579717,
  1,
  0,
  -105.751523110409,
  0.144212891593613,
  -105.734427465046,
  -105.702536673948,
  -105.846066806624,
  -105.61920988783,
  -105.767163812781,
  -105.815368917991,
  -106.097582748855,
  -105.877228137895,
  -105.678832279916,
  -105.649845957878,
  -105.727441612827,
  -105.67496043744,
  -105.753097651285,
  -106.044535203608,
  -105.575655917871,
  -105.649518912652,
  -105.585687557386,
  -105.803886248867,
  -105.56576766728,
  -105.861648310199,
  1,
  0,
  -106.164230829878,
  0.147125312175089,
  -105.953047430949,
  -106.380340268568,
  -106.276954249257,
  -106.121964179106,
  -106.159583927439,
  -106.0530748954,
  -105.938588383205,
  -106.463608711996,
  -106.211947813947,
  -106.204687535031,
  -106.269495195269,
  -106.117168767247,
  -106.278521728668,
  -106.058100446883,
  -106.050146006156,
  -106.023736944998,
  -106.294771177214,
  -106.196049139526,
  -105.949617521188,
  -106.283212275514,
  1,
  0,
  -106.809756888776,
  0.147350272802327,
  -106.759660472741,
  -107.030305071611,
  -107.023618800115,
  -106.704464297553,
  -106.780872885141,
  -106.628766077986,
  -106.929379785268,
  -106.957021710136,
  -106.685253816871,
  -106.482857599082,
  -106.984110083639,
  -106.647451868627,
  -106.767498825883,
  -106.785440200032,
  -106.991135633495,
  -106.756968519483,
  -106.890525494533,
  -106.844635531075,
  -106.712189751842,
  -106.83298135041,
  1,
  0,
  -107.650447778967,
  0.150311692167309,
  -107.680579097686,
  -107.587842611443,
  -107.841371640897,
  -107.521456951503,
  -107.727122141504,
  -107.56023947669,
  -107.903049564276,
  -107.728417675952,
  -107.645302154844,
  -107.357208977176,
  -107.286625080557,
  -107.832199695564,
  -107.710019233982,
  -107.737969403283,
  -107.578467724528,
  -107.744236029524,
  -107.707800325337,
  -107.599197930184,
  -107.584666837874,
  -107.675183026533,
  1,
  0,
  -108.562902283195,
  0.154483990326421,
  -108.650924587819,
  -108.570033622086,
  -108.713080592031,
  -108.661737258094,
  -108.752141238129,
  -108.539376345347,
  -108.793379872882,
  -108.479174351309,
  -108.566200123852,
  -108.234955358026,
  -108.350263807571,
  -108.674209432154,
  -108.548548634903,
  -108.818399459208,
  -108.430775126851,
  -108.380799230114,
  -108.663229804137,
  -108.430716500654,
  -108.492398745917,
  -108.507701572807,
  1,
  0,
  -109.461982381104,
  0.155132759464222,
  -109.532205048069,
  -109.407734638683,
  -109.247419382136,
  -109.449702109907,
  -109.642874233138,
  -109.318044958354,
  -109.406968019093,
  -109.741352177581,
  -109.48192639562,
  -109.206662732068,
  -109.460709463363,
  -109.40286130899,
  -109.545828864129,
  -109.642565910449,
  -109.34913610475,
  -109.23032295729,
  -109.670959878689,
  -109.493730760655,
  -109.654808387508,
  -109.353834291612,
  1,
  0,
  -110.588250940235,
  0.160321765023609,
  -110.877336805136,
  -110.376865529926,
  -110.467364380391,
  -110.805455469996,
  -110.74220089733,
  -110.40467775254,
  -110.362941488477,
  -110.665493433477,
  -110.676325502849,
  -110.479314130465,
  -110.831218269216,
  -110.478705415306,
  -110.664078680964,
  -110.392530565444,
  -110.669014677372,
  -110.525743981704,
  -110.422230850651,
  -110.614489478511,
  -110.622853861159,
  -110.686177633796,
  1,
  0,
  -111.213179062113,
  0.165644825009741,
  -111.154303185466,
  -111.059528782712,
  -111.229750244746,
  -111.332267732459,
  -111.436156633559,
  -111.213899910096,
  -111.170996378665,
  -111.047524990246,
  -111.316681081043,
  -111.020327684357,
  -111.177123297947,
  -111.372997346236,
  -111.373345717966,
  -111.352395356107,
  -111.104967205183,
  -111.261706697667,
  -111.19059864128,
  -110.810555719418,
  -111.521589494695,
  -111.11686514241,
  1,
  0,
  -111.303874720853,
  0.166083030700782,
  -111.269828784745,
  -111.421487108714,
  -111.294518943189,
  -111.392623873776,
  -111.433616150612,
  -111.344228556785,
  -111.253066631786,
  -111.612941139597,
  -111.69336506052,
  -111.081987257424,
  -111.104216312529,
  -111.238595387635,
  -111.383812634915,
  -111.208156350214,
  -111.173865927404,
  -111.114478427969,
  -111.21707428117,
  -111.078637731086,
  -111.356284760998,
  -111.404709096003,
  1,
  0,
  -110.886374101018,
  0.167061511768366,
  -110.821986476638,
  -111.033443695987,
  -110.813826902531,
  -111.048077345359,
  -110.859007240363,
  -110.596146527915,
  -111.123944788325,
  -111.097992558927,
  -110.943817922874,
  -111.096186657875,
  -110.679620656013,
  -110.924095131331,
  -110.680748350954,
  -110.673794224517,
  -111.12871027047,
  -110.817652977298,
  -110.928222822065,
  -110.952241291619,
  -110.794817353614,
  -110.713148825677,
  1,
  0,
  -110.432137416396,
  0.171627236145908,
  -110.686119792614,
  -110.320784420821,
  -110.44094498016,
  -110.519016408003,
  -110.489559711004,
  -110.232814192251,
  -110.11590250984,
  -110.604410381823,
  -110.276878211099,
  -110.46899680369,
  -110.489888753038,
  -110.407141590908,
  -110.541508825908,
  -110.260735165733,
  -110.499724595525,
  -110.675182275656,
  -110.413775390295,
  -110.625193100146,
  -110.497239366434,
  -110.076931852977,
  1,
  0,
  -109.601814951796,
  0.178537120236353,
  -109.659654256363,
  -109.56184343699,
  -109.654588189461,
  -109.791236286766,
  -109.793145067066,
  -109.628325116372,
  -109.3949638948,
  -109.720671868806,
  -109.649478866807,
  -109.562569723479,
  -109.186569672783,
  -109.532106116359,
  -109.63454447945,
  -109.388445917543,
  -109.799944556647,
  -109.974515682301,
  -109.594452222033,
  -109.502732939623,
  -109.631011959775,
  -109.375498782497,
  1,
  0,
  -108.194925845463,
  0.182310227439666,
  -108.269655705174,
  -108.441904841738,
  -108.174254064242,
  -108.299453461389,
  -108.253683359531,
  -108.363398819622,
  -108.298792993708,
  -108.291389570419,
  -108.235374201927,
  -107.980741580298,
  -107.792778915568,
  -107.956299178911,
  -108.051462905492,
  -108.092824710347,
  -108.272561066282,
  -108.35958486884,
  -108.128241636283,
  -108.028929414385,
  -108.544110077183,
  -108.063075537927,
  1,
  0,
  -107.15280384857,
  0.185256383423902,
  -107.324703560955,
  -107.185799840801,
  -106.778131256128,
  -107.04467046265,
  -107.234280197742,
  -107.315734938329,
  -107.244640481854,
  -107.303016840287,
  -107.121969188571,
  -106.917364413311,
  -107.132385034571,
  -107.237502241275,
  -107.085492113104,
  -107.168801462874,
  -107.207640965432,
  -107.346299681587,
  -106.866807389327,
  -107.401229257985,
  -107.33313839491,
  -106.806469249715,
  1,
  0,
  -105.865440824429,
  0.190310695112627,
  -105.718949930517,
  -105.863501814985,
  -105.74903731548,
  -105.865257811341,
  -105.750579848178,
  -106.02719622497,
  -105.924046490514,
  -105.637033465438,
  -105.588453194059,
  -105.982722219571,
  -105.580060294431,
  -106.037181288684,
  -106.028240883969,
  -106.229274022001,
  -105.953269484538,
  -105.786643138955,
  -105.787603411496,
  -105.773784611924,
  -106.26394155175,
  -105.762039485777,
  1,
  0,
  -104.370677107165,
  0.194502084618676,
  -104.390359419419,
  -104.117882535052,
  -104.367733139468,
  -104.46219622866,
  -104.662168694068,
  -104.465022228753,
  -104.206149416311,
  -104.258520183669,
  -104.231455043497,
  -104.669899035605,
  -103.972197827115,
  -104.334274856574,
  -104.690110200232,
  -104.312774914637,
  -104.283789468356,
  -104.359595674053,
  -104.424549815717,
  -104.424087504676,
  -104.639360428159,
  -104.141415529271,
  1,
  0,
  -103.413487607465,
  0.192170569276824,
  -103.069872863097,
  -103.396977144576,
  -103.483419673408,
  -103.42835001895,
  -103.456997999404,
  -103.416591048829,
  -103.891815759927,
  -103.272444702311,
  -103.465356418359,
  -103.607242976788,
  -103.62790689223,
  -103.129912043134,
  -103.496543949815,
  -103.285181542865,
  -103.221215114616,
  -103.339221636526,
  -103.59570105398,
  -103.216939166613,
  -103.540021525079,
  -103.328040618788,
  1,
  0,
  -102.307256034107,
  0.196152672497485,
  -102.258122270594,
  -102.464524470686,
  -102.518749589841,
  -102.474235088979,
  -102.474497314418,
  -102.609062179017,
  -102.201546953192,
  -102.253991724443,
  -102.203753687241,
  -102.373271044408,
  -102.608224677228,
  -102.019956692908,
  -102.38646232088,
  -102.151223705869,
  -102.101200083882,
  -102.346371470267,
  -101.984152194283,
  -101.981515643712,
  -102.461308513696,
  -102.272951056591,
  1,
  0,
  -101.894215247166,
  0.204746597816553,
  -101.766644173879,
  -102.033167468745,
  -102.204803619726,
  -101.870128532931,
  -101.873693925779,
  -102.330775468055,
  -101.755033328669,
  -101.901506084601,
  -101.406901114925,
  -101.98574553902,
  -101.888796339051,
  -101.897594615207,
  -101.7196928443,
  -101.59580635826,
  -101.845247823764,
  -101.887629039803,
  -101.929721569939,
  -101.951737406947,
  -102.177114695708,
  -101.862564994013,
  1,
  0,
  -102.098054179428,
  0.211001748594732,
  -101.742637391465,
  -102.245928748461,
  -102.213394648615,
  -102.077236705833,
  -101.86582588675,
  -102.298845910169,
  -102.033713448981,
  -101.998303204074,
  -102.015563997539,
  -101.942560666315,
  -102.019244017164,
  -102.227360120039,
  -102.003390239425,
  -101.826094759836,
  -102.482363495814,
  -102.324782382819,
  -102.364722779783,
  -102.398004207996,
  -102.061014357239,
  -101.820096620243,
  1,
  0,
  -102.286459196417,
  0.206097769843535,
  -102.325899066329,
  -102.089122802783,
  -102.375486089785,
  -102.119443323062,
  -102.686292742123,
  -102.112367124249,
  -102.37767658938,
  -102.400259589765,
  -102.231888768051,
  -102.298161290479,
  -102.198289762751,
  -102.001045658322,
  -102.259803532608,
  -102.575840760375,
  -102.675440371557,
  -102.20393802758,
  -101.912524516404,
  -102.466441218798,
  -102.196543318278,
  -102.222719375651,
  1,
  0 ;
}
