netcdf perfect_input {
dimensions:
	member = 1 ;
	metadatalength = 32 ;
	Xlocation = 36 ;
	Ylocation = 360 ;
	time = UNLIMITED ; // (1 currently)
variables:

	char MemberMetadata(member, metadatalength) ;
		MemberMetadata:long_name = "description of each member" ;

	double Xlocation(Xlocation) ;
		Xlocation:short_name = "loc1d" ;
		Xlocation:long_name = "location on unit circle" ;
		Xlocation:dimension = 1 ;
		Xlocation:valid_range = 0., 1. ;

	double Ylocation(Ylocation) ;
		Xlocation:short_name = "loc1d" ;
		Ylocation:long_name = "location on unit circle" ;
		Ylocation:dimension = 1 ;
		Ylocation:valid_range = 0., 1. ;

	double X(time, member, Xlocation) ;
		X:long_name = "slow variables X" ;

	double Y(time, member, Ylocation) ;
		Y:long_name = "fast variables Y" ;

	double time(time) ;
		time:long_name = "valid time of the model state" ;
		time:axis = "T" ;
		time:cartesian_axis = "T" ;
		time:calendar = "none" ;
		time:units = "days" ;

// global attributes:
		:title = "true state from control" ;
                :version = "$Id: perfect_input.cdl 11431 2017-04-04 17:11:44Z hendric@ucar.edu $" ;
		:model = "Lorenz_96_2scale" ;
		:model_delta_t = 0.005 ;
		:model_coupling_b = 10. ;
		:model_coupling_c = 10. ;
		:model_coupling_h = 1. ;
		:model_forcing = 15. ;
                :history = "identical to r747 (circa June 2004)" ;
data:

 MemberMetadata =
  "true state" ;

 Xlocation = 0, 0.0277777777777778, 0.0555555555555556, 0.0833333333333333, 
    0.111111111111111, 0.138888888888889, 0.166666666666667, 
    0.194444444444444, 0.222222222222222, 0.25, 0.277777777777778, 
    0.305555555555556, 0.333333333333333, 0.361111111111111, 
    0.388888888888889, 0.416666666666667, 0.444444444444444, 
    0.472222222222222, 0.5, 0.527777777777778, 0.555555555555556, 
    0.583333333333333, 0.611111111111111, 0.638888888888889, 
    0.666666666666667, 0.694444444444444, 0.722222222222222, 0.75, 
    0.777777777777778, 0.805555555555556, 0.833333333333333, 
    0.861111111111111, 0.888888888888889, 0.916666666666667, 
    0.944444444444444, 0.972222222222222 ;

 Ylocation = 0, 0.00277777777777778, 0.00555555555555556, 
    0.00833333333333333, 0.0111111111111111, 0.0138888888888889, 
    0.0166666666666667, 0.0194444444444444, 0.0222222222222222, 0.025, 
    0.0277777777777778, 0.0305555555555556, 0.0333333333333333, 
    0.0361111111111111, 0.0388888888888889, 0.0416666666666667, 
    0.0444444444444444, 0.0472222222222222, 0.05, 0.0527777777777778, 
    0.0555555555555556, 0.0583333333333333, 0.0611111111111111, 
    0.0638888888888889, 0.0666666666666667, 0.0694444444444444, 
    0.0722222222222222, 0.075, 0.0777777777777778, 0.0805555555555556, 
    0.0833333333333333, 0.0861111111111111, 0.0888888888888889, 
    0.0916666666666667, 0.0944444444444444, 0.0972222222222222, 0.1, 
    0.102777777777778, 0.105555555555556, 0.108333333333333, 
    0.111111111111111, 0.113888888888889, 0.116666666666667, 
    0.119444444444444, 0.122222222222222, 0.125, 0.127777777777778, 
    0.130555555555556, 0.133333333333333, 0.136111111111111, 
    0.138888888888889, 0.141666666666667, 0.144444444444444, 
    0.147222222222222, 0.15, 0.152777777777778, 0.155555555555556, 
    0.158333333333333, 0.161111111111111, 0.163888888888889, 
    0.166666666666667, 0.169444444444444, 0.172222222222222, 0.175, 
    0.177777777777778, 0.180555555555556, 0.183333333333333, 
    0.186111111111111, 0.188888888888889, 0.191666666666667, 
    0.194444444444444, 0.197222222222222, 0.2, 0.202777777777778, 
    0.205555555555556, 0.208333333333333, 0.211111111111111, 
    0.213888888888889, 0.216666666666667, 0.219444444444444, 
    0.222222222222222, 0.225, 0.227777777777778, 0.230555555555556, 
    0.233333333333333, 0.236111111111111, 0.238888888888889, 
    0.241666666666667, 0.244444444444444, 0.247222222222222, 0.25, 
    0.252777777777778, 0.255555555555556, 0.258333333333333, 
    0.261111111111111, 0.263888888888889, 0.266666666666667, 
    0.269444444444444, 0.272222222222222, 0.275, 0.277777777777778, 
    0.280555555555556, 0.283333333333333, 0.286111111111111, 
    0.288888888888889, 0.291666666666667, 0.294444444444444, 
    0.297222222222222, 0.3, 0.302777777777778, 0.305555555555556, 
    0.308333333333333, 0.311111111111111, 0.313888888888889, 
    0.316666666666667, 0.319444444444444, 0.322222222222222, 0.325, 
    0.327777777777778, 0.330555555555556, 0.333333333333333, 
    0.336111111111111, 0.338888888888889, 0.341666666666667, 
    0.344444444444444, 0.347222222222222, 0.35, 0.352777777777778, 
    0.355555555555556, 0.358333333333333, 0.361111111111111, 
    0.363888888888889, 0.366666666666667, 0.369444444444444, 
    0.372222222222222, 0.375, 0.377777777777778, 0.380555555555556, 
    0.383333333333333, 0.386111111111111, 0.388888888888889, 
    0.391666666666667, 0.394444444444444, 0.397222222222222, 0.4, 
    0.402777777777778, 0.405555555555556, 0.408333333333333, 
    0.411111111111111, 0.413888888888889, 0.416666666666667, 
    0.419444444444444, 0.422222222222222, 0.425, 0.427777777777778, 
    0.430555555555556, 0.433333333333333, 0.436111111111111, 
    0.438888888888889, 0.441666666666667, 0.444444444444444, 
    0.447222222222222, 0.45, 0.452777777777778, 0.455555555555556, 
    0.458333333333333, 0.461111111111111, 0.463888888888889, 
    0.466666666666667, 0.469444444444444, 0.472222222222222, 0.475, 
    0.477777777777778, 0.480555555555556, 0.483333333333333, 
    0.486111111111111, 0.488888888888889, 0.491666666666667, 
    0.494444444444444, 0.497222222222222, 0.5, 0.502777777777778, 
    0.505555555555556, 0.508333333333333, 0.511111111111111, 
    0.513888888888889, 0.516666666666667, 0.519444444444444, 
    0.522222222222222, 0.525, 0.527777777777778, 0.530555555555556, 
    0.533333333333333, 0.536111111111111, 0.538888888888889, 
    0.541666666666667, 0.544444444444444, 0.547222222222222, 0.55, 
    0.552777777777778, 0.555555555555556, 0.558333333333333, 
    0.561111111111111, 0.563888888888889, 0.566666666666667, 
    0.569444444444444, 0.572222222222222, 0.575, 0.577777777777778, 
    0.580555555555556, 0.583333333333333, 0.586111111111111, 
    0.588888888888889, 0.591666666666667, 0.594444444444444, 
    0.597222222222222, 0.6, 0.602777777777778, 0.605555555555556, 
    0.608333333333333, 0.611111111111111, 0.613888888888889, 
    0.616666666666667, 0.619444444444444, 0.622222222222222, 0.625, 
    0.627777777777778, 0.630555555555556, 0.633333333333333, 
    0.636111111111111, 0.638888888888889, 0.641666666666667, 
    0.644444444444444, 0.647222222222222, 0.65, 0.652777777777778, 
    0.655555555555556, 0.658333333333333, 0.661111111111111, 
    0.663888888888889, 0.666666666666667, 0.669444444444444, 
    0.672222222222222, 0.675, 0.677777777777778, 0.680555555555556, 
    0.683333333333333, 0.686111111111111, 0.688888888888889, 
    0.691666666666667, 0.694444444444444, 0.697222222222222, 0.7, 
    0.702777777777778, 0.705555555555556, 0.708333333333333, 
    0.711111111111111, 0.713888888888889, 0.716666666666667, 
    0.719444444444444, 0.722222222222222, 0.725, 0.727777777777778, 
    0.730555555555556, 0.733333333333333, 0.736111111111111, 
    0.738888888888889, 0.741666666666667, 0.744444444444444, 
    0.747222222222222, 0.75, 0.752777777777778, 0.755555555555556, 
    0.758333333333333, 0.761111111111111, 0.763888888888889, 
    0.766666666666667, 0.769444444444444, 0.772222222222222, 0.775, 
    0.777777777777778, 0.780555555555556, 0.783333333333333, 
    0.786111111111111, 0.788888888888889, 0.791666666666667, 
    0.794444444444444, 0.797222222222222, 0.8, 0.802777777777778, 
    0.805555555555556, 0.808333333333333, 0.811111111111111, 
    0.813888888888889, 0.816666666666667, 0.819444444444444, 
    0.822222222222222, 0.825, 0.827777777777778, 0.830555555555556, 
    0.833333333333333, 0.836111111111111, 0.838888888888889, 
    0.841666666666667, 0.844444444444444, 0.847222222222222, 0.85, 
    0.852777777777778, 0.855555555555556, 0.858333333333333, 
    0.861111111111111, 0.863888888888889, 0.866666666666667, 
    0.869444444444444, 0.872222222222222, 0.875, 0.877777777777778, 
    0.880555555555556, 0.883333333333333, 0.886111111111111, 
    0.888888888888889, 0.891666666666667, 0.894444444444444, 
    0.897222222222222, 0.9, 0.902777777777778, 0.905555555555556, 
    0.908333333333333, 0.911111111111111, 0.913888888888889, 
    0.916666666666667, 0.919444444444444, 0.922222222222222, 0.925, 
    0.927777777777778, 0.930555555555556, 0.933333333333333, 
    0.936111111111111, 0.938888888888889, 0.941666666666667, 
    0.944444444444444, 0.947222222222222, 0.95, 0.952777777777778, 
    0.955555555555556, 0.958333333333333, 0.961111111111111, 
    0.963888888888889, 0.966666666666667, 0.969444444444444, 
    0.972222222222222, 0.975, 0.977777777777778, 0.980555555555556, 
    0.983333333333333, 0.986111111111111, 0.988888888888889, 
    0.991666666666667, 0.994444444444444, 0.997222222222222 ;


 X =
   6.92459281496202,       5.18944614769092,     -0.734668101492328,    
  -3.36395090822824,      0.771317245462520,       3.22052635628041,    
   8.46038185748605,       5.47720570567362,       1.14036447745838,    
   2.07714696413133,      -1.58454958227096,      0.637603193283668,    
   1.99018983215644,       7.43063825707261,       2.49122462361896,    
  -3.73639232697119,       1.20222154686682,       7.27904068928075,    
   2.05883916402944,      -1.46526913542259,       2.42886699642269,    
   8.61987581763088,      0.119048070826218,       3.29877394053497,    
   9.13527880607689,       1.81073688975838,      -3.91930785717331,    
   3.20541406557805,       2.45732162662538,      0.655228406897632,    
   2.36986271692554,       6.30762791401110,       3.17270392986682,    
  -3.62373423498127,       1.19079862292969E-002,  2.16029301556459;    

 Y =
  0.224432521103924,     -0.117977700944283,       7.40451803774910E-002,
  0.660580694013922,      0.177934413874730,      0.235596854879660,    
 -0.235995155421895,      0.415565621008921,      0.508480435651743,    
  0.292747494912127,       5.11874084422968E-002, 0.582319616509892,    
  0.284929988267817,      0.117138247137985,       7.24950859565485E-002,
 -0.106911682415420,      0.370927251274162,      0.381810746647892,    
   6.43622019936422E-002, 0.618643173742364,      0.454070611530201,    
  -1.89571223924732E-002, -6.18944876579952E-002,  4.90997908989822E-002,
   8.78733868172423E-002, 0.395227965481599,       3.88563722602217E-002,
  -5.13282138540228E-002,-0.152663163234591,       6.01112655443800E-002,
 -0.425710140225173,      -8.45785523190943E-002, -1.04791645875188E-002,
 -0.217763377635049,      0.264288385013975,     -0.233546075038151,    
   1.84314853016578E-002, -6.66333904327314E-002,  4.61857050652470E-002,
 -0.313860280404747,      -4.62628396293726E-003,  4.34900122734427E-002,
   7.00121308593608E-002,  7.18975424245294E-002,  8.06886535626838E-002,
   3.73765049277144E-002,  2.98449595284551E-002, 0.103706911269968,    
  0.101739494226607,      -1.41693539199238E-003, 0.136927519968663,    
  0.201699226279513,      0.128880288681680,      0.100526169462929,    
  0.221839416535660,      0.143676722244464,      0.129714099183696,    
  0.465799705374190,      0.113285888810172,      -3.97511503995684E-002,
 -0.136913390984165,     -0.200463434933559,      0.744824539064179,    
  0.165128196893027,      -7.59845292167713E-002, 0.204474007675176,    
  0.502827754343558,     -0.101704311374852,      0.395967340515197,    
  0.854161102826061,       3.06122752324456E-002, -4.52616336773969E-002,
 -0.286592262547232,      0.680196176571713,      0.444699841047437,    
   6.95935171452701E-002,-0.214531259538855,       3.74984160429829E-002,
  0.503414046479722,      0.169216725781232,      -2.16932250051066E-002,
  -9.79230628545002E-002, 0.132057367913642,      0.291204804571101,    
  0.213554952111379,       8.55507841852337E-002, -3.81983351114271E-002,
   2.74300734057200E-002, 0.424330723788343,       7.62786203780202E-002,
   8.54820750172568E-002, -9.43337371323792E-002, 0.139678814618251,    
  0.304294249989458,       9.28314264079216E-002,-0.214966037369788,    
  0.130749713312603,      0.351947313222858,      -9.92999372948604E-002,
  -2.55176192131475E-002, -3.72509580680935E-002,-0.147424189304364,    
   9.97599172902704E-002,-0.149145229779087,       8.65342884755684E-002,
  -8.70649239328766E-002,  9.75811914357728E-002, -5.69791465109883E-002,
  0.114510166848968,     -0.108186545354392,      0.100768127955385,    
  -4.69320508414132E-002,  1.17123350027525E-002,  9.41312556663959E-003,
   5.17809574223413E-002,  3.61860988955552E-003,  5.32867156300316E-002,
   1.24986299549605E-002,  2.55124197549822E-002, -4.69178216943116E-002,
  -5.67261664781371E-003,  7.85812296405595E-002, 0.127394203201273,    
   9.28964698798237E-002,  5.08036754137642E-002,  2.06636843160756E-002,
  0.219285666962024,      0.195467520321880,      -1.22314167332399E-002,
  -4.55648075364063E-002, 0.312231904491472,     -0.244722577203520,    
  0.434059281985333,      0.568943149178911,      0.230447113431532,    
  -8.00674579173659E-002, 0.366732164983327,      0.235912391990593,    
   6.10871211987698E-002, 0.821482356682007,      0.476233507075293,    
  0.165230835649621,       8.62467922116348E-002,  3.77967209906622E-002,
  0.179145492371661,      0.222970900097230,      0.428414997573646,    
  0.240750905649538,     -0.297078507712352,       1.95373588366697E-002,
 -0.380702376408910,      -7.92407369020183E-002,-0.322456909810116,    
 -0.132596959738645,     -0.303791255508148,     -0.186104860797704,    
 -0.156228340513879,     -0.258579712603680,       4.76624675207858E-003,
 -0.278241468406248,      -3.90292812461024E-002,  5.39485308885602E-002,
   9.31792559461444E-002, 0.109251789160797,      0.100782917620003,    
   8.05106979593330E-002, 0.155963845981198,      0.146030286635063,    
  -2.83057652781254E-002, 0.183088268616798,      0.396028466697685,    
   1.25948361426566E-002,-0.166158400960806,      -9.26727569564734E-002,
  0.578173589941296,      0.361876250737580,      0.172059367356281,    
  0.234175127204663,      0.246114366279909,      -6.74339904648598E-002,
  0.246946359557819,      0.493565112438214,      0.248995817398965,    
  0.225021783214620,      0.341531297120857,      0.164473679597543,    
  -4.38833476148314E-002, 0.400469184085261,       8.06477202866208E-002,
  -3.52334635249885E-002,-0.111432193576759,     -0.140256304806129,    
   2.19234944558397E-002,-0.104496606976159,       4.28268859233963E-002,
 -0.138609089286285,       3.44767576315804E-002, -7.86777220715177E-002,
   8.71667683903911E-002, -8.68822928568737E-002, 0.184708690026321,    
   5.80404294082929E-002,  5.76109873918491E-002, 0.333223490522940,    
  0.170062443818334,      -6.38370888227849E-003, 0.349071131492725,    
  0.199001318468835,      -3.73824096389631E-002, -3.78189176343669E-003,
  0.555403613348991,      0.194521130052569,      0.570167820069662,    
  0.542977118115411,      0.190449242403077,      0.475620718892240,    
  0.528288107641288,      0.108383875792133,       1.04917280963676,    
  0.479604537745082,      -9.47168340598789E-002, -2.01654473136064E-002,
  -1.78972775144705E-002,  2.30939356126830E-002,-0.102684483504156,    
  -2.31607440590574E-003, -5.74240069396230E-002, -7.01793300226932E-002,
  0.109723987934054,     -0.111662854362618,       1.25752548923928E-002,
  0.155295572529050,      0.148173938508701,      0.112789239969945,    
   4.23795852987171E-002, 0.235349636061600,      0.498444088149931,    
   9.30046289675746E-002, -3.64410738765458E-002,-0.332209807036945,    
  0.447841326725433,      0.554773157467589,      0.162696397884749,    
 -0.305147968192891,       2.99937756640925E-002,  1.13781191489187,    
 -0.103513826636251,     -0.259286713339798,      0.188987504382684,    
  0.547302584019189,      -4.70947208740894E-002,  1.52958279862078E-002,
 -0.256154980593783,       8.16774848913060E-002, 0.385916368673864,    
  0.644241467115758,      0.273616495322719,      -5.24693965035327E-002,
  0.249479771320380,       3.02493091127641E-002,-0.371846934272228,    
  0.156104293813474,     -0.392212865873898,      -9.55925449783234E-002,
 -0.325976300546424,     -0.181314020346794,     -0.248213801063953,    
 -0.235427192752993,     -0.124331645107166,     -0.168260843940050,    
 -0.100409824899133,      0.117218883842394,      0.181888489263522,    
  0.124518026479678,      0.122401871749198,      0.202157465625687,    
  0.181966931644561,      0.140437710415964,      0.206912926391646,    
  0.221958956067875,      0.144458204790649,      0.122293271540285,    
  0.102467938468852,      0.105636137164089,       9.73373291180083E-002,
   9.91674175726647E-002, 0.101256662332830,      0.101759467988869,    
  0.128914744905133,       9.77696049948057E-002,  1.95169241814911E-002,
   1.91829000261203E-002,  4.27074153758634E-002,  3.22753943049854E-002,
   4.68451852638804E-002, -2.26371491934525E-002,  2.16221028840861E-002,
   2.63643223920289E-002,  4.74034585259527E-002, -3.37766153152093E-002,
   5.30394328716275E-002,  9.62878059833788E-002,  8.35747109692443E-002,
  0.155267317919757,      0.209553751177948,      0.123167059298294,    
   4.64570588663667E-002, 0.160843303573401,      0.234132189899344,    
  0.231566129588758,      0.200111545411795,       3.24284355172951E-002,
 -0.111366335769921,      -1.85573352161956E-002, 0.300155424040906,    
  0.692525370691293,      0.305192336609652,     -0.146798298270568,    
  0.270445171502140,      0.610039127972276,      0.118292301221938,    
  -9.02677380313017E-002, 0.225935130132372,      0.196348193272061,    
   5.22210881134674E-003,-0.138259787972273,      0.471998675301529,    
  0.711980017987835,      -6.50631113321427E-002,-0.195070360387866,    
 -0.323700885023372,       1.66408000652290E-002,-0.349592952721931,    
  -9.44592477271842E-002,-0.299001985591117,     -0.165678106414459,    
 -0.180364562470433,     -0.195806365613163,     -0.135530260455869,    
 -0.147351545570104,      -3.81966029140642E-002,  9.33370979952939E-002,
 -0.204218620276250,      -3.10701948841294E-002, -1.46497228629672E-002,
 -0.157900763435040,      -3.54446759470129E-003,  4.15387648649483E-002,
   5.23825254266018E-002,-0.136737229828985,       3.92205267664100E-002,
   8.52035554792090E-002,  5.28787333579182E-002, 0.148588047745194,    
  0.236527979671467,      0.139211753346888,       4.41278186243963E-002,
  -1.40518316924299E-002,  5.62282203375254E-002, 0.492322048628986 ;    

 time = 1000.0 ;

}

