netcdf sqgRestart {
dimensions:
	nx = 128 ;
	ny = 64 ;
	nz = 2 ;
	time = UNLIMITED ; // (1 currently)
variables:
	float time(time) ;
	float theta(time, nz, ny, nx) ;
		theta:description = "potential temperature" ;

// global attributes:
		:model = 1 ;
		:ntims = 1000001 ;
		:dt = 0.01f ;
		:iplot = 1000 ;
		:XL = 20.f ;
		:YL = 11.07824f ;
		:H = 1.f ;
		:Ross = 0.f ;
		:gamma = 0.f ;
		:n = 8 ;
		:tau = 0.2f ;
		:trl = 15.f ;
		:amu = 1.f ;
		:shear = 1.f ;
data:

 time = 0 ;

 theta =
  -0.2131442, -0.2042771, -0.1928141, -0.1809788, -0.1685103, -0.1531882, 
    -0.1378816, -0.1225994, -0.105348, -0.08823985, -0.07320794, -0.05902185, 
    -0.04346127, -0.02667645, -0.009235702, 0.007921606, 0.02370197, 
    0.03735104, 0.04883482, 0.05922294, 0.06847094, 0.07534771, 0.0819956, 
    0.09035011, 0.098269, 0.1035984, 0.1066184, 0.1097822, 0.1112651, 
    0.1079242, 0.1012594, 0.09411213, 0.08731365, 0.08029756, 0.07007831, 
    0.05519614, 0.04132921, 0.03268161, 0.02812767, 0.02250469, 0.01224202, 
    0.001214802, -0.00898546, -0.01799285, -0.02158374, -0.02260113, 
    -0.02561137, -0.03428957, -0.04959531, -0.0739508, -0.0983322, 
    -0.1124575, -0.1168989, -0.1157231, -0.1130084, -0.1083387, -0.100089, 
    -0.08931525, -0.07786039, -0.06612384, -0.05647705, -0.05009718, 
    -0.04262479, -0.0310514, -0.01465406, 0.01123502, 0.03949683, 0.06337157, 
    0.08482486, 0.10222, 0.113451, 0.1229797, 0.1319919, 0.1390255, 
    0.1414867, 0.1384824, 0.1302225, 0.1176693, 0.1038053, 0.09295237, 
    0.0800283, 0.06218907, 0.04309601, 0.02252457, 0.003306001, -0.01107559, 
    -0.01788871, -0.01846191, -0.01618016, -0.01428542, -0.01382303, 
    -0.009270489, 0.001432121, 0.01421255, 0.02829114, 0.04227453, 0.0552102, 
    0.06657246, 0.07626745, 0.08503187, 0.09235254, 0.09570417, 0.09455863, 
    0.09165144, 0.08704551, 0.07898918, 0.06855526, 0.05533097, 0.03945107, 
    0.02155134, 0.001563668, -0.02038947, -0.0435221, -0.06615068, 
    -0.08764049, -0.1079811, -0.1286594, -0.1494841, -0.1697769, -0.1886726, 
    -0.2052938, -0.2191008, -0.2286627, -0.2339033, -0.2350251, -0.2322058, 
    -0.2267151, -0.2201372,
  -0.2140687, -0.2048985, -0.193144, -0.180759, -0.1677208, -0.1522996, 
    -0.1366353, -0.1204167, -0.1037205, -0.08756901, -0.07175411, -0.0571555, 
    -0.04210515, -0.02525733, -0.007857867, 0.00883083, 0.02474095, 
    0.0382518, 0.04910998, 0.05907273, 0.06838875, 0.07601531, 0.08298679, 
    0.08989589, 0.09620343, 0.1020504, 0.1070423, 0.1109859, 0.1115523, 
    0.1085269, 0.1047691, 0.1010437, 0.09579873, 0.08795434, 0.07506424, 
    0.05643618, 0.03811944, 0.02423087, 0.01365539, 0.005244344, 
    -0.001338273, -0.007521868, -0.01663086, -0.02680133, -0.03027111, 
    -0.02885731, -0.02965117, -0.03594542, -0.04834956, -0.07065338, 
    -0.09513118, -0.1107818, -0.1169072, -0.1173417, -0.1147285, -0.1079573, 
    -0.09772718, -0.0861646, -0.07450635, -0.06316739, -0.05372323, 
    -0.04749328, -0.03949405, -0.02543199, -0.006606862, 0.01579162, 
    0.04195794, 0.06896937, 0.08768928, 0.1009125, 0.1130481, 0.1233782, 
    0.1320139, 0.1368907, 0.1369048, 0.1334838, 0.1302359, 0.1270041, 
    0.1153351, 0.09360102, 0.0698649, 0.04773059, 0.02605629, 0.009428561, 
    -0.0004813969, -0.008828431, -0.01761924, -0.02709611, -0.03667977, 
    -0.03863788, -0.02652767, -0.005099326, 0.01582804, 0.03154618, 
    0.04455751, 0.05628929, 0.06730503, 0.07714653, 0.08496842, 0.09044868, 
    0.09411436, 0.09715369, 0.09934111, 0.09779902, 0.09286264, 0.08606277, 
    0.07499842, 0.06063438, 0.04468045, 0.02586779, 0.004796281, -0.01652928, 
    -0.03881953, -0.0628827, -0.08597601, -0.1069065, -0.1272633, -0.1485872, 
    -0.1695823, -0.1891868, -0.2067611, -0.220241, -0.2297866, -0.235085, 
    -0.2361024, -0.2334127, -0.2279867, -0.2213802,
  -0.2146479, -0.205252, -0.193273, -0.1807739, -0.1677956, -0.15216, 
    -0.1364541, -0.1206901, -0.1031929, -0.0860477, -0.07083981, -0.05635466, 
    -0.04061483, -0.02382647, -0.006375343, 0.01099668, 0.0268625, 
    0.04009933, 0.0512149, 0.06154498, 0.07048912, 0.07698369, 0.08373129, 
    0.09237549, 0.1002318, 0.1049866, 0.1075275, 0.1103524, 0.1113686, 
    0.1084323, 0.1029136, 0.09644006, 0.08910891, 0.08082992, 0.06923926, 
    0.05306619, 0.03859526, 0.03061488, 0.02732952, 0.02238505, 0.0122841, 
    0.001246765, -0.009718329, -0.01977806, -0.02371563, -0.02496049, 
    -0.02873902, -0.03827214, -0.05376562, -0.07741851, -0.1004228, 
    -0.1126763, -0.1153311, -0.1129796, -0.1093076, -0.1036737, -0.09457869, 
    -0.08282397, -0.07032061, -0.05885545, -0.0501513, -0.04274859, 
    -0.03375909, -0.02197118, -0.005273104, 0.01992954, 0.04646587, 
    0.06864947, 0.08840694, 0.1042364, 0.1140194, 0.1225853, 0.131142, 
    0.1378831, 0.1405176, 0.1397071, 0.1340774, 0.1205856, 0.1022592, 
    0.08752495, 0.07415342, 0.05896696, 0.0446457, 0.0294733, 0.01284096, 
    -0.003249317, -0.01293205, -0.0153084, -0.01396103, -0.01261582, 
    -0.01283339, -0.008618802, 0.002759874, 0.01675081, 0.03161997, 
    0.04591769, 0.05909196, 0.07055169, 0.08020365, 0.08901083, 0.09647411, 
    0.1001765, 0.09961411, 0.09731391, 0.09328346, 0.08575369, 0.07630602, 
    0.0645967, 0.04974141, 0.03204578, 0.01241418, -0.009096242, -0.0331252, 
    -0.05780755, -0.08093379, -0.1020597, -0.1237405, -0.1464947, -0.1688706, 
    -0.1890859, -0.206774, -0.221434, -0.2313749, -0.2368573, -0.237885, 
    -0.2347233, -0.2289428, -0.2221155,
  -0.2158448, -0.2063133, -0.193993, -0.1809505, -0.1672841, -0.1514219, 
    -0.1355482, -0.1190108, -0.1018792, -0.0855823, -0.0696862, -0.05482815, 
    -0.03959808, -0.0227257, -0.005232096, 0.01158798, 0.02735064, 
    0.04052465, 0.0514159, 0.06170808, 0.07107185, 0.07850677, 0.08520278, 
    0.09161313, 0.09740371, 0.1028877, 0.1079149, 0.1120413, 0.1125532, 
    0.1093228, 0.1046986, 0.09983316, 0.09413871, 0.08667587, 0.07474139, 
    0.0578396, 0.04117021, 0.02744226, 0.01607597, 0.006625965, -0.001379088, 
    -0.009048894, -0.01903996, -0.02913462, -0.03225432, -0.03094694, 
    -0.03236999, -0.03966673, -0.05270502, -0.07435239, -0.09656037, 
    -0.1088139, -0.1118762, -0.1107087, -0.1070447, -0.09954292, -0.08974873, 
    -0.0784705, -0.0663941, -0.05583154, -0.04794847, -0.04148182, 
    -0.03284292, -0.01899296, -0.0003433451, 0.02147102, 0.04641777, 
    0.07202713, 0.08994506, 0.1023905, 0.113656, 0.1236826, 0.1328397, 
    0.1383411, 0.1382709, 0.1339214, 0.1288221, 0.1249382, 0.1162908, 
    0.0991787, 0.07803591, 0.05559042, 0.03081241, 0.007981867, -0.007671505, 
    -0.01642224, -0.02173744, -0.02831118, -0.03585844, -0.03535813, 
    -0.02107456, 0.0013372, 0.02216861, 0.0374126, 0.04993123, 0.06161214, 
    0.07298912, 0.08289787, 0.09033185, 0.09558617, 0.09940761, 0.1027621, 
    0.1054169, 0.1046118, 0.1005205, 0.09490006, 0.08539751, 0.07211743, 
    0.05694018, 0.03952938, 0.01934385, -0.002725963, -0.02583983, 
    -0.05006234, -0.07413391, -0.09688514, -0.1185971, -0.1416037, 
    -0.1653458, -0.1873729, -0.2068043, -0.2220169, -0.2326596, -0.2384557, 
    -0.2395556, -0.2364989, -0.2303635, -0.2233007,
  -0.2165613, -0.2067152, -0.1941592, -0.1810308, -0.1676537, -0.1515875, 
    -0.1355671, -0.1195321, -0.1015949, -0.08418047, -0.06891245, 
    -0.05424666, -0.03821485, -0.02135123, -0.003943726, 0.01364616, 
    0.02965265, 0.04250617, 0.05323662, 0.06349999, 0.07238995, 0.07887714, 
    0.08568254, 0.09427942, 0.1019845, 0.106383, 0.1085004, 0.1107677, 
    0.111035, 0.1078407, 0.1027744, 0.09712529, 0.09042838, 0.08214974, 
    0.06959292, 0.05178995, 0.03581382, 0.02730359, 0.02437685, 0.01979391, 
    0.0101088, -0.0004957691, -0.01154355, -0.02157664, -0.02512325, 
    -0.02712084, -0.03283917, -0.04370541, -0.05871348, -0.07952473, 
    -0.09747262, -0.1029473, -0.09994461, -0.09547082, -0.0917844, 
    -0.08718109, -0.07994524, -0.07055261, -0.06038821, -0.05116367, 
    -0.04363094, -0.03586448, -0.02681826, -0.01581407, -0.0001665279, 
    0.02391365, 0.04972224, 0.07109692, 0.08992179, 0.1053931, 0.1150853, 
    0.1235587, 0.1318142, 0.1382614, 0.1411529, 0.1416994, 0.1382128, 
    0.1263402, 0.1069265, 0.08761993, 0.06960529, 0.05259672, 0.03925982, 
    0.02895816, 0.01993249, 0.007667884, -0.00395152, -0.01004648, 
    -0.01142265, -0.01155952, -0.01257402, -0.008177757, 0.004551291, 
    0.02024032, 0.03632797, 0.05124164, 0.06456055, 0.07597647, 0.08556962, 
    0.09435464, 0.1019285, 0.1060784, 0.1062274, 0.1047958, 0.1019174, 
    0.09554808, 0.08737711, 0.07768892, 0.06556065, 0.04973656, 0.02997772, 
    0.008746795, -0.01374565, -0.03895686, -0.06563538, -0.09033421, 
    -0.1140527, -0.139017, -0.1648481, -0.1880145, -0.2072327, -0.2230268, 
    -0.2339157, -0.2399934, -0.2412538, -0.2383645, -0.2325306, -0.224856,
  -0.2182244, -0.2080833, -0.195186, -0.1813809, -0.1673877, -0.1512447, 
    -0.1348904, -0.1179392, -0.100373, -0.08382905, -0.06787711, -0.05292253, 
    -0.03749359, -0.02044275, -0.002829909, 0.01404166, 0.02967916, 0.042644, 
    0.05369397, 0.06434369, 0.07360157, 0.08058795, 0.08704709, 0.09341933, 
    0.09896408, 0.1038434, 0.1085339, 0.1127935, 0.1133877, 0.1099706, 
    0.1048893, 0.09954607, 0.09327583, 0.08503243, 0.07291177, 0.05744311, 
    0.04299627, 0.0304929, 0.01924703, 0.009418778, 0.0002008006, 
    -0.009196118, -0.02022529, -0.02966754, -0.03150485, -0.03079634, 
    -0.03405161, -0.04262362, -0.054564, -0.07153502, -0.08435698, 
    -0.08530094, -0.08311191, -0.08206955, -0.0792684, -0.0730012, 
    -0.06494578, -0.05625577, -0.04869838, -0.04296032, -0.03773393, 
    -0.03231367, -0.02484033, -0.01218674, 0.005265072, 0.0255298, 
    0.04905331, 0.07363129, 0.09117585, 0.103498, 0.1147998, 0.1248873, 
    0.1342862, 0.1404423, 0.1409755, 0.1361751, 0.1290612, 0.1227919, 
    0.1137486, 0.09959755, 0.08351348, 0.06514978, 0.04264781, 0.01788904, 
    -0.006460473, -0.02359577, -0.02955092, -0.03236508, -0.03573389, 
    -0.03089203, -0.01330921, 0.01053746, 0.03149758, 0.04609187, 0.05806664, 
    0.06991187, 0.08151627, 0.09123646, 0.09816079, 0.103151, 0.1071764, 
    0.1111399, 0.114604, 0.114673, 0.1115689, 0.1075706, 0.1005347, 
    0.08982928, 0.07663437, 0.06068977, 0.04223812, 0.02231565, 
    -0.0004690103, -0.02701596, -0.05454101, -0.08110423, -0.1061819, 
    -0.1317799, -0.1591083, -0.1858048, -0.2081101, -0.2244216, -0.2356749, 
    -0.2415504, -0.242305, -0.2389342, -0.2329676, -0.2261263,
  -0.2182848, -0.2083503, -0.1955304, -0.1817972, -0.1678009, -0.1511906, 
    -0.1346239, -0.1183767, -0.1002961, -0.0826298, -0.06719351, -0.05246329, 
    -0.03610629, -0.01889727, -0.001550928, 0.01585831, 0.03193939, 
    0.04490508, 0.05550183, 0.06537431, 0.07410917, 0.08100843, 0.08807692, 
    0.09622087, 0.10345, 0.1080177, 0.110486, 0.1124136, 0.1118986, 
    0.1084414, 0.1034765, 0.09771003, 0.09097684, 0.08318214, 0.0710808, 
    0.05268069, 0.03482619, 0.02448235, 0.02070859, 0.01591247, 0.006528487, 
    -0.003472839, -0.0143202, -0.02299903, -0.0251588, -0.0289017, 
    -0.03743809, -0.04865669, -0.05817487, -0.06681505, -0.0661388, 
    -0.0579656, -0.05298369, -0.04967682, -0.0474395, -0.04629518, 
    -0.04412502, -0.04066655, -0.03703137, -0.03264551, -0.02713923, 
    -0.020321, -0.01327865, -0.005065233, 0.007307768, 0.02857126, 0.0528558, 
    0.07327756, 0.09116185, 0.1063554, 0.1165242, 0.1257165, 0.1339203, 
    0.1398342, 0.1426278, 0.1436753, 0.1417947, 0.1329687, 0.1164372, 
    0.09609698, 0.07278322, 0.04986933, 0.03126527, 0.01737013, 0.01269235, 
    0.01128411, 0.005789235, -0.001809806, -0.00657019, -0.009320371, 
    -0.01259733, -0.00868196, 0.006237425, 0.02467119, 0.04291845, 
    0.05940091, 0.07311593, 0.08424369, 0.09370244, 0.1024436, 0.1100025, 
    0.1145467, 0.115472, 0.1151396, 0.1139659, 0.1096169, 0.103696, 
    0.0969912, 0.08867281, 0.07708336, 0.0605755, 0.03962747, 0.0153767, 
    -0.01036514, -0.03763457, -0.06634912, -0.09506323, -0.1230324, 
    -0.151674, -0.1787817, -0.2025117, -0.2225002, -0.2364914, -0.2440274, 
    -0.245228, -0.2415403, -0.2344318, -0.2262591,
  -0.2195531, -0.2091764, -0.1961542, -0.1818397, -0.167136, -0.1506206, 
    -0.1340994, -0.1168862, -0.09900266, -0.08233568, -0.06605917, 
    -0.05070981, -0.03527117, -0.01841593, -0.0007437319, 0.01647878, 
    0.03226985, 0.04498312, 0.05581442, 0.06664616, 0.07612623, 0.08293763, 
    0.08888586, 0.09503487, 0.1007022, 0.1053662, 0.1092092, 0.1127848, 
    0.1133953, 0.1101696, 0.1047841, 0.09927229, 0.09335296, 0.08518973, 
    0.07238692, 0.05672196, 0.04389739, 0.03380792, 0.0239287, 0.01455152, 
    0.004185496, -0.007654823, -0.02010359, -0.02736326, -0.02827641, 
    -0.03145137, -0.03652869, -0.03758008, -0.0364764, -0.03942682, 
    -0.03953949, -0.03872417, -0.03754286, -0.0331588, -0.02604838, 
    -0.01787218, -0.01209179, -0.008552641, -0.006831035, -0.006819084, 
    -0.007421479, -0.007516176, -0.005199671, 0.00331971, 0.01712629, 
    0.03365768, 0.05342212, 0.0758734, 0.09279159, 0.1050143, 0.1166693, 
    0.127261, 0.1367545, 0.1432464, 0.1449065, 0.1412575, 0.1337882, 
    0.124805, 0.1114343, 0.09462553, 0.0809913, 0.06788485, 0.05141594, 
    0.03516462, 0.01403928, -0.01225461, -0.02870706, -0.03371919, 
    -0.0339253, -0.02363168, 9.345263e-05, 0.02859505, 0.05019559, 
    0.06273089, 0.07305606, 0.08407618, 0.09486666, 0.1031865, 0.1098104, 
    0.1157173, 0.1203294, 0.1247114, 0.1291064, 0.1307897, 0.1294162, 
    0.1272645, 0.122862, 0.1154191, 0.105389, 0.09257203, 0.07697581, 
    0.05824266, 0.03570479, 0.01020467, -0.01802769, -0.05061299, 
    -0.08328235, -0.1128693, -0.1413886, -0.1706894, -0.1982307, -0.2192982, 
    -0.234651, -0.2436812, -0.2453014, -0.2424619, -0.2367638, -0.2285162,
  -0.219483, -0.2092427, -0.1954504, -0.1809292, -0.1670147, -0.1502052, 
    -0.1332775, -0.1172667, -0.09894347, -0.08056754, -0.06494325, 
    -0.05052549, -0.03417385, -0.01648596, 0.001195461, 0.01848224, 
    0.03421549, 0.04701654, 0.05780936, 0.06781762, 0.07624972, 0.08296715, 
    0.09024829, 0.09853835, 0.1055005, 0.1099329, 0.1125689, 0.1147452, 
    0.1142583, 0.1105161, 0.1051165, 0.09935789, 0.09285665, 0.08518998, 
    0.07380985, 0.05675575, 0.03846586, 0.0253233, 0.0183801, 0.01149415, 
    0.001040459, -0.008784261, -0.01883335, -0.0253107, -0.02878769, 
    -0.03338837, -0.03398322, -0.03628956, -0.04627426, -0.05588323, 
    -0.05636351, -0.05360105, -0.05018102, -0.04861586, -0.04864871, 
    -0.04743235, -0.04233369, -0.03285058, -0.0195103, -0.003999978, 
    0.01099318, 0.02125444, 0.02524418, 0.02492961, 0.02726215, 0.04066715, 
    0.06009895, 0.07759517, 0.09375957, 0.1083857, 0.1184686, 0.1284438, 
    0.136983, 0.1426233, 0.1451335, 0.1455076, 0.1429155, 0.1353745, 
    0.1235304, 0.108817, 0.08688705, 0.05992251, 0.03548764, 0.01151986, 
    -0.007472597, -0.01181585, -0.007471725, -0.008064926, -0.01173867, 
    -0.01678022, -0.02464011, -0.02031559, 4.917383e-05, 0.02459894, 
    0.05013014, 0.07129669, 0.08663115, 0.09882398, 0.1079828, 0.1147962, 
    0.1208766, 0.1255027, 0.1273199, 0.1284748, 0.1294942, 0.1280082, 
    0.1252331, 0.1218487, 0.1174818, 0.1106345, 0.09862595, 0.08025765, 
    0.05667573, 0.03035398, 0.0009545982, -0.03407733, -0.07197374, 
    -0.1042776, -0.1337756, -0.1652416, -0.1952319, -0.2187989, -0.2344449, 
    -0.243282, -0.2448684, -0.2411859, -0.2353894, -0.2278303,
  -0.2182912, -0.2082605, -0.1952288, -0.1796065, -0.1647376, -0.1494123, 
    -0.1326156, -0.1143982, -0.09647804, -0.08001429, -0.06360465, 
    -0.04828703, -0.03279543, -0.0155912, 0.002201051, 0.01907641, 
    0.03471022, 0.04779107, 0.05875118, 0.06909639, 0.07829513, 0.08547332, 
    0.09160133, 0.09718838, 0.1022469, 0.1071034, 0.1112157, 0.1142774, 
    0.1142685, 0.1111577, 0.1063316, 0.1010562, 0.09528706, 0.08822948, 
    0.07675149, 0.06010362, 0.04561916, 0.03710851, 0.02969873, 0.02147588, 
    0.01104023, -0.003572106, -0.01831466, -0.02451947, -0.02493937, 
    -0.02308164, -0.02888855, -0.04770572, -0.0649039, -0.07638395, 
    -0.08986683, -0.1064, -0.1192836, -0.129008, -0.1358162, -0.1399198, 
    -0.1400858, -0.1342794, -0.1225909, -0.1047959, -0.07947734, -0.04736432, 
    -0.01050961, 0.02454346, 0.04765242, 0.05695766, 0.0660584, 0.082753, 
    0.09752181, 0.1085457, 0.1199969, 0.130978, 0.1410416, 0.1473137, 
    0.149288, 0.1476732, 0.1429884, 0.1353383, 0.1194969, 0.09580619, 
    0.07509507, 0.05945754, 0.0440806, 0.03235836, 0.02721919, 0.01939487, 
    0.005469441, -0.003969774, -0.001098096, 0.01634816, 0.04363696, 
    0.070679, 0.08602346, 0.09129554, 0.09690616, 0.1027485, 0.1076731, 
    0.114936, 0.1244435, 0.1332415, 0.1395372, 0.1439245, 0.1471451, 
    0.1477154, 0.1458132, 0.1437508, 0.1406993, 0.1359792, 0.1287705, 
    0.1186799, 0.1066437, 0.09254877, 0.07376701, 0.04895113, 0.01930478, 
    -0.01669636, -0.05577512, -0.09093903, -0.1234584, -0.1600223, 
    -0.1954809, -0.2208449, -0.2364617, -0.2439, -0.2442626, -0.2390577, 
    -0.2326362, -0.226336,
  -0.2153625, -0.2039865, -0.1906769, -0.1782523, -0.1636516, -0.1453524, 
    -0.1295536, -0.1145026, -0.09568858, -0.077425, -0.06203035, -0.04700914, 
    -0.03024, -0.01310042, 0.004014969, 0.02170005, 0.03778951, 0.04999574, 
    0.06016666, 0.07040183, 0.07928558, 0.08571614, 0.09220722, 0.1004709, 
    0.1082198, 0.1130023, 0.1150111, 0.1168238, 0.1171461, 0.114193, 
    0.108768, 0.1028682, 0.09723505, 0.09094818, 0.0806849, 0.06488448, 
    0.04810365, 0.03408766, 0.02223298, 0.01084469, -0.003085196, 
    -0.01707561, -0.02659138, -0.0287623, -0.0287682, -0.03962229, 
    -0.06403226, -0.08689767, -0.1008428, -0.1162803, -0.1354081, -0.1528912, 
    -0.1690666, -0.1869894, -0.2025235, -0.2108463, -0.2093182, -0.2005226, 
    -0.1873806, -0.1713096, -0.1522519, -0.1306481, -0.1033428, -0.06294441, 
    -0.007835358, 0.04783711, 0.08105576, 0.09204787, 0.1008557, 0.1123894, 
    0.1221775, 0.132279, 0.1401801, 0.1459155, 0.1495649, 0.1497692, 
    0.1445933, 0.1336562, 0.1211396, 0.1102713, 0.09592907, 0.07591781, 
    0.05483071, 0.03392122, 0.009651888, -0.01987883, -0.03833022, 
    -0.04424148, -0.05192266, -0.06080569, -0.05692262, -0.02461319, 
    0.01884653, 0.05022803, 0.07262556, 0.09224725, 0.1106585, 0.1219989, 
    0.1203771, 0.1057023, 0.08023353, 0.04826903, 0.01694832, -0.005761263, 
    -0.01668184, -0.01628452, -0.003263148, 0.02100731, 0.05173182, 
    0.07975347, 0.09456486, 0.09285299, 0.07993655, 0.06016143, 0.03271666, 
    -0.001255482, -0.04200625, -0.08280234, -0.1189765, -0.1546835, 
    -0.1890008, -0.216198, -0.2349307, -0.2462892, -0.2467077, -0.2385679, 
    -0.2286008, -0.221873,
  -0.2084073, -0.2019022, -0.1864733, -0.1702564, -0.158909, -0.1429259, 
    -0.1241141, -0.1085566, -0.09252524, -0.07432523, -0.05684781, 
    -0.04334652, -0.0294435, -0.01130056, 0.007826507, 0.02396707, 
    0.03797205, 0.05078739, 0.0626398, 0.07308927, 0.08112827, 0.08763096, 
    0.09448621, 0.1007983, 0.1053069, 0.1093167, 0.1135165, 0.1176757, 
    0.1187675, 0.1154883, 0.1103738, 0.1061928, 0.1021586, 0.09635933, 
    0.08662263, 0.07113171, 0.0531005, 0.03981434, 0.03123583, 0.02430536, 
    0.01578617, 0.003049381, -0.009992391, -0.01328577, -0.01577711, 
    -0.04209751, -0.07829814, -0.1016728, -0.1222858, -0.1512577, -0.1821945, 
    -0.2120979, -0.2444949, -0.2771189, -0.3018061, -0.3147838, -0.3158665, 
    -0.3035993, -0.2789022, -0.245396, -0.2075407, -0.1704309, -0.1405565, 
    -0.1170723, -0.08678767, -0.03400642, 0.03661269, 0.090523, 0.1103796, 
    0.1164726, 0.124145, 0.1354182, 0.1477133, 0.1538001, 0.1548834, 
    0.1538144, 0.1510678, 0.1471011, 0.1362166, 0.114763, 0.08967045, 
    0.06381419, 0.03868639, 0.01734326, -0.001745943, -0.00891931, 
    0.0005173124, 0.01043228, 0.01967439, 0.03421875, 0.04058523, 0.03469378, 
    0.03002844, 0.04698657, 0.08371021, 0.1071425, 0.09289348, 0.04531957, 
    -0.01758778, -0.079414, -0.1278483, -0.1562285, -0.1668734, -0.1679108, 
    -0.1644067, -0.1578677, -0.1508933, -0.1408593, -0.1193507, -0.07713224, 
    -0.01734386, 0.03651814, 0.06102642, 0.05704939, 0.03780054, 0.006870896, 
    -0.03167403, -0.07157725, -0.1093628, -0.1478986, -0.1871979, -0.2114314, 
    -0.2276383, -0.2408003, -0.2424254, -0.2385156, -0.2282306, -0.2151701,
  -0.1951647, -0.1897573, -0.1808947, -0.1619485, -0.145234, -0.1338404, 
    -0.1201481, -0.1022255, -0.08302253, -0.0668726, -0.05310464, 
    -0.03897867, -0.02233756, -0.005195171, 0.01112902, 0.02713598, 
    0.04207503, 0.05477126, 0.06552632, 0.0743145, 0.08158048, 0.08873229, 
    0.0967813, 0.1043216, 0.110107, 0.1151943, 0.1195233, 0.1223122, 
    0.1220908, 0.1190854, 0.1154324, 0.1117389, 0.1066748, 0.1005546, 
    0.0925886, 0.07925187, 0.06169409, 0.04824801, 0.03877184, 0.02614351, 
    0.008997917, -0.01079302, -0.02946908, -0.03700507, -0.04349066, 
    -0.07442102, -0.1069921, -0.1236292, -0.1468454, -0.1813238, -0.2180108, 
    -0.26139, -0.3107261, -0.3570919, -0.3904494, -0.4093488, -0.4164295, 
    -0.4128355, -0.3958372, -0.3586723, -0.3019903, -0.2381036, -0.1801665, 
    -0.1371477, -0.1077814, -0.0813719, -0.03616875, 0.03621703, 0.09711412, 
    0.1239224, 0.131699, 0.1375764, 0.1449646, 0.15211, 0.1549657, 0.1552668, 
    0.1515536, 0.1397879, 0.1236388, 0.1074067, 0.08827861, 0.06924435, 
    0.05410009, 0.03840365, 0.02816508, 0.02468414, 0.01252321, -0.004034147, 
    0.0007403567, 0.02491806, 0.05369342, 0.09093627, 0.1261482, 0.1426282, 
    0.1164183, 0.03470998, -0.06443582, -0.1401156, -0.1803292, -0.1933726, 
    -0.192811, -0.1902986, -0.1884296, -0.1830769, -0.1717454, -0.1562134, 
    -0.1380063, -0.1246435, -0.1230611, -0.1284145, -0.1161545, -0.06773609, 
    -0.0046933, 0.02999707, 0.02919033, 0.007004127, -0.0293512, -0.06863515, 
    -0.103725, -0.1440372, -0.1827074, -0.2049828, -0.228629, -0.2398765, 
    -0.2331368, -0.2290566, -0.2244553, -0.20994,
  -0.1888077, -0.1773925, -0.1642338, -0.1483971, -0.1333468, -0.1197678, 
    -0.1050583, -0.08760712, -0.07075131, -0.05794838, -0.04481822, 
    -0.0289939, -0.01296146, 0.0005856454, 0.01390423, 0.03065104, 
    0.04803257, 0.05928882, 0.06601422, 0.07528596, 0.0869979, 0.09500577, 
    0.09813394, 0.1014739, 0.1082432, 0.1157302, 0.1195848, 0.1215561, 
    0.1238187, 0.1240804, 0.1206879, 0.1161159, 0.1124418, 0.1095722, 
    0.1034877, 0.09027166, 0.07140496, 0.0552516, 0.04310638, 0.02967612, 
    0.01666337, 0.005546115, -0.007353336, -0.01745477, -0.03233233, 
    -0.07138033, -0.1049427, -0.1216743, -0.1503924, -0.1959929, -0.251844, 
    -0.3130782, -0.3688543, -0.4114637, -0.4369455, -0.4528516, -0.4646377, 
    -0.4675022, -0.4610803, -0.4441816, -0.3991426, -0.3180457, -0.231051, 
    -0.1674719, -0.1262955, -0.09618771, -0.07099533, -0.02433914, 
    0.04742406, 0.1046139, 0.1323998, 0.1428267, 0.1490767, 0.1560053, 
    0.1619432, 0.1619985, 0.1569471, 0.1514715, 0.1420311, 0.1243144, 
    0.1046394, 0.08568725, 0.06400731, 0.04162743, 0.02111613, -0.002274632, 
    -0.02846309, -0.04207074, -0.03903766, -0.03119105, -0.009343237, 
    0.03837495, 0.07113391, 0.03497658, -0.06220765, -0.1522982, -0.1910305, 
    -0.197301, -0.205339, -0.2288506, -0.2588163, -0.2805145, -0.2875994, 
    -0.2826003, -0.2674445, -0.243994, -0.2157868, -0.1830007, -0.1491119, 
    -0.126554, -0.1207337, -0.111157, -0.07173448, -0.02032912, 0.005082458, 
    0.002122, -0.02203126, -0.06267418, -0.1053706, -0.1455586, -0.1702121, 
    -0.1975602, -0.2298958, -0.2369283, -0.2324246, -0.2225007, -0.2115709, 
    -0.2006969,
  -0.1764779, -0.1626674, -0.1433474, -0.1256955, -0.1148186, -0.1030451, 
    -0.08658871, -0.07032216, -0.05731773, -0.04516992, -0.0304749, 
    -0.01550578, -0.003834695, 0.007590909, 0.02456372, 0.04360137, 
    0.05492036, 0.05978274, 0.06888801, 0.08329683, 0.09229042, 0.09304059, 
    0.09623312, 0.1082958, 0.1202676, 0.1236806, 0.1221268, 0.1248993, 
    0.1317771, 0.1333009, 0.126827, 0.1209212, 0.1205469, 0.1201291, 
    0.1120994, 0.09661873, 0.08018719, 0.06741641, 0.0562509, 0.04125547, 
    0.02789326, 0.01782621, -0.002553836, -0.02569559, -0.03200815, 
    -0.05991966, -0.1041133, -0.124244, -0.1513489, -0.2068445, -0.2675492, 
    -0.3228627, -0.3735576, -0.4155614, -0.4526386, -0.4936583, -0.5321026, 
    -0.5495411, -0.5338237, -0.4954594, -0.4610789, -0.4016436, -0.2921833, 
    -0.1951363, -0.1431848, -0.1114394, -0.0810537, -0.05152887, 
    -0.005360588, 0.05933824, 0.1136276, 0.1419979, 0.1558098, 0.1645363, 
    0.1684005, 0.1668288, 0.1597812, 0.1478976, 0.1376325, 0.1277896, 
    0.1076197, 0.07982627, 0.05340652, 0.02811405, 0.00682037, -0.01395951, 
    -0.02673642, -0.02245053, -0.01604713, -0.02326087, -0.0125604, 
    0.03980847, 0.03327707, -0.05958916, -0.1492861, -0.1862858, -0.2074316, 
    -0.2479683, -0.2991309, -0.3396257, -0.3627875, -0.3766921, -0.3853701, 
    -0.3810144, -0.358687, -0.3249701, -0.288088, -0.2523551, -0.2160509, 
    -0.1772546, -0.1433309, -0.120477, -0.09689528, -0.05785151, -0.02686869, 
    -0.02203265, -0.03639383, -0.06941465, -0.1109062, -0.1396618, 
    -0.1667519, -0.2076674, -0.2235785, -0.2272805, -0.2311634, -0.2188439, 
    -0.2032081, -0.1886402,
  -0.1666536, -0.147284, -0.1301581, -0.115848, -0.1007761, -0.08471918, 
    -0.07167479, -0.05922875, -0.04462585, -0.02995354, -0.01726192, 
    -0.007131591, 0.00373828, 0.01844211, 0.03446657, 0.04690901, 0.05558923, 
    0.06553637, 0.0785312, 0.08889453, 0.09238166, 0.09527382, 0.1041629, 
    0.1145638, 0.117487, 0.1153385, 0.1191057, 0.1316425, 0.1409661, 
    0.1366469, 0.1269971, 0.1275688, 0.1345842, 0.1320136, 0.1189488, 
    0.1062454, 0.09773733, 0.08391489, 0.06411022, 0.0490161, 0.04341765, 
    0.03214966, 0.006338045, -0.02025759, -0.02864849, -0.04459259, 
    -0.08886868, -0.1203838, -0.1348818, -0.1810969, -0.2474818, -0.3079742, 
    -0.3636902, -0.4153959, -0.4566033, -0.5024674, -0.5571657, -0.5999866, 
    -0.6141865, -0.5804898, -0.507269, -0.4557214, -0.3661785, -0.2393695, 
    -0.161376, -0.1268229, -0.09969014, -0.05750459, -0.01382483, 0.03225922, 
    0.08011705, 0.1164763, 0.1389925, 0.1535581, 0.1580199, 0.1561226, 
    0.1560408, 0.1563931, 0.1477786, 0.1251105, 0.09937031, 0.07562946, 
    0.05569752, 0.04135575, 0.02279418, 0.003439173, 0.0006997511, 
    0.007404443, 0.004037827, 0.004030123, 0.01956835, 0.0422539, 
    -0.03104924, -0.1541331, -0.2152174, -0.2458162, -0.291153, -0.3349628, 
    -0.3698528, -0.4091267, -0.453086, -0.4928209, -0.5219897, -0.5351503, 
    -0.522368, -0.480517, -0.4222446, -0.3601859, -0.2988403, -0.2412306, 
    -0.1906358, -0.1474552, -0.1107401, -0.07904519, -0.05334024, 
    -0.04562866, -0.05376442, -0.07419902, -0.1034421, -0.1361251, 
    -0.1812293, -0.2140446, -0.2187953, -0.2287693, -0.2278195, -0.2083274, 
    -0.1943351, -0.1836621,
  -0.1515099, -0.1358744, -0.1207929, -0.1078133, -0.09225777, -0.07333651, 
    -0.05703053, -0.04439659, -0.03143805, -0.01667635, -0.003722988, 
    0.006494116, 0.01921652, 0.03509961, 0.04902879, 0.05861448, 0.06787582, 
    0.07931453, 0.08910763, 0.09337304, 0.09829911, 0.1081214, 0.1174942, 
    0.1203667, 0.1225722, 0.1311503, 0.1434043, 0.1482, 0.1444506, 0.1400665, 
    0.1444711, 0.1514555, 0.1490368, 0.1367738, 0.1304043, 0.1274226, 
    0.1168593, 0.09269038, 0.07484354, 0.0685028, 0.06151839, 0.04055962, 
    0.01803398, 0.001867414, -0.01114966, -0.03683122, -0.06855083, 
    -0.09902695, -0.114161, -0.1428439, -0.1996512, -0.2640404, -0.3154428, 
    -0.3686503, -0.418859, -0.4678422, -0.5147405, -0.5585127, -0.5797843, 
    -0.6014853, -0.5658978, -0.4863682, -0.4208698, -0.2937861, -0.1897036, 
    -0.1339459, -0.108226, -0.07691182, -0.02952185, 0.02419842, 0.06655645, 
    0.1010736, 0.1244782, 0.1412644, 0.1516541, 0.1679657, 0.1780965, 
    0.1672551, 0.1521933, 0.1375201, 0.1238108, 0.1056531, 0.08638382, 
    0.06090594, 0.03684916, 0.02148016, 0.01497652, 0.00468567, -0.004658047, 
    0.01015209, 0.05018137, 0.05273866, -0.07823944, -0.2005581, -0.2297529, 
    -0.268047, -0.3248231, -0.379388, -0.4401935, -0.4931786, -0.5262709, 
    -0.5535352, -0.5803047, -0.6032867, -0.6213613, -0.6168215, -0.5702572, 
    -0.4974322, -0.4190391, -0.3373879, -0.2580906, -0.192899, -0.1374505, 
    -0.09433706, -0.0740863, -0.06759164, -0.06288037, -0.0705139, 
    -0.1005882, -0.1465524, -0.1903871, -0.2096489, -0.214361, -0.2273507, 
    -0.2254994, -0.2003832, -0.1776044, -0.1650734,
  -0.1314632, -0.1199929, -0.1076291, -0.09658596, -0.08415014, -0.06931886, 
    -0.05295458, -0.03601485, -0.01896102, -0.002675362, 0.01291886, 
    0.02611616, 0.03914379, 0.05309196, 0.06729029, 0.07803643, 0.08890216, 
    0.1002471, 0.1110391, 0.1170673, 0.1227518, 0.1279245, 0.1341474, 
    0.1382405, 0.1441617, 0.1504597, 0.1570674, 0.1584204, 0.1621272, 
    0.1693366, 0.1773167, 0.1726225, 0.1635581, 0.1605928, 0.1677624, 
    0.1605521, 0.1359691, 0.1096543, 0.1066854, 0.1078395, 0.09374821, 
    0.06581052, 0.05510734, 0.05062297, 0.03077991, -0.007185608, 
    -0.02653015, -0.03519007, -0.05765311, -0.09055131, -0.1292152, 
    -0.1826718, -0.2468061, -0.305879, -0.3552409, -0.3972642, -0.4458007, 
    -0.4876195, -0.5061798, -0.5224226, -0.568156, -0.5102802, -0.4449209, 
    -0.3488151, -0.2311895, -0.1551072, -0.1077729, -0.07818375, -0.05300421, 
    -0.02017204, 0.02450325, 0.07016633, 0.1068147, 0.1292745, 0.1433753, 
    0.1616026, 0.172341, 0.1720694, 0.1654036, 0.1398944, 0.1320214, 
    0.120249, 0.0966984, 0.06695755, 0.04866692, 0.03312473, 0.01621562, 
    -0.001303945, 0.002866477, 0.03377778, 0.08104737, 0.03963942, 
    -0.1377427, -0.2252554, -0.2371152, -0.3075309, -0.3802994, -0.4323078, 
    -0.4782448, -0.5066585, -0.5259503, -0.5532215, -0.5806412, -0.6086447, 
    -0.6489888, -0.6891562, -0.7001779, -0.6518592, -0.5600545, -0.4665447, 
    -0.3608226, -0.2564147, -0.1791055, -0.1250311, -0.0885995, -0.08398473, 
    -0.0876535, -0.08926649, -0.1117304, -0.1554435, -0.1923182, -0.2048058, 
    -0.2055049, -0.2136675, -0.2085413, -0.1813664, -0.15705, -0.1427351,
  -0.1302558, -0.1310879, -0.1320901, -0.1338282, -0.1322946, -0.1251028, 
    -0.1110706, -0.09296491, -0.06925297, -0.04019058, -0.00844764, 
    0.01912492, 0.04330555, 0.06290866, 0.08032548, 0.09339166, 0.1038485, 
    0.1117345, 0.1221937, 0.130968, 0.1391095, 0.1446143, 0.1530175, 
    0.1593718, 0.1656129, 0.1697242, 0.1772414, 0.1827711, 0.1884407, 
    0.1881338, 0.1873754, 0.1848173, 0.1877844, 0.1882123, 0.1823272, 
    0.1617104, 0.1431157, 0.1342987, 0.1337203, 0.1206202, 0.09683581, 
    0.08258533, 0.07830647, 0.06960866, 0.04205893, 0.01542717, -0.005335391, 
    -0.007310048, -0.0274328, -0.05334194, -0.08600003, -0.1076154, 
    -0.153301, -0.2087378, -0.2729318, -0.323658, -0.3718872, -0.3995783, 
    -0.4389974, -0.4557583, -0.5310637, -0.5349498, -0.4620363, -0.4013551, 
    -0.300413, -0.2162039, -0.1522518, -0.1093504, -0.07348334, -0.04874197, 
    -0.02538757, -0.000425145, 0.0319127, 0.06586215, 0.1018968, 0.1293181, 
    0.1420698, 0.1484743, 0.1590957, 0.1470449, 0.1414465, 0.1209994, 
    0.1062162, 0.08155852, 0.05932887, 0.03891587, 0.02567242, 0.01285177, 
    0.01373113, 0.0460653, 0.08932665, 0.01650815, -0.1632603, -0.2052933, 
    -0.2363631, -0.3373887, -0.3844231, -0.4260492, -0.4812688, -0.4898622, 
    -0.4776128, -0.4895101, -0.4998924, -0.4996665, -0.5194065, -0.5836759, 
    -0.6649598, -0.7314055, -0.7037967, -0.6120253, -0.5122659, -0.3846568, 
    -0.2560174, -0.1750024, -0.1301525, -0.1009637, -0.09912243, -0.1088369, 
    -0.1237207, -0.1552836, -0.1855514, -0.1954466, -0.1943672, -0.1981247, 
    -0.1851136, -0.159247, -0.1441321, -0.1350267,
  -0.1636541, -0.1837759, -0.2019018, -0.2145235, -0.217531, -0.2136216, 
    -0.2033888, -0.1860099, -0.1590954, -0.1266097, -0.08997729, -0.05184833, 
    -0.01213975, 0.02457319, 0.05548947, 0.07793601, 0.09686291, 0.1114987, 
    0.1223161, 0.1288859, 0.1350392, 0.1409732, 0.1489997, 0.1562923, 
    0.1646443, 0.1726886, 0.1816597, 0.1886836, 0.1948909, 0.1988139, 
    0.2022773, 0.2032008, 0.2008263, 0.1933377, 0.184356, 0.1736487, 
    0.1614273, 0.1484376, 0.1378152, 0.1289333, 0.1192991, 0.1151279, 
    0.104098, 0.09797712, 0.06526947, 0.05684316, 0.03135969, 0.02978337, 
    0.008326575, 2.4423e-05, -0.02858049, -0.05149747, -0.08061777, 
    -0.1174634, -0.1787105, -0.2331991, -0.2801304, -0.3171314, -0.3621632, 
    -0.3912994, -0.4529493, -0.5175942, -0.4703249, -0.4332456, -0.3730499, 
    -0.3158696, -0.2621778, -0.2231096, -0.1852773, -0.153101, -0.1134543, 
    -0.07867339, -0.04103613, -0.009212457, 0.02310347, 0.05026937, 
    0.08941059, 0.1286807, 0.1535022, 0.1433467, 0.1548831, 0.1492069, 
    0.1381388, 0.1165336, 0.08676251, 0.06178448, 0.05162175, 0.0388035, 
    0.02096887, 0.05104922, 0.100075, 0.007444285, -0.167364, -0.1984266, 
    -0.2608088, -0.3485764, -0.3698565, -0.4282403, -0.4467107, -0.4191996, 
    -0.4321843, -0.4526916, -0.4376868, -0.4176791, -0.4199341, -0.4606881, 
    -0.5396113, -0.6484266, -0.7556593, -0.7415068, -0.6497903, -0.5464257, 
    -0.404094, -0.2620402, -0.1798196, -0.1441797, -0.1205735, -0.1184551, 
    -0.1300538, -0.1500442, -0.1663198, -0.1713624, -0.1789986, -0.1836046, 
    -0.1628284, -0.1377648, -0.1345804, -0.1472923,
  -0.2018697, -0.2298556, -0.2423573, -0.2458038, -0.2425872, -0.2342113, 
    -0.223989, -0.2142095, -0.2014932, -0.1804303, -0.1529701, -0.123657, 
    -0.0914022, -0.05793405, -0.02746096, -0.00212489, 0.01716812, 
    0.03435741, 0.04914998, 0.06081205, 0.07081389, 0.08365931, 0.09794024, 
    0.1118466, 0.1250828, 0.1403687, 0.1535246, 0.1644743, 0.1727154, 
    0.1810285, 0.1836693, 0.183335, 0.1811108, 0.1794741, 0.1691613, 
    0.1547907, 0.140523, 0.1360203, 0.1305876, 0.1227223, 0.1111042, 
    0.1053984, 0.09521826, 0.08520848, 0.06167509, 0.05931082, 0.02673078, 
    0.03796966, 0.007265776, 0.005379081, -0.0004346669, -0.007430747, 
    -0.02461587, -0.05863172, -0.1006699, -0.1493024, -0.1913765, -0.2331924, 
    -0.2801861, -0.3224532, -0.3593597, -0.4738726, -0.4636953, -0.4482131, 
    -0.426082, -0.4079402, -0.3922083, -0.3845891, -0.378083, -0.3687801, 
    -0.3491053, -0.3167867, -0.2665616, -0.2050472, -0.1331477, -0.06684092, 
    -0.01265159, 0.0216105, 0.06499883, 0.112675, 0.1505426, 0.1426031, 
    0.1410263, 0.1354836, 0.1192154, 0.1027028, 0.08517924, 0.07227242, 
    0.04743334, 0.05935604, 0.104713, 0.02767738, -0.1359845, -0.1730385, 
    -0.2436061, -0.3135885, -0.3394114, -0.3880469, -0.3952924, -0.4104849, 
    -0.4194174, -0.3983158, -0.3805541, -0.3582434, -0.3490891, -0.3555385, 
    -0.4015343, -0.4590111, -0.6007655, -0.7652498, -0.7718127, -0.6890128, 
    -0.5772762, -0.4247402, -0.2767123, -0.1922586, -0.157246, -0.1360842, 
    -0.1279701, -0.1347138, -0.1437132, -0.1560442, -0.1692746, -0.1682701, 
    -0.1455256, -0.1270418, -0.1322886, -0.1627779,
  -0.2284679, -0.2375185, -0.2309563, -0.2220865, -0.2143489, -0.2042426, 
    -0.190781, -0.1755208, -0.1646323, -0.158152, -0.1465739, -0.1307258, 
    -0.1176221, -0.1007023, -0.08517732, -0.07196763, -0.06199034, 
    -0.05374342, -0.04807272, -0.04175469, -0.03500946, -0.02271493, 
    -0.003526777, 0.02403771, 0.0532632, 0.08280797, 0.1085987, 0.1303309, 
    0.142818, 0.1527683, 0.1591185, 0.1621224, 0.1559013, 0.1487347, 
    0.1392752, 0.13041, 0.1168725, 0.105994, 0.09528275, 0.09176251, 
    0.08488826, 0.07895607, 0.07071729, 0.06752512, 0.05659527, 0.04280906, 
    0.02851146, 0.03130302, 0.004539937, 0.03343084, 0.01909463, 0.004266575, 
    -0.008962914, -0.03966917, -0.06058224, -0.08953495, -0.1091811, 
    -0.1543538, -0.2074503, -0.2602805, -0.2951173, -0.4437349, -0.4526519, 
    -0.4370678, -0.4536863, -0.4765053, -0.5167754, -0.5578218, -0.6065833, 
    -0.6430429, -0.6526209, -0.6323992, -0.5824111, -0.5113745, -0.4245569, 
    -0.3288917, -0.2195288, -0.1125499, -0.03476828, 0.01154018, 0.07137159, 
    0.1175878, 0.137273, 0.13632, 0.1329664, 0.1307073, 0.1221752, 0.1159603, 
    0.09023563, 0.0846328, 0.1243109, 0.08207726, -0.08617114, -0.1501534, 
    -0.2152014, -0.2800309, -0.3113528, -0.3450967, -0.3675871, -0.3648188, 
    -0.3416905, -0.3260324, -0.2951619, -0.2770864, -0.2809519, -0.2647376, 
    -0.2656009, -0.3060072, -0.3805548, -0.5647231, -0.757228, -0.7927096, 
    -0.7232991, -0.6076214, -0.4487896, -0.3022345, -0.2107655, -0.1687596, 
    -0.1382715, -0.1203819, -0.1173605, -0.1288941, -0.1430316, -0.1300765, 
    -0.113792, -0.1202511, -0.151095, -0.196245,
  -0.200654, -0.2008953, -0.1973935, -0.1971764, -0.1991892, -0.1957651, 
    -0.1845242, -0.1646227, -0.1379272, -0.1148351, -0.1043963, -0.09463601, 
    -0.09108698, -0.0873719, -0.07998997, -0.07603079, -0.07733769, 
    -0.07654144, -0.0723855, -0.06656095, -0.06288688, -0.05740685, 
    -0.05037998, -0.03955658, -0.02067286, 0.005420048, 0.02915571, 
    0.05180741, 0.06588231, 0.06952016, 0.06388193, 0.05824313, 0.04855943, 
    0.03058184, 0.005329985, -0.01344562, -0.02897465, -0.04472003, 
    -0.05952213, -0.06637862, -0.07665077, -0.08447485, -0.08484667, 
    -0.08222815, -0.09617153, -0.1050181, -0.1091363, -0.1216622, -0.1151223, 
    -0.07404597, -0.07389113, -0.04125765, -0.02640936, -0.03396077, 
    -0.03087777, -0.06224268, -0.07926843, -0.1216747, -0.1509525, 
    -0.1886371, -0.2109164, -0.3504729, -0.3963487, -0.3941455, -0.455613, 
    -0.5221629, -0.6409408, -0.7981746, -0.9616665, -1.092248, -1.173363, 
    -1.187919, -1.138426, -1.025957, -0.8658704, -0.6856294, -0.5222861, 
    -0.3809161, -0.2327724, -0.09413113, -0.01692094, 0.0332735, 0.1119162, 
    0.1575556, 0.1574869, 0.1557846, 0.1568264, 0.1572791, 0.1436524, 
    0.1317058, 0.1478637, 0.1472608, 0.00387525, -0.09520637, -0.147783, 
    -0.2132531, -0.2532806, -0.2761588, -0.3091134, -0.3289068, -0.3167232, 
    -0.2792358, -0.2548828, -0.2532173, -0.2288118, -0.2010959, -0.1670736, 
    -0.1799895, -0.235496, -0.3452985, -0.5493665, -0.7525045, -0.8115889, 
    -0.7584665, -0.6374682, -0.4740694, -0.3298735, -0.234619, -0.1810737, 
    -0.1356739, -0.1025963, -0.1032773, -0.1134272, -0.08937042, -0.07268886, 
    -0.09613758, -0.1398896, -0.1815283,
  -0.1673931, -0.1762511, -0.1838241, -0.1820529, -0.1774822, -0.176234, 
    -0.1691341, -0.1497672, -0.1176174, -0.07924534, -0.05778695, 
    -0.04942564, -0.04766987, -0.05341694, -0.05928918, -0.06613375, 
    -0.07502665, -0.07990813, -0.07783958, -0.07283695, -0.06958957, 
    -0.06192221, -0.03919275, -0.01639897, -0.01488842, -0.0181004, 
    -0.01926079, -0.02032068, -0.02657835, -0.03995059, -0.05353592, 
    -0.06479114, -0.08283005, -0.104192, -0.1151415, -0.1212343, -0.1405068, 
    -0.1606308, -0.1613232, -0.1559122, -0.1639276, -0.1662761, -0.1573913, 
    -0.1596734, -0.1729387, -0.1714413, -0.1716245, -0.1849852, -0.17537, 
    -0.1525484, -0.1648803, -0.163338, -0.1643668, -0.1473199, -0.09793689, 
    -0.09250408, -0.07920782, -0.1180327, -0.1285896, -0.1487332, -0.1582943, 
    -0.2616727, -0.3722009, -0.3792224, -0.4313969, -0.5583402, -0.7899458, 
    -1.05646, -1.304395, -1.465533, -1.543468, -1.578846, -1.591093, 
    -1.567717, -1.481594, -1.297801, -1.01882, -0.7179338, -0.4942366, 
    -0.3229047, -0.1360565, -0.006761547, 0.05170687, 0.1377259, 0.1918206, 
    0.1997884, 0.197637, 0.1989314, 0.1908196, 0.1880165, 0.2030586, 
    0.2180656, 0.1119822, -0.02912699, -0.08471974, -0.1427592, -0.1927402, 
    -0.2132094, -0.2437281, -0.2674789, -0.2482076, -0.240999, -0.218232, 
    -0.2013501, -0.1860787, -0.16666, -0.1256292, -0.09961822, -0.1088041, 
    -0.1868449, -0.319032, -0.5187892, -0.7410415, -0.8178334, -0.7898332, 
    -0.6702126, -0.4984112, -0.3480774, -0.246526, -0.1808891, -0.1189249, 
    -0.07657828, -0.08439013, -0.0643459, -0.03791657, -0.06644686, 
    -0.1218315, -0.157204,
  -0.122133, -0.1277565, -0.1331153, -0.1394206, -0.1461949, -0.1447923, 
    -0.1269988, -0.1075986, -0.08458558, -0.04760791, -0.01867968, 
    -0.01086207, -0.01486626, -0.0249138, -0.03951123, -0.05426657, 
    -0.06416246, -0.06231597, -0.0540515, -0.05167572, -0.060165, 
    -0.06405374, -0.04496851, 0.008618444, 0.04278034, 0.03620335, 
    0.02246262, 0.003990412, -0.02567677, -0.05899792, -0.08005516, 
    -0.1004383, -0.1308931, -0.158415, -0.1759793, -0.2037514, -0.2383056, 
    -0.2532467, -0.2547925, -0.2715264, -0.2901035, -0.2905798, -0.2898095, 
    -0.2997109, -0.2963485, -0.276298, -0.269006, -0.2747251, -0.246204, 
    -0.2015413, -0.1727426, -0.1444677, -0.1486099, -0.2041434, -0.2110285, 
    -0.2003519, -0.1440701, -0.1568967, -0.1632299, -0.1477334, -0.1353955, 
    -0.1705011, -0.2912773, -0.2941051, -0.3531762, -0.5427349, -0.8228166, 
    -1.157604, -1.398711, -1.471785, -1.492187, -1.511861, -1.537015, 
    -1.564763, -1.599365, -1.613682, -1.546647, -1.30505, -0.9057701, 
    -0.5524248, -0.3500167, -0.1434204, 0.03103282, 0.1006805, 0.1787755, 
    0.2438904, 0.2523692, 0.2455255, 0.2400364, 0.2426399, 0.257158, 
    0.2853492, 0.2341885, 0.08543295, 0.002850578, -0.04082213, -0.1014868, 
    -0.127033, -0.1434327, -0.1751641, -0.192469, -0.1809329, -0.1355322, 
    -0.1331996, -0.1346768, -0.1214374, -0.1033518, -0.0706567, -0.02891727, 
    -0.02771416, -0.1376694, -0.2623179, -0.48575, -0.7043719, -0.7967429, 
    -0.8030531, -0.6869043, -0.5033206, -0.3461596, -0.2328691, -0.1459078, 
    -0.06183717, -0.02647375, -0.03341142, -0.01080382, -0.02784193, 
    -0.07895714, -0.112574,
  -0.06376509, -0.08347515, -0.09179099, -0.09857422, -0.1061951, 
    -0.09636842, -0.07267427, -0.05572825, -0.04597919, -0.03367009, 
    -0.02065969, -0.01273274, -0.01426019, -0.02063892, -0.0265194, 
    -0.02456328, -0.01814511, -0.0003342722, 0.0158915, 0.01500142, 
    0.0006597564, 0.007462053, 0.01624308, 0.03758566, 0.07197356, 
    0.05735909, 0.02161635, -0.02211624, -0.08075237, -0.1378315, -0.1761738, 
    -0.2156083, -0.2664465, -0.31349, -0.3465206, -0.3819237, -0.4204327, 
    -0.4418941, -0.4397698, -0.4423802, -0.4589683, -0.4728113, -0.4789127, 
    -0.4906689, -0.4982316, -0.4913323, -0.4812636, -0.4782599, -0.4550142, 
    -0.4156387, -0.3690794, -0.2952342, -0.1932136, -0.1574638, -0.1643084, 
    -0.1772801, -0.1702708, -0.1604862, -0.2048488, -0.1977261, -0.170077, 
    -0.1063599, -0.1816337, -0.2235828, -0.2444111, -0.4160134, -0.7090861, 
    -1.090286, -1.305813, -1.349184, -1.348099, -1.39512, -1.43258, 
    -1.471463, -1.503839, -1.520464, -1.545012, -1.558137, -1.423299, 
    -1.010603, -0.5465474, -0.3066433, -0.09759925, 0.09857523, 0.1647941, 
    0.2365103, 0.3004377, 0.3104571, 0.2976207, 0.3039933, 0.3292413, 
    0.3616506, 0.341959, 0.2100183, 0.09124756, 0.0525552, -0.00620088, 
    -0.04612058, -0.04679624, -0.05941696, -0.08190925, -0.08705217, 
    -0.07437611, -0.05610679, -0.06259608, -0.0632277, -0.05810263, 
    -0.02990179, 0.01471944, 0.05663262, 0.008769495, -0.08518068, 
    -0.2269091, -0.4769869, -0.6783242, -0.7954189, -0.8017459, -0.6668855, 
    -0.4669182, -0.3087506, -0.1803885, -0.06630038, 0.0261661, 0.03939748, 
    0.03660772, 0.02719507, -0.01789818, -0.0433673,
  -0.007216893, -0.01532783, -0.01765077, -0.03876241, -0.0459162, 
    -0.03096741, -0.02026644, -0.02547713, -0.03045344, -0.03023308, 
    -0.02980798, -0.02857459, -0.01835241, -0.001870915, 0.00992186, 
    0.02003927, 0.03558639, 0.06593192, 0.074036, 0.04393548, 0.02120129, 
    0.06185643, 0.0966151, 0.08573414, 0.08223815, 0.0460067, -0.01283552, 
    -0.08254349, -0.1595215, -0.229278, -0.2801256, -0.3178607, -0.3534632, 
    -0.3952676, -0.4378162, -0.475841, -0.5131304, -0.5549764, -0.5860157, 
    -0.5971274, -0.6017287, -0.6091239, -0.6182083, -0.6335274, -0.6547733, 
    -0.6619141, -0.6484624, -0.6340717, -0.6259055, -0.6062666, -0.5671793, 
    -0.504394, -0.4143186, -0.3036648, -0.2166676, -0.1604873, -0.1411322, 
    -0.09372634, -0.1048569, -0.1661472, -0.1961063, -0.1315221, -0.09215833, 
    -0.1504182, -0.1286654, -0.2210427, -0.4818964, -0.8570667, -1.138339, 
    -1.213211, -1.202386, -1.250914, -1.297867, -1.313592, -1.381917, 
    -1.443168, -1.48195, -1.486494, -1.490727, -1.402577, -0.9962894, 
    -0.4697133, -0.2132176, -0.0002946397, 0.1953575, 0.2492032, 0.2999869, 
    0.3502798, 0.3759364, 0.3819711, 0.3917237, 0.4267111, 0.4487172, 
    0.3554336, 0.2165991, 0.1632077, 0.1190887, 0.06635954, 0.05819402, 
    0.04774998, 0.02160903, 0.01054851, 0.009051632, 0.009518575, 0.01486699, 
    -0.003686899, -0.04106514, -0.003549566, 0.07976817, 0.110347, 0.1016474, 
    0.0357134, -0.07311536, -0.2443274, -0.4778327, -0.6733135, -0.7905605, 
    -0.7686899, -0.5897405, -0.3776285, -0.2161372, -0.07680309, 0.05259033, 
    0.1191034, 0.1242082, 0.1154499, 0.07230398, 0.02581513,
  0.08039972, 0.07174958, 0.0520245, 0.01782018, 0.006340824, 0.003901541, 
    -0.001722142, -0.0121245, -0.02094115, -0.0193842, -0.006892003, 
    0.005954243, 0.01838101, 0.03368631, 0.05156405, 0.07173893, 0.09424596, 
    0.1075932, 0.08991987, 0.0691091, 0.0824647, 0.1451048, 0.1816351, 
    0.146187, 0.08238675, -0.0001710504, -0.07723237, -0.1484579, -0.2199684, 
    -0.2893768, -0.3472746, -0.3913642, -0.4253594, -0.4542903, -0.4815733, 
    -0.5135064, -0.5504378, -0.587914, -0.6244243, -0.6591359, -0.6892754, 
    -0.704852, -0.7066891, -0.7049712, -0.7185229, -0.7423508, -0.7553418, 
    -0.7422593, -0.7261715, -0.7293337, -0.7223057, -0.6618834, -0.5567073, 
    -0.4490483, -0.3326553, -0.2115322, -0.1410428, -0.08829687, 
    -0.005095161, -0.008169591, -0.08528384, -0.135944, -0.06524631, 
    -0.05383094, -0.06289481, -0.03332898, -0.1935628, -0.5157772, 
    -0.8545886, -1.041772, -1.064565, -1.070543, -1.117567, -1.122206, 
    -1.154451, -1.258578, -1.3429, -1.402646, -1.426573, -1.408561, 
    -1.306637, -0.8711427, -0.3296187, -0.08597246, 0.130991, 0.310736, 
    0.3422655, 0.3757397, 0.4136807, 0.4597619, 0.4873325, 0.5044378, 
    0.5356631, 0.4800074, 0.3426099, 0.2642544, 0.2299565, 0.1784085, 
    0.1579196, 0.1552967, 0.1432972, 0.1247674, 0.09761849, 0.0971682, 
    0.106538, 0.0974452, 0.03347812, 0.04071192, 0.1434406, 0.1795568, 
    0.154812, 0.09143317, 0.01870283, -0.06547554, -0.2616764, -0.4770378, 
    -0.6708902, -0.765672, -0.6633269, -0.4447838, -0.2289911, -0.06792901, 
    0.07424277, 0.1758048, 0.2102484, 0.198311, 0.1533068, 0.1099972,
  0.1725229, 0.1479565, 0.1252837, 0.09667714, 0.07489812, 0.04223048, 
    0.01896066, 0.008410983, 0.00151898, 0.001130328, 0.009351179, 
    0.01795663, 0.02650485, 0.04055557, 0.06728689, 0.09875138, 0.1158596, 
    0.1068288, 0.1054186, 0.1332363, 0.168382, 0.2038745, 0.1937806, 
    0.1288691, 0.04507267, -0.03617455, -0.1047551, -0.1693868, -0.2347505, 
    -0.2955709, -0.3440782, -0.3869522, -0.4358917, -0.4903184, -0.5354384, 
    -0.5708847, -0.6097602, -0.6461039, -0.6661786, -0.6721986, -0.6935689, 
    -0.7282388, -0.7516584, -0.7448606, -0.7244351, -0.7260375, -0.7401071, 
    -0.7494248, -0.7372608, -0.7305789, -0.73543, -0.7214847, -0.6445991, 
    -0.524236, -0.4201034, -0.2970601, -0.1616177, -0.1075336, -0.0428694, 
    0.04157835, 0.06300958, -0.0124041, -0.05977619, -0.002546765, 
    0.008465819, 0.05088722, 0.06077515, -0.1385561, -0.4443417, -0.7383196, 
    -0.8893616, -0.9155857, -0.926974, -0.9624279, -0.9969624, -1.107853, 
    -1.216172, -1.268676, -1.325582, -1.340958, -1.310906, -1.165807, 
    -0.6769312, -0.1547071, 0.05948345, 0.2791657, 0.4341032, 0.4672151, 
    0.4979714, 0.5477192, 0.5864216, 0.5995914, 0.6230564, 0.5954713, 
    0.4931895, 0.3998935, 0.3548441, 0.3027653, 0.276909, 0.2636153, 
    0.2464218, 0.2319199, 0.2200052, 0.1897394, 0.177998, 0.1666026, 
    0.145562, 0.1902222, 0.2144923, 0.1904743, 0.1536585, 0.1092298, 
    0.06786971, 0.00424777, -0.1374027, -0.2992449, -0.5079855, -0.6855469, 
    -0.6618856, -0.4690816, -0.2353788, -0.03175189, 0.1182162, 0.2260619, 
    0.2842739, 0.2833152, 0.2535557, 0.2172806,
  0.2684249, 0.2515041, 0.2184716, 0.1720217, 0.1399333, 0.09123859, 
    0.06080502, 0.05667286, 0.04086446, 0.02068038, 0.01256979, 0.01787845, 
    0.03203835, 0.05437754, 0.08635862, 0.1161535, 0.1286573, 0.1424239, 
    0.1812378, 0.2126225, 0.2205893, 0.2109309, 0.1676311, 0.1047562, 
    0.03030073, -0.05221896, -0.1353487, -0.2106562, -0.2789799, -0.3385982, 
    -0.3849192, -0.414308, -0.4362355, -0.4690499, -0.5144911, -0.564737, 
    -0.6223693, -0.6807979, -0.7345678, -0.7584665, -0.7533792, -0.7434386, 
    -0.747413, -0.7658542, -0.7667713, -0.7471535, -0.7226162, -0.7035376, 
    -0.6992577, -0.7093565, -0.7113012, -0.6740659, -0.6228085, -0.5365232, 
    -0.4218448, -0.3350879, -0.2163069, -0.1225326, -0.0618775, 0.01917584, 
    0.1074938, 0.1357393, 0.04956415, 0.0172667, 0.05933603, 0.09992363, 
    0.1770265, 0.1554868, -0.02868411, -0.2987023, -0.5676802, -0.7239491, 
    -0.7697172, -0.7677, -0.7828585, -0.8464949, -1.004861, -1.147651, 
    -1.206822, -1.2389, -1.231457, -1.183906, -0.9914039, -0.4549569, 
    0.022264, 0.2080476, 0.4145143, 0.5619047, 0.6113287, 0.6627156, 
    0.7004776, 0.7106972, 0.7084339, 0.6849977, 0.6112685, 0.5276367, 
    0.4719648, 0.4202956, 0.3856265, 0.3775674, 0.3729418, 0.360648, 
    0.3302296, 0.3001634, 0.2556709, 0.2252008, 0.2742264, 0.2765487, 
    0.2111431, 0.1502153, 0.1042937, 0.06656015, 0.03847602, 0.003115878, 
    -0.08234412, -0.213071, -0.3999089, -0.5741605, -0.6087509, -0.441784, 
    -0.1990914, 0.01744082, 0.1888513, 0.2844748, 0.3609519, 0.3718814, 
    0.3510263, 0.3196179,
  0.3795265, 0.3725083, 0.3094023, 0.2496298, 0.2234942, 0.1706749, 
    0.1329518, 0.1143229, 0.08384241, 0.05910587, 0.03991253, 0.04492022, 
    0.07457321, 0.1082027, 0.1373018, 0.1698347, 0.2056796, 0.2410546, 
    0.2552381, 0.2423248, 0.2169252, 0.174275, 0.1095693, 0.03120501, 
    -0.05415704, -0.1409308, -0.2235603, -0.2953433, -0.3552904, -0.4087854, 
    -0.4612063, -0.505911, -0.5336438, -0.5560468, -0.581223, -0.609784, 
    -0.6367961, -0.6560448, -0.6919507, -0.7423037, -0.7882662, -0.7941356, 
    -0.7613024, -0.7197263, -0.706077, -0.7097906, -0.7090552, -0.673564, 
    -0.6243845, -0.6142826, -0.665423, -0.6246672, -0.544275, -0.5173645, 
    -0.4467328, -0.3395444, -0.2360458, -0.1290983, -0.03494367, 0.04668204, 
    0.1283361, 0.2127445, 0.1596452, 0.06828185, 0.07725818, 0.1219261, 
    0.2084694, 0.2987659, 0.266411, 0.1154315, -0.1273706, -0.3787364, 
    -0.5515958, -0.6191322, -0.6285702, -0.660136, -0.74705, -0.9168556, 
    -1.048648, -1.129649, -1.144562, -1.111473, -1.038613, -0.8028693, 
    -0.2531366, 0.1809032, 0.3461125, 0.5210782, 0.6725006, 0.7376926, 
    0.7762372, 0.8020642, 0.8045182, 0.7814348, 0.7242806, 0.6645846, 
    0.6053536, 0.5512601, 0.5057598, 0.4907985, 0.4778471, 0.4666892, 
    0.4333102, 0.389282, 0.3414153, 0.3408403, 0.3143616, 0.2363769, 
    0.1617395, 0.07723923, 0.01249197, -0.01060458, -0.01868536, -0.05977356, 
    -0.150673, -0.2470532, -0.3524627, -0.4946776, -0.5161461, -0.3702163, 
    -0.1249404, 0.08796338, 0.278368, 0.3732816, 0.4454486, 0.4858027, 
    0.4600572, 0.42087,
  0.4942888, 0.4775218, 0.4047205, 0.345324, 0.3113062, 0.251014, 0.2170477, 
    0.1863666, 0.1344575, 0.103784, 0.09221441, 0.1048147, 0.1405077, 
    0.1866713, 0.2210363, 0.239752, 0.2564712, 0.2638605, 0.24551, 0.2056919, 
    0.1512015, 0.08373607, 0.003513873, -0.08541029, -0.1723827, -0.2503516, 
    -0.3164128, -0.3744193, -0.4223382, -0.4594466, -0.4920159, -0.533015, 
    -0.5764021, -0.6191379, -0.6507511, -0.68348, -0.7157903, -0.7267668, 
    -0.7167274, -0.6960481, -0.6970927, -0.7311072, -0.7509521, -0.708238, 
    -0.6372916, -0.610428, -0.6425859, -0.633294, -0.567057, -0.5212827, 
    -0.58582, -0.5531639, -0.4586037, -0.4479281, -0.4442406, -0.3762596, 
    -0.2633305, -0.1367102, -0.02383752, 0.06662238, 0.1345886, 0.2190507, 
    0.2210613, 0.1340609, 0.098409, 0.1127551, 0.1917471, 0.3262758, 
    0.4003382, 0.3687521, 0.2480058, 0.03066902, -0.2016263, -0.3862934, 
    -0.4560908, -0.4961264, -0.5813477, -0.762286, -0.9230132, -0.9890231, 
    -1.015099, -1.029253, -0.9782757, -0.8847454, -0.6371903, -0.115103, 
    0.3049231, 0.4660893, 0.5882511, 0.7211243, 0.8088246, 0.8477861, 
    0.8539719, 0.829394, 0.7900983, 0.7489033, 0.7074395, 0.6570482, 
    0.6040007, 0.5943335, 0.6072063, 0.5713677, 0.4912457, 0.4710793, 
    0.4627199, 0.370434, 0.2541728, 0.1706519, 0.07940105, -0.01548516, 
    -0.0927653, -0.1328076, -0.1219708, -0.1039021, -0.1347209, -0.2094845, 
    -0.3164079, -0.4377171, -0.421418, -0.267189, -0.02369098, 0.182551, 
    0.3693969, 0.4910387, 0.5481901, 0.5947217, 0.5728192, 0.5244951,
  0.6047856, 0.574514, 0.5192019, 0.4564781, 0.400991, 0.3424577, 0.3182818, 
    0.2709283, 0.1964742, 0.1637359, 0.1630355, 0.1791933, 0.2008755, 
    0.232731, 0.2548297, 0.2561218, 0.2445633, 0.2206796, 0.1767491, 
    0.1053997, 0.01325813, -0.08631703, -0.1825164, -0.2730356, -0.3534071, 
    -0.4153313, -0.4562553, -0.4869225, -0.5128206, -0.533762, -0.5501341, 
    -0.5710493, -0.599337, -0.6342238, -0.6478432, -0.6554679, -0.6747126, 
    -0.7061844, -0.7175295, -0.6974204, -0.6505727, -0.6168231, -0.6229637, 
    -0.6164216, -0.5688667, -0.5205256, -0.5360605, -0.5447085, -0.5015342, 
    -0.4461492, -0.4662087, -0.4329825, -0.4019012, -0.401968, -0.3790129, 
    -0.3331926, -0.2543388, -0.1279336, -0.005290568, 0.07537106, 0.1471853, 
    0.2123253, 0.265384, 0.2171575, 0.1369158, 0.09932521, 0.1197259, 
    0.2288066, 0.3964059, 0.4941508, 0.4874742, 0.3494895, 0.1507722, 
    -0.08667607, -0.2545402, -0.3326117, -0.418529, -0.5849811, -0.7844777, 
    -0.8771383, -0.9120039, -0.9155276, -0.9130225, -0.8398846, -0.7376224, 
    -0.5205274, -0.07161041, 0.3571362, 0.5625219, 0.6472026, 0.7161336, 
    0.7827849, 0.8288886, 0.8478751, 0.837166, 0.8101181, 0.7755332, 
    0.7374372, 0.7085094, 0.6914204, 0.6571069, 0.6104877, 0.5904392, 
    0.5460264, 0.4111825, 0.2760541, 0.1828622, 0.08473295, -0.007667396, 
    -0.07979946, -0.1349839, -0.177095, -0.1877611, -0.1681716, -0.1442319, 
    -0.1657984, -0.2550229, -0.3529671, -0.328867, -0.1655061, 0.08405682, 
    0.2970304, 0.4650741, 0.5937457, 0.6586537, 0.6956729, 0.6852914, 
    0.6391954,
  0.7087302, 0.6776686, 0.6321465, 0.5577645, 0.5017943, 0.4495794, 
    0.3982583, 0.3623801, 0.2947348, 0.2351938, 0.2262919, 0.2400961, 
    0.2366577, 0.2377413, 0.2326918, 0.2068669, 0.1610542, 0.09304379, 
    0.004797202, -0.09361089, -0.1932184, -0.284381, -0.3613051, -0.4216985, 
    -0.466052, -0.4951988, -0.5110267, -0.5191654, -0.5300663, -0.5447376, 
    -0.5658261, -0.5892903, -0.611255, -0.6342216, -0.6396162, -0.6259903, 
    -0.6069834, -0.6090741, -0.6254954, -0.6149187, -0.5719646, -0.5172188, 
    -0.5064365, -0.5113929, -0.4783615, -0.4348518, -0.4369833, -0.4446033, 
    -0.4104037, -0.352437, -0.3422485, -0.3305433, -0.3297736, -0.3158261, 
    -0.2965266, -0.2687251, -0.213213, -0.1344763, 0.004626639, 0.08663492, 
    0.1432287, 0.1909259, 0.2474076, 0.2633719, 0.2115827, 0.1292327, 
    0.06125937, 0.07218999, 0.1851788, 0.3797914, 0.5686684, 0.5560832, 
    0.4193441, 0.2007899, -0.03270525, -0.1637374, -0.2815852, -0.4670934, 
    -0.6360438, -0.7166893, -0.7939043, -0.8110913, -0.8079034, -0.7918887, 
    -0.7119182, -0.6101038, -0.4547456, -0.1291259, 0.268672, 0.5562904, 
    0.6981652, 0.7604461, 0.7910571, 0.8076636, 0.8101771, 0.8035437, 
    0.7908493, 0.7831038, 0.7690032, 0.7397417, 0.7021152, 0.6575462, 
    0.5557367, 0.395725, 0.2648131, 0.1845157, 0.09599825, 0.002596524, 
    -0.07604137, -0.1266141, -0.1482778, -0.1604287, -0.1671637, -0.158814, 
    -0.131477, -0.1277835, -0.1879145, -0.2576156, -0.2333351, -0.08248022, 
    0.1784941, 0.4002589, 0.5593977, 0.6864172, 0.759262, 0.7850975, 
    0.7785133, 0.7444633,
  0.8039651, 0.7770206, 0.7352042, 0.6613106, 0.6067711, 0.5516341, 
    0.4936883, 0.4779044, 0.4018019, 0.3271542, 0.3096097, 0.3126835, 
    0.2834678, 0.2405158, 0.1956212, 0.1287474, 0.04067475, -0.05502385, 
    -0.1454349, -0.227294, -0.3020844, -0.3688035, -0.4253879, -0.4686845, 
    -0.5007582, -0.5166158, -0.5142355, -0.502486, -0.5046031, -0.5246513, 
    -0.5507175, -0.5615603, -0.5644653, -0.5708019, -0.5765028, -0.5644805, 
    -0.5402804, -0.5179336, -0.5131746, -0.5022909, -0.4496635, -0.3922111, 
    -0.3859629, -0.4023502, -0.3784795, -0.3395695, -0.3249224, -0.3236642, 
    -0.2840162, -0.2305726, -0.2432631, -0.2711183, -0.2399741, -0.217519, 
    -0.2330974, -0.2334798, -0.1728216, -0.1424361, -0.07545713, 0.03926715, 
    0.1320431, 0.1837188, 0.2265139, 0.27471, 0.2760285, 0.221638, 0.1568992, 
    0.07879192, 0.04813819, 0.126795, 0.3679316, 0.6081903, 0.6107607, 
    0.4180119, 0.1553558, -0.007251449, -0.1469315, -0.344265, -0.5062271, 
    -0.5905346, -0.649864, -0.6878772, -0.6982259, -0.6915766, -0.67145, 
    -0.6008407, -0.5042525, -0.4016703, -0.2261832, 0.03879444, 0.3136641, 
    0.5268288, 0.6635881, 0.7420592, 0.7799841, 0.7908091, 0.7824962, 
    0.7550047, 0.7052308, 0.6363831, 0.546421, 0.4342194, 0.3271011, 
    0.2539895, 0.1862741, 0.1015429, 0.00768932, -0.07776074, -0.1310218, 
    -0.1481579, -0.1403725, -0.135163, -0.1308205, -0.1172051, -0.07609003, 
    -0.06626932, -0.1100484, -0.1601827, -0.1389554, -0.02322895, 0.227192, 
    0.4801098, 0.6372901, 0.7581038, 0.8285891, 0.8605499, 0.8636217, 
    0.8369141,
  0.8859372, 0.8598702, 0.8193895, 0.7638259, 0.7110438, 0.6517936, 
    0.5864658, 0.5622275, 0.5233431, 0.443716, 0.3863952, 0.3838413, 
    0.355094, 0.2761848, 0.18879, 0.09128329, -0.006011514, -0.09894361, 
    -0.1857564, -0.2611129, -0.3257177, -0.3833014, -0.4299539, -0.4603045, 
    -0.4763111, -0.484588, -0.4753023, -0.4528309, -0.4520274, -0.4767042, 
    -0.507886, -0.5185698, -0.5071912, -0.4897636, -0.4852524, -0.4765307, 
    -0.4470255, -0.4081063, -0.3785705, -0.3565333, -0.314718, -0.2904844, 
    -0.2943395, -0.2967036, -0.2710263, -0.2334211, -0.2028158, -0.2034505, 
    -0.2077804, -0.1874037, -0.1647013, -0.1700907, -0.1683705, -0.1638901, 
    -0.1493387, -0.1373806, -0.1042906, -0.06687872, -0.07646462, 
    -0.04808664, 0.04398729, 0.1265506, 0.1731448, 0.196915, 0.2238875, 
    0.2238132, 0.2048375, 0.154614, 0.1422998, 0.1460969, 0.2259837, 
    0.5621531, 0.7457235, 0.566828, 0.2970131, 0.1176185, -0.05171249, 
    -0.2526022, -0.399526, -0.4817902, -0.5462568, -0.5820432, -0.5939511, 
    -0.5948819, -0.5818025, -0.5612624, -0.5089163, -0.4266579, -0.3419858, 
    -0.2530734, -0.1388571, -0.003007874, 0.1330794, 0.2467581, 0.3272787, 
    0.3700376, 0.380224, 0.3701857, 0.3494854, 0.3197452, 0.2879865, 0.26519, 
    0.2427396, 0.186243, 0.09705911, 0.006857473, -0.05754882, -0.09491368, 
    -0.1141239, -0.126341, -0.1137847, -0.0907529, -0.06162135, -0.04718181, 
    -0.02750587, -0.01393392, -0.02623171, -0.06036241, -0.06143966, 
    0.01237274, 0.2131834, 0.4967587, 0.6858118, 0.8062114, 0.8828628, 
    0.919575, 0.9271594, 0.9107071,
  0.9454147, 0.9213084, 0.8834018, 0.8528637, 0.8094079, 0.7440838, 
    0.6852142, 0.6483818, 0.6251124, 0.5583566, 0.4877257, 0.4635544, 
    0.4446543, 0.3591776, 0.2394885, 0.1286246, 0.02823565, -0.07312925, 
    -0.1692536, -0.2436849, -0.2986404, -0.3464828, -0.3858741, -0.4092337, 
    -0.4188884, -0.4225988, -0.4132648, -0.3904275, -0.3951674, -0.4225735, 
    -0.4428401, -0.4433102, -0.4210733, -0.3993831, -0.3904684, -0.3728276, 
    -0.3317571, -0.2861664, -0.2510922, -0.2283819, -0.207948, -0.2009647, 
    -0.1919414, -0.1861799, -0.1599505, -0.1310005, -0.1342174, -0.1546227, 
    -0.1409269, -0.1081417, -0.09717201, -0.1074612, -0.08671929, 
    -0.04579622, -0.01559539, -0.005096268, 0.008644849, 0.04499838, 
    0.05622076, 0.04587201, 0.09587841, 0.1473587, 0.1910617, 0.1847127, 
    0.1573675, 0.1744485, 0.1931938, 0.2297713, 0.2204039, 0.2649067, 
    0.2933299, 0.6074744, 0.8504531, 0.6312463, 0.3794816, 0.2045149, 
    0.01746844, -0.1829609, -0.3135282, -0.3857687, -0.4307219, -0.4744428, 
    -0.4965932, -0.5033203, -0.4972778, -0.4799752, -0.457371, -0.4219573, 
    -0.3671361, -0.2987758, -0.2219996, -0.1490273, -0.08221111, -0.01826327, 
    0.04405673, 0.09737217, 0.1437802, 0.1840302, 0.2201533, 0.2434041, 
    0.243683, 0.2122536, 0.1551445, 0.08236448, 0.008794941, -0.04818903, 
    -0.07167821, -0.08011152, -0.07678474, -0.06802458, -0.04821865, 
    -0.02666011, -0.0002614148, 0.02752388, 0.05044651, 0.05266391, 
    0.04507893, 0.03700383, 0.02551614, 0.05196273, 0.157194, 0.410125, 
    0.6658388, 0.8132405, 0.8976734, 0.9467587, 0.9644917, 0.9620201,
  0.9772737, 0.9566401, 0.9247933, 0.9075987, 0.8804334, 0.826207, 0.7753999, 
    0.7246782, 0.7067218, 0.6656398, 0.580489, 0.5365434, 0.5220467, 
    0.4484603, 0.3314729, 0.2174307, 0.1059972, -0.006142434, -0.1057167, 
    -0.1766627, -0.2393097, -0.2982589, -0.3406726, -0.3532037, -0.3525767, 
    -0.3538785, -0.3380473, -0.3198886, -0.3347349, -0.363464, -0.3759924, 
    -0.3567137, -0.3198698, -0.3075553, -0.3002437, -0.2737043, -0.222409, 
    -0.1700232, -0.1301539, -0.1187863, -0.1182966, -0.1143983, -0.1080685, 
    -0.1033113, -0.08030051, -0.07974754, -0.08549564, -0.07818492, 
    -0.05349284, -0.03147269, 0.004450634, 0.03479075, 0.06243467, 0.0749258, 
    0.07638162, 0.07018042, 0.09310218, 0.1147039, 0.1340477, 0.1379321, 
    0.1922701, 0.2466527, 0.3063443, 0.301234, 0.2708958, 0.3038482, 
    0.3158005, 0.3905766, 0.399062, 0.4286354, 0.4181938, 0.7619278, 
    0.9133552, 0.6275881, 0.4262026, 0.2459345, 0.04409733, -0.1290989, 
    -0.2334257, -0.301268, -0.338757, -0.3715261, -0.396793, -0.4183565, 
    -0.4144728, -0.4044176, -0.3953311, -0.3785452, -0.3331169, -0.2876661, 
    -0.2467521, -0.2008702, -0.1360266, -0.06895114, -0.0006201193, 
    0.05846468, 0.1076113, 0.1470777, 0.1772715, 0.1803321, 0.1561716, 
    0.1125999, 0.06543941, 0.01576526, -0.02164409, -0.04447103, -0.04569916, 
    -0.03448541, -0.01898267, -0.002167124, 0.02577042, 0.05432808, 
    0.07296909, 0.08379523, 0.1033915, 0.1178611, 0.117338, 0.1190635, 
    0.108526, 0.117714, 0.1476534, 0.2667966, 0.512947, 0.7433034, 0.8696645, 
    0.9321326, 0.9686136, 0.9834886,
  0.9595025, 0.9577621, 0.9486118, 0.9356105, 0.9151068, 0.8791253, 
    0.8494958, 0.816498, 0.7803952, 0.7388012, 0.6650003, 0.6201766, 
    0.5900108, 0.5221782, 0.4211028, 0.3125106, 0.1931579, 0.07177114, 
    -0.0230935, -0.1092792, -0.1954642, -0.257813, -0.2876162, -0.282703, 
    -0.2760513, -0.2854683, -0.2662621, -0.2439235, -0.2728835, -0.308619, 
    -0.3041157, -0.25949, -0.2270007, -0.2245562, -0.2154217, -0.1830211, 
    -0.129394, -0.07177661, -0.03490986, -0.0362592, -0.03237552, -0.0327674, 
    -0.03204063, -0.01303694, -0.0158428, -0.02224817, -0.002571853, 
    0.02585608, 0.07210365, 0.104625, 0.1127699, 0.09857586, 0.09237678, 
    0.0941612, 0.1048331, 0.1202983, 0.1610621, 0.181872, 0.184608, 0.180937, 
    0.2253921, 0.2675428, 0.3117242, 0.2989203, 0.3335262, 0.3842733, 
    0.5035111, 0.5777295, 0.5923231, 0.5596321, 0.6152174, 0.9687345, 
    0.863324, 0.5927921, 0.4355476, 0.2383568, 0.05549056, -0.07407245, 
    -0.1715511, -0.237896, -0.2660874, -0.2822674, -0.3064859, -0.3374319, 
    -0.3466527, -0.3370324, -0.3211805, -0.3231818, -0.306601, -0.2552422, 
    -0.1940362, -0.1557999, -0.1231452, -0.07708164, -0.02717588, 0.02093867, 
    0.06875543, 0.1056055, 0.1246433, 0.11808, 0.09218943, 0.05682864, 
    0.02513999, -0.001170669, -0.01672965, -0.01534576, 0.002834763, 
    0.02163392, 0.04215343, 0.06734558, 0.09669931, 0.1199407, 0.1379579, 
    0.1529239, 0.1704725, 0.1830662, 0.1886574, 0.1992009, 0.2018058, 
    0.1929251, 0.1948292, 0.2174607, 0.3142551, 0.5119116, 0.7208571, 
    0.8544446, 0.9208915, 0.9500834,
  0.8722702, 0.8972936, 0.9140912, 0.9124033, 0.8975389, 0.8800386, 
    0.8870637, 0.8918015, 0.8438974, 0.7945285, 0.7375374, 0.6930943, 
    0.6443321, 0.566146, 0.4811376, 0.3802303, 0.2517189, 0.134876, 
    0.0285572, -0.08794159, -0.1782696, -0.2276951, -0.2347875, -0.2189115, 
    -0.2093681, -0.2134862, -0.1947814, -0.1825933, -0.2213009, -0.2452795, 
    -0.2213976, -0.1734696, -0.1541487, -0.1539763, -0.1469867, -0.1110227, 
    -0.04466435, 0.02796928, 0.06481663, 0.05343271, 0.04298296, 0.03149639, 
    0.03227292, 0.04354292, 0.04495116, 0.06039811, 0.08091085, 0.1328488, 
    0.1764238, 0.1425128, 0.07100599, 0.05477678, 0.07841697, 0.1144594, 
    0.1360675, 0.1653652, 0.2022339, 0.2385873, 0.2457353, 0.2528611, 
    0.2799544, 0.3089546, 0.3223121, 0.3528194, 0.427735, 0.4949179, 
    0.6204765, 0.6883626, 0.7044721, 0.6352069, 0.9049617, 1.019819, 
    0.7327974, 0.5711884, 0.392072, 0.2028427, 0.05922282, -0.03186613, 
    -0.1142215, -0.1718559, -0.2042626, -0.2147308, -0.2340111, -0.2577458, 
    -0.2684897, -0.2728133, -0.2725464, -0.2598158, -0.2418511, -0.2157216, 
    -0.1792556, -0.1255588, -0.07906942, -0.03650555, 0.007575691, 
    0.04435487, 0.07220986, 0.0954372, 0.09842706, 0.07973987, 0.05315649, 
    0.03376984, 0.01854251, 0.007527575, 0.007314064, 0.0199092, 0.03976508, 
    0.06685114, 0.09998593, 0.1340529, 0.16536, 0.1894437, 0.2098143, 
    0.2240871, 0.2337458, 0.2404242, 0.2532351, 0.2715181, 0.2787892, 
    0.2710488, 0.2563173, 0.2589598, 0.2771302, 0.3218416, 0.443716, 
    0.6134558, 0.7523603, 0.8317923,
  0.6745245, 0.7395376, 0.7851769, 0.8134245, 0.8456185, 0.881918, 0.9199706, 
    0.9382977, 0.8765859, 0.8278576, 0.7959436, 0.7427123, 0.6746625, 
    0.5920192, 0.5156161, 0.4022272, 0.2735413, 0.1575638, 0.02431945, 
    -0.09277702, -0.1599804, -0.1830007, -0.1709549, -0.1606064, -0.1534536, 
    -0.1469585, -0.1316748, -0.1375154, -0.1716451, -0.1771102, -0.1451347, 
    -0.1048504, -0.09474218, -0.09343635, -0.08438183, -0.03714425, 
    0.05153013, 0.1326078, 0.1539929, 0.113203, 0.0971432, 0.1052286, 
    0.09835935, 0.09725072, 0.1116849, 0.1282037, 0.1879296, 0.2324722, 
    0.1643786, 0.05233708, 0.007222179, 0.05348228, 0.1259896, 0.1880509, 
    0.230527, 0.2780336, 0.3049935, 0.3146638, 0.3144892, 0.3344889, 
    0.3457999, 0.3494331, 0.3651592, 0.4400546, 0.5095283, 0.5811821, 
    0.7113853, 0.7520288, 0.7047198, 0.9141421, 1.091907, 0.8427062, 
    0.6497748, 0.502702, 0.3088472, 0.1659602, 0.0750203, 0.0005358756, 
    -0.07139535, -0.1164086, -0.1415314, -0.1605052, -0.1743004, -0.193401, 
    -0.204781, -0.2063854, -0.2070681, -0.2046303, -0.1977807, -0.1683806, 
    -0.128382, -0.07811417, -0.02756429, 0.004993991, 0.03077926, 0.06084001, 
    0.08125436, 0.08865444, 0.0821566, 0.065937, 0.04863701, 0.03166416, 
    0.01702942, 0.0118164, 0.01765118, 0.03590246, 0.0641514, 0.09859731, 
    0.1393117, 0.1798384, 0.2120038, 0.23706, 0.2634262, 0.2893541, 
    0.3056259, 0.3134919, 0.326018, 0.3430066, 0.346673, 0.3428315, 
    0.3361844, 0.3297176, 0.3322395, 0.3390175, 0.3490956, 0.3997402, 
    0.4954144, 0.5936579,
  0.5117896, 0.5554398, 0.604651, 0.6845981, 0.7944321, 0.8863958, 0.9336934, 
    0.9410363, 0.8821142, 0.8676155, 0.8371212, 0.7609205, 0.6867089, 
    0.6083208, 0.5155573, 0.3828791, 0.2591258, 0.1195124, -0.02363588, 
    -0.101973, -0.1283994, -0.130555, -0.1162908, -0.1114123, -0.1003641, 
    -0.08669703, -0.08028378, -0.09879583, -0.1218297, -0.1207688, 
    -0.08894552, -0.0556676, -0.04626697, -0.0439418, -0.03476634, 
    0.03068966, 0.1439794, 0.2229322, 0.230795, 0.1788466, 0.1466901, 
    0.139373, 0.132679, 0.1535072, 0.1709904, 0.2118538, 0.2607127, 
    0.1964109, 0.07705633, 0.01455135, 0.02870964, 0.1268815, 0.2338958, 
    0.2985257, 0.3621872, 0.4250869, 0.4601601, 0.4652165, 0.4700077, 
    0.4681197, 0.4489069, 0.4341249, 0.4702433, 0.5372941, 0.6204043, 
    0.7211749, 0.7879195, 0.7970441, 0.9807855, 1.121874, 0.8946114, 
    0.6958776, 0.567295, 0.3791308, 0.2394239, 0.1549473, 0.08295497, 
    0.01377115, -0.0297243, -0.06285752, -0.1022371, -0.1241062, -0.1233782, 
    -0.1302355, -0.147495, -0.1584584, -0.1556828, -0.1420472, -0.1373372, 
    -0.1270741, -0.1008009, -0.05364246, 0.003091201, 0.0472042, 0.07475062, 
    0.08835123, 0.09514264, 0.09091433, 0.07302789, 0.05433454, 0.04039396, 
    0.02143451, 0.003861763, -0.005321324, -5.77122e-05, 0.01773664, 
    0.05093834, 0.09944326, 0.1522798, 0.1992514, 0.2418149, 0.2803786, 
    0.3124988, 0.3373179, 0.3616791, 0.3856404, 0.401159, 0.4066492, 
    0.409978, 0.4186677, 0.4222975, 0.4149517, 0.3966019, 0.397827, 
    0.4116875, 0.4014878, 0.4058529, 0.453173,
  0.5345438, 0.546647, 0.5965824, 0.7157282, 0.8379246, 0.8949775, 0.9246593, 
    0.9230452, 0.8912082, 0.8982739, 0.8307763, 0.7477138, 0.6861104, 
    0.5966803, 0.4691634, 0.338041, 0.1929487, 0.02713549, -0.07157636, 
    -0.09195191, -0.0947455, -0.09180969, -0.0721501, -0.0609105, 
    -0.05011996, -0.04747333, -0.04534869, -0.05926736, -0.08008536, 
    -0.08259046, -0.04910511, -0.01657243, -0.007959548, -0.008359835, 
    0.009891342, 0.09866501, 0.2235065, 0.2860937, 0.2686674, 0.2166914, 
    0.2013242, 0.1822991, 0.1786749, 0.2008154, 0.21414, 0.2588124, 
    0.2431532, 0.1531775, 0.09786518, 0.06012891, 0.09871693, 0.2376159, 
    0.3344234, 0.4163945, 0.522254, 0.6123965, 0.6572626, 0.6555169, 
    0.6259854, 0.5861619, 0.5569346, 0.5588618, 0.5983209, 0.66833, 
    0.7533227, 0.8459529, 0.94103, 1.088447, 1.118575, 0.8896293, 0.7128696, 
    0.5885409, 0.4091465, 0.2799747, 0.2075501, 0.1409993, 0.07651186, 
    0.03989349, 0.01021662, -0.02776146, -0.06550409, -0.09029627, 
    -0.09614578, -0.09913732, -0.1090509, -0.1096163, -0.106712, -0.1056163, 
    -0.1090264, -0.09076305, -0.06052705, -0.02684303, 0.01765203, 
    0.05675599, 0.07984921, 0.08685534, 0.08570872, 0.07755055, 0.06339912, 
    0.05106021, 0.02628472, -0.003455848, -0.01736329, -0.02347651, 
    -0.02425313, -0.01259241, 0.01726875, 0.06261061, 0.1200664, 0.181247, 
    0.2377291, 0.2849697, 0.3260704, 0.3652496, 0.4016034, 0.4319659, 
    0.4530922, 0.4660717, 0.4750737, 0.4858965, 0.4953847, 0.4976999, 
    0.492408, 0.481077, 0.4672275, 0.453089, 0.4645878, 0.5007473,
  0.5892334, 0.6341575, 0.7077293, 0.7924875, 0.8531984, 0.8866831, 
    0.9108621, 0.9048684, 0.9142003, 0.8765346, 0.7821749, 0.7322083, 
    0.6538562, 0.5295452, 0.3979534, 0.2461841, 0.06486166, -0.04705888, 
    -0.07078269, -0.06653143, -0.0666995, -0.05146465, -0.03476476, 
    -0.02929453, -0.01991108, -0.01320451, -0.0110769, -0.02417307, 
    -0.04136402, -0.04294289, -0.01704392, 0.008473936, 0.01507615, 
    0.02142272, 0.04711725, 0.1453075, 0.2726346, 0.3197728, 0.3014865, 
    0.2514639, 0.2223764, 0.195892, 0.2004012, 0.2354399, 0.2418983, 
    0.2568303, 0.2180879, 0.170579, 0.1483133, 0.09238485, 0.1860555, 
    0.3292327, 0.416356, 0.5352305, 0.6699777, 0.788623, 0.8453826, 
    0.8287681, 0.7714905, 0.7212055, 0.6934003, 0.7046283, 0.774443, 
    0.873603, 0.9815297, 1.083114, 1.141208, 1.044442, 0.8288522, 0.6932843, 
    0.5693922, 0.406875, 0.298235, 0.2307874, 0.1732766, 0.1252132, 
    0.09259111, 0.06633382, 0.0345623, 0.007673547, -0.0212985, -0.05360657, 
    -0.07143795, -0.0742593, -0.08430766, -0.0935066, -0.0886516, 
    -0.06925328, -0.06580305, -0.06664164, -0.0519458, -0.02529509, 
    0.01491695, 0.0548073, 0.07788892, 0.08530162, 0.08429261, 0.07297193, 
    0.05562675, 0.03353233, 0.005958695, -0.006850272, -0.02023964, 
    -0.04321345, -0.05632087, -0.0570247, -0.0422687, -0.007404864, 
    0.04765519, 0.1161664, 0.1906355, 0.2584555, 0.3125052, 0.3565778, 
    0.3982317, 0.4382487, 0.4733046, 0.5013771, 0.5217251, 0.5359865, 
    0.5479439, 0.562322, 0.5681511, 0.5644972, 0.5524194, 0.5470741, 
    0.5557159, 0.5664266,
  0.6904751, 0.7311405, 0.7688367, 0.8057613, 0.8469248, 0.8844684, 
    0.9010957, 0.9126834, 0.8896627, 0.8054088, 0.751375, 0.6820467, 
    0.5617369, 0.4349655, 0.2739812, 0.08826024, -0.03077155, -0.05835252, 
    -0.0543561, -0.0465628, -0.0355123, -0.01538116, -0.007306203, 
    0.0003665164, 0.00932027, 0.01474921, 0.01491714, 0.003922142, 
    -0.01120372, -0.02254506, -0.00863472, 0.01844202, 0.02824868, 
    0.03821624, 0.06688491, 0.1635116, 0.2970491, 0.3340049, 0.3046131, 
    0.2776152, 0.2577987, 0.2289055, 0.2120938, 0.245873, 0.2575549, 
    0.2605504, 0.246831, 0.2331021, 0.1657474, 0.1308808, 0.2749534, 
    0.3806015, 0.4671441, 0.5953864, 0.7506055, 0.9026951, 0.9704744, 
    0.9392555, 0.8661101, 0.8233825, 0.8554051, 0.9573171, 1.062434, 
    1.126905, 1.140129, 1.062818, 0.8984841, 0.7391573, 0.6417909, 0.5196433, 
    0.3858405, 0.2970126, 0.2276632, 0.1738842, 0.148801, 0.1350013, 
    0.1052075, 0.07331689, 0.05092829, 0.03222024, -0.0004102215, -0.0357751, 
    -0.05511319, -0.05866863, -0.06456083, -0.07187399, -0.07563708, 
    -0.06731705, -0.06019092, -0.05366635, -0.03234614, -0.009608559, 
    0.01213964, 0.03358943, 0.05161938, 0.06148333, 0.05993218, 0.05460627, 
    0.04611118, 0.02798565, 0.008918323, -0.00739079, -0.03546555, 
    -0.05589005, -0.06908407, -0.07900704, -0.07973943, -0.07315688, 
    -0.04806742, 0.0002907068, 0.07005264, 0.1547625, 0.2389416, 0.3112121, 
    0.3669287, 0.4124609, 0.4534841, 0.4906613, 0.5242556, 0.5539108, 
    0.5746651, 0.5886762, 0.6049556, 0.6245949, 0.6416203, 0.6584726, 
    0.6632944, 0.6686546,
  0.7553786, 0.7837706, 0.8053432, 0.8315997, 0.8634392, 0.8858525, 
    0.8903451, 0.861801, 0.8008033, 0.7515823, 0.6791343, 0.5647189, 
    0.4390514, 0.2720741, 0.0881629, -0.02253104, -0.05868043, -0.05698209, 
    -0.04012401, -0.0281113, -0.01140965, 0.00366177, 0.009126469, 
    0.02352751, 0.03259424, 0.03269065, 0.03341348, 0.02690767, 0.01353925, 
    -0.00749357, -0.01190221, 0.01078403, 0.02439589, 0.0395206, 0.07176252, 
    0.149741, 0.2870522, 0.3432824, 0.3179178, 0.3022012, 0.2792968, 
    0.2509258, 0.2288887, 0.2532833, 0.2712003, 0.2600004, 0.2413515, 
    0.2362749, 0.1643459, 0.1828406, 0.3275592, 0.4106047, 0.4863071, 
    0.5934854, 0.736267, 0.8977662, 1.031688, 1.070876, 1.0608, 1.070018, 
    1.105868, 1.119901, 1.08506, 0.9942307, 0.8631682, 0.7314732, 0.6400886, 
    0.5590287, 0.4480853, 0.3499028, 0.2777119, 0.209542, 0.1719934, 
    0.1557679, 0.1452106, 0.1296806, 0.1119165, 0.09369101, 0.07416859, 
    0.0508531, 0.02489982, 0.001860887, -0.02746233, -0.05081586, 
    -0.06014601, -0.06617989, -0.07044234, -0.0621401, -0.04655244, 
    -0.04812774, -0.04455116, -0.02333297, 0.003193706, 0.02759006, 
    0.04369096, 0.05156371, 0.05538586, 0.05515574, 0.04405314, 0.02145933, 
    0.008077756, -0.0009093285, -0.02026339, -0.03469407, -0.04670119, 
    -0.06375808, -0.07875563, -0.0892925, -0.09281264, -0.0816834, 
    -0.05078771, 0.005370259, 0.0836157, 0.1734999, 0.2626442, 0.3374969, 
    0.3949378, 0.4403291, 0.4797613, 0.5178019, 0.5549676, 0.5867871, 
    0.6134381, 0.6386418, 0.6623504, 0.6859189, 0.7104917, 0.7320684,
  0.7616335, 0.785585, 0.8097879, 0.8309544, 0.8424213, 0.8382525, 0.8099422, 
    0.7644342, 0.7190862, 0.6461939, 0.5397426, 0.408375, 0.2345571, 
    0.0646846, -0.02865284, -0.05542732, -0.06011453, -0.04485049, 
    -0.02729419, -0.01536707, 0.004250683, 0.01819686, 0.02329472, 
    0.03576195, 0.04188653, 0.04271067, 0.05213493, 0.0492796, 0.03920711, 
    0.02178524, 0.001669563, 0.0134936, 0.02463962, 0.03986577, 0.07516935, 
    0.1262896, 0.2445912, 0.3467037, 0.3363465, 0.3087305, 0.3011224, 
    0.2892549, 0.2615118, 0.2501562, 0.2716464, 0.2768207, 0.2507766, 
    0.2443509, 0.1857669, 0.2310558, 0.3464258, 0.4164774, 0.4798858, 
    0.5413659, 0.6438448, 0.7606068, 0.8794966, 0.9652336, 1.006413, 
    0.9988004, 0.9489571, 0.8674656, 0.7714269, 0.6771753, 0.6031008, 
    0.5380415, 0.459031, 0.3742067, 0.3099785, 0.2476604, 0.1947408, 
    0.1687601, 0.1591395, 0.1387327, 0.1290025, 0.1316193, 0.1288147, 
    0.1037985, 0.0774412, 0.05990427, 0.03923049, 0.01506006, -0.008792505, 
    -0.02920508, -0.04089055, -0.04753542, -0.06029595, -0.07524899, 
    -0.06449167, -0.04441609, -0.03596434, -0.0248204, -0.008378215, 
    0.004068203, 0.01817807, 0.02937578, 0.0356238, 0.03826213, 0.03678191, 
    0.03074077, 0.0253884, 0.01133475, -0.006703034, -0.01450044, 
    -0.02746238, -0.05101359, -0.07329249, -0.09121349, -0.104631, 
    -0.1134999, -0.1162288, -0.1043069, -0.07017733, -0.0124343, 0.0662488, 
    0.1595419, 0.2525486, 0.3324061, 0.3956112, 0.445023, 0.4882488, 
    0.5295402, 0.569585, 0.6074066, 0.6448275, 0.6796567, 0.7101746, 0.7366015,
  0.7113176, 0.7347251, 0.749332, 0.7525475, 0.7429242, 0.7221985, 0.6944383, 
    0.6541378, 0.5825696, 0.4761208, 0.3333216, 0.1601008, 0.02221939, 
    -0.04657042, -0.06753593, -0.06320113, -0.04952165, -0.03030927, 
    -0.01296435, 0.0009419583, 0.0191118, 0.03013719, 0.03454903, 0.04614776, 
    0.05397274, 0.06099289, 0.07544689, 0.06662971, 0.05881588, 0.05155399, 
    0.02356484, 0.020804, 0.0262717, 0.03707934, 0.07044926, 0.1087199, 
    0.1800423, 0.308093, 0.3703675, 0.3340411, 0.2998547, 0.3011723, 
    0.2864227, 0.2488067, 0.2427177, 0.2635155, 0.252318, 0.2329102, 
    0.2016894, 0.2679085, 0.3578556, 0.411397, 0.4755165, 0.5050151, 
    0.5453393, 0.5984709, 0.6517545, 0.6859064, 0.6940115, 0.6759503, 
    0.6409323, 0.5933535, 0.5427334, 0.4891637, 0.4280695, 0.3633145, 
    0.3115071, 0.2639461, 0.2109799, 0.18135, 0.1694343, 0.1555117, 
    0.1503333, 0.1430248, 0.1380048, 0.1287615, 0.1254425, 0.1161068, 
    0.09812441, 0.0733208, 0.04645606, 0.02926444, 0.01283441, -0.01495253, 
    -0.03843599, -0.04477763, -0.04400219, -0.04959271, -0.05691727, 
    -0.05494709, -0.04692456, -0.03717281, -0.0177787, 0.001008891, 
    0.01240937, 0.02311915, 0.03376868, 0.03728703, 0.03574049, 0.03243417, 
    0.03053653, 0.02601618, 0.01828206, 0.008900613, -0.003948361, 
    -0.01987252, -0.03914836, -0.0584996, -0.07565024, -0.09192096, 
    -0.107003, -0.1206635, -0.1297293, -0.1256877, -0.102145, -0.05469866, 
    0.01692607, 0.1053344, 0.1994936, 0.2888079, 0.3648621, 0.4269405, 
    0.4781891, 0.5223788, 0.5636977, 0.6054202, 0.6459364, 0.6812606,
  0.5927449, 0.612492, 0.6246278, 0.6275246, 0.6200628, 0.5986617, 0.5521847, 
    0.4701777, 0.3525402, 0.2062649, 0.0619825, -0.03008742, -0.06586807, 
    -0.07630537, -0.07429435, -0.0620396, -0.0419062, -0.01365279, 
    0.002288871, 0.01319527, 0.03180555, 0.04362805, 0.04982537, 0.05804702, 
    0.06342014, 0.07733876, 0.09232792, 0.07678554, 0.07467345, 0.07692501, 
    0.05135322, 0.03021102, 0.01675091, 0.01877712, 0.04718123, 0.09487684, 
    0.1399368, 0.2261225, 0.3353217, 0.3739821, 0.3317431, 0.3106248, 
    0.3041574, 0.2908527, 0.2535622, 0.2456457, 0.2315423, 0.2231785, 
    0.2264682, 0.2748635, 0.3625886, 0.3946857, 0.443555, 0.4702063, 
    0.4891825, 0.5063879, 0.5215154, 0.5301108, 0.5289949, 0.5116755, 
    0.4812713, 0.4391243, 0.3904098, 0.3405671, 0.3009264, 0.2620575, 
    0.2167166, 0.1764556, 0.1633537, 0.1545148, 0.1418208, 0.1412392, 
    0.1548809, 0.1524922, 0.1388368, 0.1338852, 0.1378427, 0.1294847, 
    0.108281, 0.09042927, 0.06761818, 0.04422011, 0.02920887, 0.01251047, 
    -0.009631231, -0.02817179, -0.04185657, -0.04702327, -0.04988968, 
    -0.04822986, -0.03665568, -0.02366706, -0.0179824, -0.007831126, 
    0.004695617, 0.01241933, 0.02114056, 0.03265063, 0.03780843, 0.03863803, 
    0.04012886, 0.04141769, 0.03615659, 0.02610585, 0.01393691, 0.001004636, 
    -0.01667562, -0.03704095, -0.05429678, -0.07308008, -0.09107979, 
    -0.1066078, -0.1213739, -0.1338885, -0.1426512, -0.1436012, -0.1326761, 
    -0.1034526, -0.05290743, 0.01946223, 0.1087565, 0.2044467, 0.2957356, 
    0.3749488, 0.4387466, 0.4897446, 0.5316116, 0.5660959,
  0.3998064, 0.4256418, 0.4349729, 0.4261314, 0.3940042, 0.3340604, 
    0.2477157, 0.1439728, 0.03950448, -0.03949978, -0.07996023, -0.0959972, 
    -0.1002058, -0.08612062, -0.07034737, -0.05243085, -0.02693508, 
    -0.006689455, 0.008147553, 0.0288862, 0.04277623, 0.04654838, 0.05784269, 
    0.07063821, 0.06977683, 0.07320372, 0.08444051, 0.08861375, 0.09585079, 
    0.08248179, 0.06882872, 0.05627878, 0.03009325, 0.01242276, 0.01078925, 
    0.04944907, 0.09752208, 0.1548798, 0.2372686, 0.3299268, 0.3718323, 
    0.3560957, 0.3049338, 0.2944327, 0.2658726, 0.2573111, 0.2413073, 
    0.2604865, 0.252088, 0.2619413, 0.3514048, 0.3751871, 0.4123899, 
    0.4265493, 0.4313502, 0.4316183, 0.4292824, 0.417333, 0.3999344, 
    0.3712369, 0.3423456, 0.3084306, 0.2795224, 0.2472331, 0.2088671, 
    0.1644417, 0.1512647, 0.1437773, 0.1297195, 0.1126311, 0.1199987, 
    0.1250984, 0.1305646, 0.1416916, 0.1500586, 0.1461276, 0.1327498, 
    0.1210003, 0.1075068, 0.09472032, 0.07089297, 0.04173052, 0.02068114, 
    0.0081334, -0.005211558, -0.01875286, -0.02854356, -0.02928571, 
    -0.0347463, -0.04388926, -0.04495154, -0.02892775, -0.01086853, 
    0.0007138848, 0.01233773, 0.02584717, 0.03164691, 0.03731374, 0.04375491, 
    0.04604618, 0.04207288, 0.04421452, 0.04742444, 0.03891051, 0.02689418, 
    0.01842728, 0.002183646, -0.01823783, -0.0362533, -0.05835953, 
    -0.08073035, -0.09735488, -0.1137165, -0.1311306, -0.1442802, -0.1526206, 
    -0.1618384, -0.1690837, -0.1706268, -0.1600409, -0.1324842, -0.08330014, 
    -0.01479764, 0.06747231, 0.1535843, 0.2340602, 0.3028711, 0.3585523,
  0.03348726, 0.05674309, 0.06343292, 0.05151203, 0.02330545, -0.01509604, 
    -0.05746867, -0.09328566, -0.1104392, -0.1168297, -0.1226785, -0.1168249, 
    -0.1039909, -0.08881161, -0.06906813, -0.04188632, -0.01985614, 
    -0.005996108, 0.01309283, 0.03188176, 0.04086523, 0.04840517, 0.06043045, 
    0.06798527, 0.0705616, 0.07500352, 0.08146372, 0.09412111, 0.1008601, 
    0.07776747, 0.07164377, 0.06368992, 0.04269036, 0.02413584, 0.006322697, 
    0.02004243, 0.05352626, 0.09776423, 0.1452473, 0.2148306, 0.3001141, 
    0.3603278, 0.3662043, 0.3451608, 0.2975174, 0.28177, 0.2685898, 
    0.2944875, 0.2535115, 0.2657742, 0.3363225, 0.3426003, 0.3637057, 
    0.3680843, 0.3633128, 0.3503976, 0.3357036, 0.3157458, 0.3042628, 
    0.2845513, 0.2656838, 0.2400214, 0.2054465, 0.1631635, 0.1366354, 
    0.118867, 0.1215911, 0.1076262, 0.116772, 0.1115981, 0.1126377, 
    0.1190075, 0.1288185, 0.1410578, 0.1412, 0.1378639, 0.1392028, 0.1300182, 
    0.1063558, 0.09618752, 0.08304034, 0.0575882, 0.03496323, 0.01558832, 
    -0.002849232, -0.01798739, -0.03237217, -0.04454347, -0.04861445, 
    -0.03888851, -0.03017347, -0.02536368, -0.0165507, -0.003494203, 
    0.004257798, 0.01239267, 0.02295651, 0.03358132, 0.04225177, 0.05303966, 
    0.05777985, 0.05539522, 0.0513787, 0.04663917, 0.03655332, 0.02433336, 
    0.008679986, -0.01337516, -0.03155559, -0.04585615, -0.06772676, 
    -0.09082872, -0.1077937, -0.1236132, -0.1418909, -0.1555127, -0.1678797, 
    -0.1786745, -0.1877562, -0.1950374, -0.1996901, -0.1988656, -0.1898124, 
    -0.169199, -0.1359677, -0.09200779, -0.04513437, -0.001662739,
  -0.1652932, -0.1556365, -0.1498077, -0.1463602, -0.1456312, -0.1459963, 
    -0.14474, -0.143241, -0.1429047, -0.1363269, -0.1238409, -0.1085085, 
    -0.0953742, -0.08080614, -0.05892758, -0.03632834, -0.0175302, 
    0.001264572, 0.02136054, 0.03330184, 0.04277547, 0.05642256, 0.0641461, 
    0.06356999, 0.07366849, 0.09269334, 0.1057923, 0.1106278, 0.104798, 
    0.08872505, 0.08586831, 0.07288235, 0.05298445, 0.03008358, 0.005363189, 
    -0.005368911, 0.008845985, 0.05176818, 0.09598236, 0.1368992, 0.1860148, 
    0.2540066, 0.3241547, 0.3627958, 0.3611301, 0.3378666, 0.3012452, 
    0.2833824, 0.2624357, 0.3015417, 0.32356, 0.3235629, 0.3259008, 0.319751, 
    0.3069575, 0.2905054, 0.2810302, 0.2639225, 0.2516227, 0.2322013, 
    0.2089029, 0.1778758, 0.1412196, 0.112502, 0.09921139, 0.07923119, 
    0.09260171, 0.09133302, 0.09117063, 0.09423314, 0.1055586, 0.12127, 
    0.1268135, 0.1276399, 0.1291037, 0.1287739, 0.1287204, 0.1196269, 
    0.1030262, 0.08952831, 0.06890235, 0.04847832, 0.03025853, 0.01139584, 
    -0.004764222, -0.01400754, -0.01792933, -0.02474708, -0.03597726, 
    -0.04328369, -0.04000641, -0.0258695, -0.00910835, 0.006411493, 
    0.01810289, 0.02452944, 0.03193526, 0.04447295, 0.05507097, 0.06113559, 
    0.0629219, 0.06348352, 0.06408963, 0.06042975, 0.04824248, 0.0345158, 
    0.02416897, 0.008472621, -0.01555553, -0.03546387, -0.05400488, 
    -0.07936171, -0.09924902, -0.1140762, -0.1349788, -0.1500997, -0.1625283, 
    -0.1804928, -0.1953499, -0.2030371, -0.2111521, -0.2175652, -0.2186033, 
    -0.2156924, -0.2123864, -0.2063348, -0.1945666, -0.1790613,
  -0.2056967, -0.1975701, -0.1922488, -0.1872132, -0.1814079, -0.1760887, 
    -0.1712081, -0.1618006, -0.1471261, -0.130141, -0.1169847, -0.1064287, 
    -0.09273528, -0.07352965, -0.05073572, -0.03071553, -0.0123608, 
    0.006265166, 0.02199838, 0.033699, 0.04562094, 0.05697709, 0.06362139, 
    0.06736649, 0.07536495, 0.08497889, 0.09388103, 0.09704864, 0.09357073, 
    0.09668711, 0.09856264, 0.07997282, 0.06183531, 0.04568437, 0.02361172, 
    -0.004896864, -0.02179871, -0.01025458, 0.02246344, 0.06986041, 
    0.1187114, 0.1650915, 0.2144423, 0.2707296, 0.3221903, 0.3524369, 
    0.3587559, 0.3498418, 0.3378852, 0.317081, 0.2857389, 0.285338, 
    0.2835844, 0.2766508, 0.2622213, 0.2408116, 0.2309589, 0.2186783, 
    0.2077779, 0.18745, 0.1562025, 0.136236, 0.1086118, 0.07905282, 
    0.07263473, 0.06371087, 0.06479158, 0.06989588, 0.07995054, 0.08983624, 
    0.0989359, 0.1111633, 0.1211855, 0.1382659, 0.1538064, 0.1534878, 
    0.1455899, 0.1314079, 0.1167592, 0.1023275, 0.07799757, 0.05377296, 
    0.03424044, 0.01523247, -0.002113424, -0.01621034, -0.02924559, 
    -0.03784739, -0.03741335, -0.03297034, -0.02929891, -0.02156547, 
    -0.01020035, -0.0002095103, 0.009855494, 0.02117601, 0.03390044, 
    0.04716951, 0.05750273, 0.06502101, 0.06918199, 0.06908534, 0.06755157, 
    0.0663709, 0.05739294, 0.04314493, 0.03323251, 0.01804914, -0.005654573, 
    -0.02350825, -0.03898069, -0.06416619, -0.08537909, -0.1018345, -0.12386, 
    -0.140312, -0.1547282, -0.1742409, -0.1918926, -0.2046513, -0.2169302, 
    -0.2275063, -0.2318236, -0.2313639, -0.2307069, -0.2295118, -0.2250798, 
    -0.216008,
  -0.2197051, -0.2124156, -0.2047819, -0.1985478, -0.1920827, -0.1839945, 
    -0.1734388, -0.1582893, -0.1417452, -0.1261344, -0.1114423, -0.09852637, 
    -0.08333161, -0.06383547, -0.04424105, -0.02534641, -0.005324662, 
    0.01193335, 0.02556076, 0.0388403, 0.05067959, 0.05790358, 0.06362364, 
    0.07267346, 0.08256699, 0.08582284, 0.08390914, 0.08329105, 0.08807545, 
    0.09895234, 0.09391615, 0.0765709, 0.0674184, 0.05583008, 0.03814377, 
    0.01430666, -0.005334724, -0.01361404, -0.01396276, 0.00242186, 
    0.03533128, 0.08125597, 0.1318281, 0.1785432, 0.2226142, 0.2645833, 
    0.2947337, 0.3073213, 0.2995641, 0.2810512, 0.265811, 0.2581226, 
    0.2507933, 0.238626, 0.2267126, 0.2057324, 0.1955627, 0.1811267, 
    0.1622746, 0.1515194, 0.1231993, 0.09820122, 0.07942513, 0.05913228, 
    0.05055395, 0.04783089, 0.05536346, 0.07711971, 0.09369689, 0.09807914, 
    0.09910762, 0.112332, 0.1339513, 0.1490871, 0.1491836, 0.139978, 
    0.1284346, 0.1156652, 0.1061441, 0.09090494, 0.07121885, 0.05287283, 
    0.0311436, 0.01274461, 0.0006480068, -0.009013712, -0.01622717, 
    -0.02249916, -0.03250808, -0.0407113, -0.0371299, -0.02258885, 
    -0.004637174, 0.01144223, 0.02528758, 0.03646317, 0.04692841, 0.05754094, 
    0.06426337, 0.06704824, 0.07078205, 0.07590252, 0.07808955, 0.07422934, 
    0.06496222, 0.05277394, 0.04029278, 0.02686712, 0.007984653, -0.01303545, 
    -0.03354862, -0.05691725, -0.07784796, -0.09820241, -0.1174958, 
    -0.1328472, -0.1494728, -0.1672219, -0.1836265, -0.1997176, -0.2141912, 
    -0.2234738, -0.2293584, -0.2333585, -0.2346215, -0.232746, -0.2290603, 
    -0.2249422,
  -0.2198998, -0.2131844, -0.2054735, -0.1983021, -0.1905136, -0.1809393, 
    -0.1698541, -0.1548703, -0.1355365, -0.1191423, -0.1072984, -0.09383316, 
    -0.07620323, -0.05766249, -0.03927086, -0.02035162, -0.001930386, 
    0.01411802, 0.02725269, 0.03948158, 0.05154318, 0.06007759, 0.06525912, 
    0.0723124, 0.08329448, 0.0936407, 0.1013741, 0.1080958, 0.1117034, 
    0.1081716, 0.09290384, 0.08289504, 0.07698594, 0.06066206, 0.03788972, 
    0.0113398, -0.004952619, -0.0134987, -0.02090866, -0.02003236, 
    -0.01153024, 0.00666118, 0.03991903, 0.08645637, 0.1353153, 0.1795339, 
    0.2130473, 0.2314083, 0.2352056, 0.2307732, 0.2241782, 0.219613, 
    0.2103427, 0.1953577, 0.1860726, 0.1665249, 0.1534467, 0.1471766, 
    0.1262897, 0.1120825, 0.09689799, 0.07637495, 0.06070057, 0.04628193, 
    0.03539418, 0.03917451, 0.0563955, 0.07973796, 0.09876925, 0.09923619, 
    0.09725881, 0.1146919, 0.1334407, 0.1321026, 0.1240814, 0.1279221, 
    0.1295114, 0.121119, 0.1083163, 0.09063528, 0.07073408, 0.04923286, 
    0.03059188, 0.01371052, -0.003592089, -0.01745158, -0.0271254, 
    -0.0330666, -0.03300864, -0.02903915, -0.02501194, -0.01827636, 
    -0.008010427, 0.00323011, 0.01598397, 0.02876642, 0.0402948, 0.0505549, 
    0.0595675, 0.06825389, 0.07730918, 0.0823582, 0.07897627, 0.07302253, 
    0.06791263, 0.0590353, 0.04616564, 0.03032196, 0.01076451, -0.008098438, 
    -0.02588555, -0.04634607, -0.06750256, -0.08845696, -0.1076041, 
    -0.1252976, -0.1429886, -0.1608381, -0.1793406, -0.1964594, -0.2106763, 
    -0.2223418, -0.2300155, -0.234084, -0.2356048, -0.2343438, -0.2308113, 
    -0.2256882,
  -0.2205098, -0.2135686, -0.2044377, -0.1958684, -0.1873182, -0.1761101, 
    -0.1622237, -0.1460298, -0.1300331, -0.1156838, -0.100147, -0.08478012, 
    -0.0693405, -0.05237366, -0.03405073, -0.01509199, 0.002810359, 
    0.01761546, 0.03141008, 0.0442898, 0.05449257, 0.06191048, 0.06838964, 
    0.07573584, 0.08374207, 0.09036399, 0.09964164, 0.1134081, 0.119021, 
    0.1060723, 0.08995076, 0.08551005, 0.07801849, 0.06594948, 0.05159314, 
    0.03016154, 0.01308864, 0.000332579, -0.01220734, -0.027855, -0.03771008, 
    -0.0354623, -0.02588601, -0.003585063, 0.03123551, 0.07356019, 0.11565, 
    0.1503533, 0.1702218, 0.1747437, 0.1759906, 0.1754822, 0.1647666, 
    0.1518381, 0.1454619, 0.1329861, 0.1158284, 0.1067666, 0.09544592, 
    0.07860942, 0.06426595, 0.04747942, 0.02824041, 0.01785417, 0.02116191, 
    0.03730905, 0.06380877, 0.08747777, 0.09147054, 0.08770084, 0.09582329, 
    0.1143858, 0.1270137, 0.1340852, 0.148549, 0.1572897, 0.1471356, 
    0.1347187, 0.1213036, 0.09827828, 0.07544956, 0.05801256, 0.03892169, 
    0.01853953, 0.00346075, -0.007075384, -0.01552321, -0.02325502, 
    -0.03263577, -0.03932697, -0.0348055, -0.0193318, -0.0007781908, 
    0.01509938, 0.02870489, 0.03980493, 0.04992375, 0.05947133, 0.06759317, 
    0.07408944, 0.07941751, 0.08375391, 0.08363362, 0.07846436, 0.07330053, 
    0.06504115, 0.05029592, 0.03411264, 0.01675733, -0.002033643, 
    -0.02242827, -0.04417109, -0.06615925, -0.08711848, -0.1053787, 
    -0.1225087, -0.139149, -0.1567359, -0.1747457, -0.1916934, -0.2070863, 
    -0.2187544, -0.2266113, -0.2313384, -0.2331326, -0.2319624, -0.2287841, 
    -0.2250341,
  -0.2173688, -0.210402, -0.2015792, -0.1926786, -0.1834732, -0.1712267, 
    -0.1575547, -0.1426034, -0.125285, -0.1093266, -0.09535614, -0.08111487, 
    -0.06485773, -0.04777362, -0.02977573, -0.01144385, 0.005107276, 
    0.01977823, 0.03374808, 0.04593181, 0.05536917, 0.06223353, 0.06904821, 
    0.07881624, 0.09041843, 0.09750941, 0.09783655, 0.09559156, 0.09582132, 
    0.09551723, 0.09516221, 0.09321888, 0.08426426, 0.07381292, 0.05659585, 
    0.03028052, 0.008072048, -0.003632382, -0.006101616, -0.008315712, 
    -0.01697911, -0.03466493, -0.04957397, -0.04903005, -0.03760983, 
    -0.0173907, 0.01043066, 0.04128419, 0.06956501, 0.08870061, 0.09812418, 
    0.1009916, 0.09765051, 0.09070174, 0.08623489, 0.08223586, 0.07226797, 
    0.0591141, 0.04693888, 0.03369704, 0.01935668, 0.009381749, 0.006103575, 
    0.009275854, 0.01864177, 0.03425273, 0.04759809, 0.0554316, 0.06400007, 
    0.07673949, 0.09488726, 0.1146543, 0.1318182, 0.1474278, 0.154835, 
    0.1460786, 0.129799, 0.1156039, 0.09906316, 0.08267778, 0.06752437, 
    0.04845288, 0.02746509, 0.009031892, -0.005337708, -0.01690768, 
    -0.02574366, -0.03043796, -0.02933829, -0.0254358, -0.0221101, 
    -0.01582015, -0.005312525, 0.006336138, 0.01931216, 0.03186979, 
    0.04390969, 0.05540673, 0.0655934, 0.07564066, 0.08287154, 0.08376838, 
    0.08074595, 0.07812048, 0.07322165, 0.0632641, 0.05173298, 0.03738473, 
    0.01922539, 0.0001538331, -0.01933139, -0.03951796, -0.06047678, 
    -0.08084124, -0.1004149, -0.118575, -0.1360216, -0.1540258, -0.1726229, 
    -0.1900944, -0.2051539, -0.2176192, -0.2260481, -0.2308431, -0.2327951, 
    -0.2314097, -0.2277237, -0.2228221,
  -0.2165065, -0.2091498, -0.1994938, -0.1897301, -0.1796337, -0.1666086, 
    -0.1519695, -0.136151, -0.1205062, -0.1056692, -0.09013789, -0.07536903, 
    -0.06002931, -0.04320132, -0.02574639, -0.008201439, 0.008796999, 
    0.02366571, 0.03670103, 0.04810885, 0.0579503, 0.06552502, 0.07114039, 
    0.07727053, 0.08536169, 0.09512491, 0.10443, 0.1076791, 0.1067826, 
    0.1044131, 0.09944968, 0.0916604, 0.08244286, 0.07226601, 0.05615667, 
    0.03551763, 0.01851614, 0.008212775, 0.0005726814, -0.007632598, 
    -0.01408479, -0.01925381, -0.03041756, -0.0495621, -0.06502718, 
    -0.07095757, -0.06851193, -0.05859455, -0.04470418, -0.02914253, 
    -0.0148956, -0.004766956, 0.001169011, 0.002054557, 8.247048e-05, 
    -0.0005640909, -0.0004211217, -0.002393976, -0.006794222, -0.01180337, 
    -0.01549035, -0.02045619, -0.0274362, -0.03259332, -0.03286166, 
    -0.02448195, -0.004081905, 0.02329767, 0.04776651, 0.07388496, 0.1000131, 
    0.1210891, 0.1389601, 0.145692, 0.1366978, 0.1266816, 0.1249099, 
    0.1247856, 0.1175472, 0.1013259, 0.08156486, 0.0616833, 0.0406679, 
    0.02160874, 0.006559178, -0.005917519, -0.01579891, -0.02396424, 
    -0.03356467, -0.03980687, -0.03390759, -0.01705059, 0.002112895, 
    0.01782018, 0.03160631, 0.04329471, 0.05354637, 0.0634125, 0.07140711, 
    0.07718669, 0.08099188, 0.08372244, 0.08596054, 0.08406036, 0.0770914, 
    0.06744553, 0.05446941, 0.03872152, 0.02159896, 0.002792634, -0.01741427, 
    -0.03838722, -0.06012045, -0.08143714, -0.1005423, -0.1179334, 
    -0.1348706, -0.1524424, -0.1705506, -0.188056, -0.2038801, -0.2159065, 
    -0.2242536, -0.2292326, -0.2309861, -0.2295242, -0.2258812, -0.2215575,
  -0.2141691, -0.2067741, -0.1973436, -0.1875048, -0.1769537, -0.1632734, 
    -0.1489461, -0.1341303, -0.1173854, -0.1012785, -0.08687446, -0.07242098, 
    -0.05658523, -0.04028718, -0.02286742, -0.004922934, 0.0112426, 
    0.02552353, 0.03835009, 0.04938477, 0.05896648, 0.0669686, 0.0748295, 
    0.08463322, 0.09319291, 0.09789152, 0.1028345, 0.110628, 0.1191411, 
    0.1190844, 0.1071871, 0.09500502, 0.08813761, 0.08139165, 0.07024685, 
    0.05246612, 0.03142634, 0.01528251, 0.00671494, 0.001066506, 
    -0.006744951, -0.01405481, -0.02133116, -0.03094208, -0.04266816, 
    -0.0575422, -0.07174918, -0.08268809, -0.08976066, -0.09495321, 
    -0.09795479, -0.09851177, -0.0960414, -0.09211673, -0.08853416, 
    -0.08589092, -0.08326454, -0.07994875, -0.07720307, -0.0769757, 
    -0.08060262, -0.08570982, -0.08889327, -0.08605081, -0.07315738, 
    -0.04663122, -0.01383497, 0.01866537, 0.05140972, 0.08140045, 0.104067, 
    0.1205837, 0.1324574, 0.1365129, 0.1390802, 0.1472319, 0.1471791, 
    0.1325855, 0.1108806, 0.08921623, 0.06839162, 0.04639298, 0.02556258, 
    0.007617644, -0.006482638, -0.01707975, -0.0242689, -0.02742842, 
    -0.02594316, -0.02259384, -0.01980583, -0.0136895, -0.003076404, 
    0.008585557, 0.0215213, 0.03447934, 0.04668577, 0.05813104, 0.06799179, 
    0.07702414, 0.08413853, 0.08656426, 0.08515674, 0.08200255, 0.07561634, 
    0.06599867, 0.05491757, 0.04071352, 0.0233496, 0.004471038, -0.01505812, 
    -0.03549537, -0.05679705, -0.07747164, -0.09705189, -0.1155039, 
    -0.1335132, -0.1515685, -0.1702402, -0.1879733, -0.2032038, -0.2158944, 
    -0.2246791, -0.2295837, -0.231268, -0.2295592, -0.225478, -0.2201085,
  -0.213854, -0.2061846, -0.1960325, -0.1853956, -0.1741118, -0.1601656, 
    -0.1453352, -0.1296903, -0.1139871, -0.09871245, -0.08301537, 
    -0.06836338, -0.05352179, -0.03705478, -0.01961499, -0.002465621, 
    0.0137422, 0.02820012, 0.04090409, 0.05180617, 0.06079827, 0.06745789, 
    0.07297578, 0.0803751, 0.08979283, 0.09862325, 0.103628, 0.104337, 
    0.1036299, 0.0999947, 0.09518217, 0.09372076, 0.08997606, 0.07986553, 
    0.06415614, 0.04264045, 0.02352402, 0.01332065, 0.006713688, 
    -0.0002976954, -0.007529974, -0.01297736, -0.01850647, -0.02567133, 
    -0.03398716, -0.04510501, -0.05745202, -0.06886181, -0.08271766, 
    -0.09803301, -0.1057045, -0.1113223, -0.1172279, -0.1213248, -0.1229584, 
    -0.1211604, -0.1169109, -0.1123111, -0.1083243, -0.1037241, -0.09844739, 
    -0.09589682, -0.09317894, -0.08283765, -0.06723984, -0.04567519, 
    -0.01217698, 0.02742034, 0.0586679, 0.08376026, 0.105613, 0.1234807, 
    0.1373891, 0.1459757, 0.1501166, 0.1430004, 0.125724, 0.1131271, 
    0.1034304, 0.08905739, 0.07314527, 0.05765027, 0.04058743, 0.02368582, 
    0.008610904, -0.004783541, -0.01578978, -0.0249805, -0.03495818, 
    -0.04040664, -0.03292668, -0.01494357, 0.004511893, 0.02044681, 
    0.0344824, 0.04632045, 0.05653798, 0.06627749, 0.07442348, 0.0801513, 
    0.08401146, 0.08714779, 0.08881912, 0.08550664, 0.07895524, 0.07122663, 
    0.05875162, 0.0425145, 0.02508235, 0.006495275, -0.01335164, -0.03447988, 
    -0.05656966, -0.07810974, -0.09744443, -0.1155891, -0.133269, -0.1511502, 
    -0.1692728, -0.1869625, -0.2032187, -0.2157405, -0.224209, -0.2288992, 
    -0.2304311, -0.2288357, -0.2246765, -0.2195442,
  -0.2126213, -0.2046098, -0.1946795, -0.1842317, -0.1726283, -0.1580748, 
    -0.143635, -0.1289665, -0.1119455, -0.0952407, -0.08081309, -0.06681724, 
    -0.05105225, -0.03436623, -0.0172032, -0.0001188815, 0.01598365, 
    0.0305696, 0.04261619, 0.052725, 0.06260866, 0.07125079, 0.0787362, 
    0.08704555, 0.09477867, 0.1008894, 0.1058116, 0.109554, 0.1115576, 
    0.1089866, 0.1029203, 0.09577967, 0.08754204, 0.07995921, 0.07058863, 
    0.05559829, 0.03955805, 0.02715677, 0.01879206, 0.01232761, 0.003425479, 
    -0.006613821, -0.01499933, -0.02014658, -0.02296093, -0.02908263, 
    -0.03993982, -0.05601093, -0.07603934, -0.09859678, -0.1123551, 
    -0.117188, -0.1192092, -0.1193694, -0.1189308, -0.1167612, -0.1122229, 
    -0.1055825, -0.09883358, -0.09149942, -0.08419999, -0.08118294, 
    -0.08213717, -0.07696395, -0.06243717, -0.03538629, -2.1182e-05, 
    0.03445557, 0.06625453, 0.09179509, 0.1101347, 0.1266969, 0.1382853, 
    0.1406455, 0.1364523, 0.1323654, 0.132295, 0.1301221, 0.117651, 
    0.09868777, 0.07675529, 0.05287075, 0.02985382, 0.009069651, 
    -0.006500185, -0.01689062, -0.02272633, -0.02424082, -0.02234861, 
    -0.01971805, -0.01768723, -0.01185676, -0.001309127, 0.01030868, 
    0.02352296, 0.03700072, 0.04944207, 0.06057805, 0.07031619, 0.07967959, 
    0.08687991, 0.08886987, 0.08719382, 0.08452819, 0.07903286, 0.06939327, 
    0.05784393, 0.04417435, 0.02774835, 0.008913912, -0.01114374, 
    -0.03168703, -0.05325891, -0.0747676, -0.09492431, -0.1135537, 
    -0.1321179, -0.150927, -0.1699192, -0.1877227, -0.2030744, -0.216049, 
    -0.2252001, -0.2301705, -0.2314262, -0.2292284, -0.2248356, -0.2191305,
  -0.2130156, -0.204666, -0.193917, -0.1827852, -0.1708229, -0.1561852, 
    -0.1410643, -0.1254115, -0.1095101, -0.09386314, -0.07802093, 
    -0.06344695, -0.04876428, -0.03230342, -0.01484928, 0.002060529, 
    0.01808507, 0.03225246, 0.04411945, 0.05429052, 0.06307197, 0.06974263, 
    0.076106, 0.08468315, 0.09364799, 0.1004275, 0.1050575, 0.1095377, 
    0.1128846, 0.111502, 0.1064688, 0.1001817, 0.09331933, 0.08503897, 
    0.0706839, 0.04914135, 0.02941528, 0.01746666, 0.00977084, 0.003145337, 
    -0.002615124, -0.008220106, -0.01618725, -0.02464151, -0.02778161, 
    -0.02900943, -0.03408703, -0.04451886, -0.05850005, -0.08074954, 
    -0.1033579, -0.115716, -0.1210344, -0.122844, -0.1226795, -0.1191709, 
    -0.1120745, -0.103504, -0.09579681, -0.08769567, -0.07744606, 
    -0.07220563, -0.07116285, -0.06142802, -0.04445063, -0.02204828, 
    0.0104878, 0.04678117, 0.07364845, 0.09364033, 0.109864, 0.1223697, 
    0.1319206, 0.1380628, 0.1431402, 0.1438884, 0.1354264, 0.1207852, 
    0.1026495, 0.08299065, 0.06586635, 0.05044049, 0.03462645, 0.02113664, 
    0.009065083, -0.004024558, -0.0159705, -0.02601364, -0.03607097, 
    -0.04059082, -0.0318321, -0.0127328, 0.007471859, 0.02355665, 0.03736314, 
    0.04918104, 0.05967456, 0.06959979, 0.07758407, 0.08309375, 0.08684243, 
    0.08956479, 0.09133075, 0.08902352, 0.08269332, 0.07441206, 0.06251144, 
    0.04753166, 0.03010999, 0.01053719, -0.009396121, -0.02998785, 
    -0.05243034, -0.07496893, -0.09499512, -0.1135933, -0.1319357, 
    -0.1504653, -0.1691432, -0.1873829, -0.2038551, -0.2164541, -0.2252678, 
    -0.2301778, -0.2314353, -0.2292937, -0.2246969, -0.219227,
  -0.2124209, -0.2039422, -0.1932301, -0.1821155, -0.1700351, -0.1550262, 
    -0.1401494, -0.1252443, -0.1081741, -0.09120601, -0.07638086, -0.0623709, 
    -0.04689258, -0.03015589, -0.01273767, 0.00431022, 0.02007131, 
    0.03414705, 0.04599561, 0.05633378, 0.06599337, 0.07384391, 0.08076324, 
    0.08842029, 0.09578517, 0.101822, 0.1059294, 0.1088065, 0.1091708, 
    0.1048632, 0.09836575, 0.09263393, 0.08721107, 0.08058788, 0.07086593, 
    0.05665204, 0.04216796, 0.03190947, 0.02573645, 0.01942423, 0.009398401, 
    -0.001289994, -0.01062387, -0.01811031, -0.02087626, -0.02245161, 
    -0.02650553, -0.03651106, -0.05309564, -0.07820332, -0.1021738, 
    -0.115113, -0.1194197, -0.1188583, -0.1169302, -0.1134111, -0.1066797, 
    -0.0972323, -0.08740285, -0.07722597, -0.06740162, -0.06194103, 
    -0.0586074, -0.04952333, -0.03418921, -0.007866696, 0.02415081, 
    0.05260335, 0.0779354, 0.09857594, 0.1130528, 0.1249747, 0.1349, 
    0.1412039, 0.1412341, 0.1349911, 0.1269389, 0.1202681, 0.1114315, 
    0.09944785, 0.08205962, 0.05951566, 0.03669339, 0.01452479, -0.003426872, 
    -0.01517043, -0.0207305, -0.02134818, -0.01903364, -0.01675233, 
    -0.01554835, -0.01040676, 0.000133276, 0.01218212, 0.02572203, 
    0.03942963, 0.05206889, 0.06336892, 0.07297178, 0.08179498, 0.08936432, 
    0.09223062, 0.09038678, 0.08744313, 0.08271143, 0.07387188, 0.0624125, 
    0.04862633, 0.03263509, 0.01455209, -0.00568226, -0.02723753, 
    -0.04932075, -0.07108365, -0.09201041, -0.1116677, -0.1311536, 
    -0.1505512, -0.1698949, -0.188203, -0.2040998, -0.2172973, -0.2265416, 
    -0.2316658, -0.2328772, -0.2302758, -0.2252584, -0.2191488,
  -0.2131878, -0.2043508, -0.1930715, -0.1813558, -0.1687875, -0.1536909, 
    -0.1383781, -0.1225223, -0.1061604, -0.09019928, -0.07446764, 
    -0.05997035, -0.04504878, -0.02834874, -0.01104299, 0.005655646, 
    0.02175057, 0.03565578, 0.04673764, 0.0565566, 0.06566809, 0.0730079, 
    0.07994418, 0.08781498, 0.09534675, 0.1016516, 0.1064185, 0.1105497, 
    0.1123841, 0.1104037, 0.1070264, 0.1028276, 0.09615348, 0.08705491, 
    0.07338956, 0.0533644, 0.03403458, 0.02091599, 0.01171911, 0.004413992, 
    -0.00121215, -0.006703138, -0.01533756, -0.02513096, -0.0285106, 
    -0.02750775, -0.02886245, -0.03550687, -0.04796517, -0.07024208, 
    -0.0949692, -0.1113823, -0.1185607, -0.1197819, -0.1181842, -0.1129826, 
    -0.1041359, -0.09375744, -0.08345431, -0.07265131, -0.06214243, 
    -0.05654685, -0.05107918, -0.03811495, -0.02015308, 0.002582353, 
    0.03137098, 0.06158207, 0.08277892, 0.0980185, 0.1121653, 0.1238738, 
    0.1323861, 0.1365288, 0.1375109, 0.1363635, 0.1337109, 0.1271622, 
    0.1102573, 0.08622643, 0.06427884, 0.04589194, 0.0286974, 0.01556349, 
    0.005892038, -0.004993502, -0.01626639, -0.02661544, -0.03677416, 
    -0.0402635, -0.0298965, -0.009568721, 0.01110727, 0.02709389, 0.04056999, 
    0.05242002, 0.06309617, 0.07292566, 0.08104649, 0.08656287, 0.09018266, 
    0.09304476, 0.09481674, 0.09281284, 0.08728416, 0.07951708, 0.06762006, 
    0.05289581, 0.03631052, 0.01691001, -0.003752895, -0.02453991, 
    -0.04698344, -0.07054126, -0.09183624, -0.1111327, -0.1303114, 
    -0.1500029, -0.1694267, -0.1881673, -0.205173, -0.2181653, -0.2272301, 
    -0.232196, -0.2332987, -0.2308754, -0.2258627, -0.2199085,
  -0.2449929, -0.2392884, -0.2324482, -0.2240469, -0.2143291, -0.202827, 
    -0.1888396, -0.173116, -0.1547283, -0.133271, -0.1105209, -0.08933939, 
    -0.06877743, -0.04836127, -0.02835062, -0.01034009, 0.005295783, 
    0.01846017, 0.03098533, 0.04326922, 0.05442377, 0.0638371, 0.07141474, 
    0.0767365, 0.08270966, 0.08853684, 0.09443625, 0.09826045, 0.09577654, 
    0.09130248, 0.09004989, 0.08962412, 0.08818743, 0.08719844, 0.08573461, 
    0.08178321, 0.07489228, 0.06834906, 0.06320795, 0.05421805, 0.0423921, 
    0.03257495, 0.0244329, 0.0159958, 0.006407201, -0.004754871, -0.01720938, 
    -0.03034914, -0.04368502, -0.05702665, -0.0698944, -0.08340666, 
    -0.0973624, -0.1097644, -0.1170023, -0.1187208, -0.1214039, -0.1249546, 
    -0.1083063, -0.07124652, -0.03709273, -0.02111065, -0.03886221, 
    -0.09789464, -0.168264, -0.2054659, -0.1992757, -0.1666826, -0.1286623, 
    -0.06154938, 0.05634288, 0.1149195, 0.1057072, 0.122903, 0.136345, 
    0.144941, 0.1546072, 0.1551152, 0.1546813, 0.1509999, 0.1418307, 
    0.1252345, 0.1044551, 0.08383954, 0.06492504, 0.04806867, 0.03207666, 
    0.01179975, -0.006366894, -0.02076851, -0.02784687, -0.02267939, 
    -0.01580304, -0.01369786, -0.01300824, -0.01111984, -0.006981909, 
    -0.0008651018, 0.006618023, 0.01664984, 0.02901834, 0.0424763, 
    0.05546892, 0.06680381, 0.07877359, 0.09032345, 0.09510216, 0.09249464, 
    0.0880582, 0.08268877, 0.07308131, 0.05890746, 0.04165544, 0.02136502, 
    -0.003093064, -0.02972931, -0.05453542, -0.08189395, -0.1094573, 
    -0.1316266, -0.1536782, -0.1691314, -0.1846146, -0.2037138, -0.2229995, 
    -0.2374371, -0.2442036, -0.2470003,
  -0.2447772, -0.2406219, -0.2344304, -0.2269427, -0.2169771, -0.2039015, 
    -0.1882389, -0.1694666, -0.1496278, -0.1299099, -0.1099561, -0.08835271, 
    -0.0671756, -0.04692274, -0.02853858, -0.01138769, 0.004868835, 
    0.02026001, 0.03333704, 0.04398528, 0.05271474, 0.06060153, 0.06811708, 
    0.07672402, 0.0850203, 0.09240095, 0.09775789, 0.09894727, 0.09439534, 
    0.09152631, 0.0910663, 0.08959179, 0.08924764, 0.08882028, 0.08512092, 
    0.079312, 0.07453507, 0.07151473, 0.06426015, 0.05108273, 0.03989452, 
    0.03131515, 0.02349725, 0.01546699, 0.006444454, -0.004784942, 
    -0.01771179, -0.03136125, -0.04473907, -0.05853626, -0.07342261, 
    -0.08645609, -0.09589526, -0.1040635, -0.1133991, -0.1229614, -0.1282379, 
    -0.129954, -0.1281114, -0.1112542, -0.07670696, -0.0368527, 
    -0.0001826622, 0.0212121, 0.01646313, -0.00626304, -0.02152047, 
    -0.0100769, 0.03407839, 0.08477464, 0.09462152, 0.08559869, 0.1073282, 
    0.1276884, 0.1332995, 0.143929, 0.1520325, 0.1577222, 0.1578912, 
    0.1515793, 0.141403, 0.127368, 0.1094851, 0.08734921, 0.06331491, 
    0.03960091, 0.01942286, 0.007912755, -0.001016945, -0.008271128, 
    -0.0152523, -0.02535574, -0.0302439, -0.02742282, -0.02064604, 
    -0.01288846, -0.004318893, 0.00538373, 0.01517028, 0.0252319, 0.03432083, 
    0.04226702, 0.05070728, 0.06023857, 0.06728104, 0.07117602, 0.07720204, 
    0.08384673, 0.084558, 0.07999364, 0.0725497, 0.06052089, 0.04411483, 
    0.0230082, -0.001133174, -0.02738103, -0.05486608, -0.07919678, 
    -0.1034828, -0.1297088, -0.1502188, -0.1730434, -0.1949547, -0.210741, 
    -0.2219168, -0.2319586, -0.2413409, -0.2454314,
  -0.2453417, -0.2392756, -0.2320976, -0.2233599, -0.2132018, -0.2011405, 
    -0.1866015, -0.1703886, -0.1517451, -0.1301548, -0.1073971, -0.08615965, 
    -0.06565788, -0.04521942, -0.02519363, -0.006993741, 0.008709729, 
    0.02165255, 0.03329211, 0.04446708, 0.05530903, 0.06592587, 0.07510237, 
    0.08087204, 0.08606692, 0.09132504, 0.09675866, 0.09977803, 0.09700829, 
    0.09274282, 0.09102044, 0.08930311, 0.08663598, 0.08579049, 0.08564806, 
    0.08293673, 0.07626894, 0.06942484, 0.06397456, 0.05426013, 0.04107291, 
    0.03029716, 0.02185872, 0.01313201, 0.003012598, -0.008407623, 
    -0.02087158, -0.03381452, -0.04704198, -0.06037433, -0.07313384, 
    -0.08621487, -0.09948403, -0.1103155, -0.1157963, -0.1175561, -0.1183363, 
    -0.1190295, -0.1192089, -0.1198066, -0.1144863, -0.09770383, -0.07170298, 
    -0.03956002, -0.006007366, 0.02316862, 0.04393873, 0.0562295, 0.05768666, 
    0.05412461, 0.06580131, 0.09172137, 0.1104431, 0.122312, 0.1343508, 
    0.1452631, 0.1541071, 0.1573725, 0.1565317, 0.1521886, 0.1426125, 0.1267, 
    0.1070026, 0.0878104, 0.06909931, 0.05040389, 0.03110623, 0.009099633, 
    -0.007692665, -0.01829663, -0.02185546, -0.01614508, -0.01115504, 
    -0.01079109, -0.01072519, -0.008526176, -0.003695071, 0.003008425, 
    0.01094502, 0.02128989, 0.03391629, 0.04793096, 0.06153515, 0.07343927, 
    0.08707246, 0.1010977, 0.1063925, 0.1036905, 0.09994596, 0.09118536, 
    0.07311104, 0.05174839, 0.03324664, 0.01764238, -0.0001631379, 
    -0.02405569, -0.05140594, -0.07953957, -0.1045554, -0.1273281, 
    -0.1511923, -0.1672467, -0.1842388, -0.2041812, -0.2235589, -0.2378506, 
    -0.2446014, -0.2474596,
  -0.2454558, -0.2411367, -0.2345949, -0.226649, -0.2161757, -0.2027175, 
    -0.1866567, -0.1675788, -0.1473235, -0.1272923, -0.1071126, -0.08546969, 
    -0.06422955, -0.04403031, -0.02579004, -0.008987054, 0.006819338, 
    0.0219613, 0.03536133, 0.04689623, 0.05644382, 0.06393156, 0.06984511, 
    0.07739935, 0.08605675, 0.09386085, 0.09897599, 0.0998096, 0.09505114, 
    0.09180366, 0.09121165, 0.09046045, 0.09120601, 0.0903213, 0.08358836, 
    0.07425514, 0.06772077, 0.06483749, 0.05786963, 0.0455845, 0.03604691, 
    0.02779996, 0.01978247, 0.01190066, 0.00254029, -0.009534098, 
    -0.02345168, -0.03767157, -0.05084928, -0.06399543, -0.07813478, 
    -0.09033781, -0.09898441, -0.1066387, -0.1147508, -0.1220691, -0.12579, 
    -0.1243066, -0.1178113, -0.1083336, -0.0987339, -0.08966181, -0.07753277, 
    -0.06275409, -0.04634368, -0.02974782, -0.01400301, 0.002360821, 
    0.0260818, 0.05442095, 0.07487491, 0.08835047, 0.1061665, 0.1250411, 
    0.1347388, 0.1443806, 0.1531555, 0.1572687, 0.1572841, 0.1518111, 
    0.1421914, 0.1278651, 0.1090604, 0.08603702, 0.0627979, 0.04181974, 
    0.0246029, 0.01352453, 0.002111524, -0.008738399, -0.01760945, 
    -0.02616815, -0.02777546, -0.02266591, -0.01503117, -0.007144004, 
    0.001311138, 0.01094225, 0.02101681, 0.03147817, 0.04094239, 0.04912302, 
    0.05802438, 0.06876564, 0.07563051, 0.07647838, 0.08281662, 0.0904949, 
    0.07866837, 0.05542372, 0.04198578, 0.03565639, 0.02312955, 0.0003244877, 
    -0.02179132, -0.03453387, -0.04773675, -0.07225904, -0.1006861, 
    -0.1249397, -0.1466052, -0.1714676, -0.1936144, -0.210275, -0.2219173, 
    -0.2326195, -0.2422985, -0.2463449,
  -0.2461347, -0.2395985, -0.2321798, -0.2231718, -0.2126026, -0.1999646, 
    -0.1849571, -0.1683359, -0.149474, -0.1277402, -0.104887, -0.08356407, 
    -0.06309015, -0.04272434, -0.02267629, -0.004311681, 0.011712, 
    0.02494368, 0.03656586, 0.04710206, 0.05684859, 0.06682271, 0.07685743, 
    0.08414292, 0.08966848, 0.0945972, 0.1001572, 0.1026165, 0.09876484, 
    0.09436435, 0.09212375, 0.08773994, 0.08090216, 0.07538265, 0.07364839, 
    0.07328364, 0.0692822, 0.06398614, 0.05711447, 0.04518366, 0.03212787, 
    0.02168921, 0.01258401, 0.003843844, -0.005293682, -0.01550072, 
    -0.02696882, -0.03972098, -0.05354958, -0.06719151, -0.07942968, 
    -0.09184201, -0.1041642, -0.1134626, -0.1176857, -0.1186667, -0.1185947, 
    -0.1192124, -0.1180227, -0.1136405, -0.1050181, -0.09257576, -0.07716464, 
    -0.05918726, -0.03984346, -0.01961744, 0.000585705, 0.01908147, 
    0.03360549, 0.04663831, 0.06520411, 0.0867933, 0.1073231, 0.1235873, 
    0.1341067, 0.1448903, 0.1544023, 0.159584, 0.1602198, 0.1559127, 
    0.1463029, 0.1304049, 0.1110564, 0.09177768, 0.0712743, 0.04968923, 
    0.0288374, 0.008235663, -0.004976556, -0.01208332, -0.01451803, 
    -0.01054634, -0.007891696, -0.008593763, -0.008262448, -0.005112924, 
    0.0007833764, 0.008155301, 0.01655955, 0.02722883, 0.04031599, 
    0.05518688, 0.06979707, 0.08130566, 0.09536937, 0.1177067, 0.1289059, 
    0.1054608, 0.08302367, 0.1073485, 0.1540509, 0.1826319, 0.179521, 
    0.1415489, 0.06966472, -0.0124191, -0.06073477, -0.07319051, -0.09387369, 
    -0.1235119, -0.1459896, -0.1641031, -0.1832681, -0.2041306, -0.2242559, 
    -0.2383848, -0.2453395, -0.2483419,
  -0.2465206, -0.2421219, -0.2351868, -0.2266372, -0.2157341, -0.2019426, 
    -0.1855692, -0.1661054, -0.1454696, -0.1251039, -0.1047659, -0.08301964, 
    -0.06169549, -0.04137501, -0.02314079, -0.006496698, 0.008900404, 
    0.02362418, 0.0367054, 0.04836431, 0.05875566, 0.06734554, 0.07324139, 
    0.07949027, 0.08739969, 0.09561731, 0.09958237, 0.09855588, 0.09375851, 
    0.08914405, 0.08277065, 0.07727636, 0.08002573, 0.08628571, 0.08799876, 
    0.0845056, 0.08194237, 0.0811119, 0.07227049, 0.05399724, 0.03485209, 
    0.01985581, 0.007552013, -0.003739923, -0.0148403, -0.02713472, 
    -0.0393047, -0.05048423, -0.06111995, -0.07269187, -0.08593079, 
    -0.0970448, -0.1045112, -0.1111911, -0.1182578, -0.124033, -0.125941, 
    -0.1227246, -0.1160546, -0.1080232, -0.09936082, -0.09039295, 
    -0.07917754, -0.0658943, -0.05056366, -0.03487309, -0.01989958, 
    -0.004065186, 0.01848599, 0.04480866, 0.06630147, 0.08486871, 0.1055999, 
    0.1241271, 0.1350525, 0.146549, 0.1562693, 0.1594838, 0.1584297, 
    0.1530689, 0.1435098, 0.1291009, 0.1102931, 0.08760057, 0.06582531, 
    0.04636514, 0.0288846, 0.01529616, 0.0008408129, -0.01133912, 
    -0.01849268, -0.02339939, -0.02175596, -0.01524498, -0.007545784, 
    -4.481524e-05, 0.008164109, 0.01780593, 0.02827305, 0.03898885, 
    0.0485358, 0.05651488, 0.06544868, 0.07882787, 0.09204325, 0.08802948, 
    0.06461087, 0.06690387, 0.1379315, 0.2346287, 0.2929218, 0.3100459, 
    0.3089161, 0.2974437, 0.2618256, 0.1745367, 0.03665427, -0.07001211, 
    -0.09354371, -0.1125407, -0.1430418, -0.1665493, -0.1917271, -0.2091187, 
    -0.2218305, -0.2332524, -0.2433334, -0.2473146,
  -0.2466018, -0.2399339, -0.2322349, -0.2232798, -0.212105, -0.1990263, 
    -0.183458, -0.1666151, -0.1474692, -0.1256937, -0.1026292, -0.08129311, 
    -0.06077611, -0.04060382, -0.02057478, -0.00226894, 0.0140194, 
    0.02749139, 0.03949638, 0.05013871, 0.05952729, 0.06826018, 0.077724, 
    0.08602433, 0.09326267, 0.09728985, 0.1021317, 0.1055772, 0.09890512, 
    0.08932355, 0.08613934, 0.087352, 0.08588132, 0.07595006, 0.06368195, 
    0.05493739, 0.05055859, 0.0568716, 0.07257634, 0.06855705, 0.04635212, 
    0.03320948, 0.02253036, 0.00779623, -0.007729938, -0.02376323, 
    -0.03949037, -0.05444266, -0.06778959, -0.07926202, -0.09000565, 
    -0.101531, -0.1122685, -0.1196081, -0.1225122, -0.1224964, -0.1222404, 
    -0.1223156, -0.1201665, -0.1145018, -0.1056214, -0.09403554, -0.08041325, 
    -0.06551438, -0.04992849, -0.03275822, -0.01381554, 0.004997522, 
    0.02208216, 0.03950854, 0.06131279, 0.08342618, 0.1050258, 0.1242985, 
    0.135514, 0.1451228, 0.1544241, 0.1610636, 0.1639746, 0.1603818, 
    0.1508546, 0.1346834, 0.1142631, 0.09305309, 0.07058376, 0.04831835, 
    0.02907299, 0.01123223, 0.0003303587, -0.006616272, -0.01114423, 
    -0.009825855, -0.008179992, -0.007893205, -0.005751319, -0.000979729, 
    0.006020553, 0.01393541, 0.02274782, 0.03395399, 0.04809967, 0.06501797, 
    0.08295251, 0.09647401, 0.1028889, 0.1047602, 0.1160809, 0.1693553, 
    0.2641913, 0.3338807, 0.3507873, 0.3433163, 0.3278605, 0.3111934, 
    0.3021138, 0.2858846, 0.2217205, 0.06429958, -0.08348075, -0.1130326, 
    -0.1343483, -0.1607832, -0.1791329, -0.2041995, -0.224023, -0.239114, 
    -0.2457991, -0.2495497,
  -0.2477368, -0.2430526, -0.2354984, -0.2263794, -0.2151787, -0.2011819, 
    -0.1844615, -0.1646672, -0.1436588, -0.1230554, -0.1025702, -0.08078343, 
    -0.05932778, -0.0388709, -0.02048188, -0.003835559, 0.01143771, 
    0.02592623, 0.03877461, 0.05012058, 0.06052923, 0.06997669, 0.07701887, 
    0.08319552, 0.08887866, 0.09579626, 0.1003696, 0.09202322, 0.07966027, 
    0.07794949, 0.07487705, 0.06680423, 0.05872059, 0.05745216, 0.06364742, 
    0.05996992, 0.03558532, 0.01755209, 0.02761335, 0.04664815, 0.04781229, 
    0.02435047, -0.003488857, -0.02318571, -0.03517336, -0.04603926, 
    -0.05716417, -0.0688903, -0.07904798, -0.09041771, -0.1015367, 
    -0.1093003, -0.1143843, -0.1207213, -0.1271372, -0.1305563, -0.1314643, 
    -0.1269781, -0.1206083, -0.1128328, -0.1048842, -0.09614085, -0.08541301, 
    -0.07208569, -0.05655903, -0.04066184, -0.02605355, -0.01044956, 
    0.01147245, 0.03743348, 0.05950794, 0.0805617, 0.1037013, 0.1235634, 
    0.1345594, 0.1485205, 0.161331, 0.1655371, 0.1635661, 0.1577878, 
    0.1481903, 0.1336249, 0.1139479, 0.09164967, 0.06986648, 0.04951769, 
    0.0303764, 0.01653068, 0.00239259, -0.007438891, -0.01173609, 
    -0.01324127, -0.009826303, -0.00320147, 0.0027242, 0.009381138, 
    0.01747818, 0.02828184, 0.0390748, 0.04948803, 0.05717904, 0.06300367, 
    0.06716362, 0.0738336, 0.08239617, 0.09521469, 0.1204518, 0.1810701, 
    0.2611314, 0.3217078, 0.3569598, 0.3799284, 0.3658096, 0.3192177, 
    0.2875405, 0.2748573, 0.2578236, 0.2094045, 0.04169121, -0.1082073, 
    -0.127673, -0.1601318, -0.1876998, -0.2068217, -0.2214057, -0.2336712, 
    -0.2439812, -0.2479709,
  -0.246994, -0.2393537, -0.232703, -0.2226862, -0.2115992, -0.1973127, 
    -0.1820453, -0.1644034, -0.1456489, -0.1232803, -0.1005781, -0.07871872, 
    -0.05868489, -0.03824192, -0.01878384, -0.0002170503, 0.0156858, 
    0.02962232, 0.04135562, 0.05257446, 0.0618829, 0.07068972, 0.07891582, 
    0.08685072, 0.09422334, 0.09985615, 0.09908501, 0.1003651, 0.1047734, 
    0.09230666, 0.06870526, 0.06475285, 0.0815164, 0.1179855, 0.1471738, 
    0.1413622, 0.07897297, 0.002322793, 0.001214519, 0.02333895, 
    -0.004324369, -0.03561209, -0.04356686, -0.04792742, -0.05434695, 
    -0.06336308, -0.0738005, -0.08640482, -0.0979518, -0.1090702, -0.1179233, 
    -0.1279798, -0.135546, -0.1394568, -0.1399702, -0.1370952, -0.1375715, 
    -0.135893, -0.1341231, -0.1268074, -0.1183377, -0.1055513, -0.09221365, 
    -0.07727969, -0.06309089, -0.04612924, -0.02736692, -0.007618323, 
    0.01003888, 0.03001505, 0.05383107, 0.07779166, 0.1008287, 0.1246739, 
    0.1381343, 0.1478341, 0.1554016, 0.1621149, 0.166018, 0.1639329, 
    0.1543994, 0.1380934, 0.1163794, 0.09564959, 0.07386907, 0.0541201, 
    0.03685754, 0.02000004, 0.007899113, -0.0007566176, -0.006909002, 
    -0.005921952, -0.004424207, -0.002701625, 0.001768477, 0.008744933, 
    0.01444769, 0.0190265, 0.02380196, 0.03451092, 0.05018723, 0.07088535, 
    0.09168248, 0.1109235, 0.1275707, 0.1476516, 0.1748315, 0.2053285, 
    0.2421511, 0.2792203, 0.3063109, 0.3007148, 0.2626124, 0.2175127, 
    0.1962272, 0.2095537, 0.2313119, 0.2179799, 0.1601291, -0.02988261, 
    -0.1337926, -0.1444213, -0.1783674, -0.1999301, -0.2250351, -0.2378644, 
    -0.2474372, -0.2493671,
  -0.2487018, -0.2427768, -0.2349681, -0.2252234, -0.2142941, -0.1997359, 
    -0.1829537, -0.1626081, -0.1416081, -0.1205988, -0.1003277, -0.07831466, 
    -0.05703884, -0.03622803, -0.01792541, -0.0009478927, 0.01414633, 
    0.02881414, 0.04146814, 0.05295763, 0.06310615, 0.07262085, 0.07985635, 
    0.08568317, 0.08968888, 0.0906316, 0.09045358, 0.09110498, 0.07189919, 
    0.05661188, 0.07544404, 0.1171742, 0.1550769, 0.1787839, 0.1702875, 
    0.1616342, 0.1235079, 0.01367362, -0.02290507, -0.02325805, -0.010844, 
    0.0174382, 0.02901369, 0.02116929, 0.004492626, -0.01720585, -0.04053176, 
    -0.06349382, -0.08500509, -0.1068098, -0.1259166, -0.1413552, -0.1517799, 
    -0.1612024, -0.1677009, -0.1675263, -0.1665533, -0.1571184, -0.1493708, 
    -0.1383282, -0.1304464, -0.1199995, -0.1095362, -0.09438655, -0.07631379, 
    -0.05809292, -0.04226714, -0.02609926, -0.002785653, 0.02437922, 
    0.04857677, 0.07212862, 0.09961173, 0.1228537, 0.1337352, 0.147644, 
    0.1655179, 0.17333, 0.1733917, 0.1673467, 0.1580307, 0.1411038, 
    0.1205629, 0.0970476, 0.07609141, 0.05469784, 0.03636919, 0.02075926, 
    0.007304676, -0.00277615, -0.005892605, -0.008461434, -0.003792448, 
    0.001424162, 0.005129928, 0.007124362, 0.0173282, 0.03591429, 0.06028139, 
    0.07493918, 0.07969591, 0.06709721, 0.05281763, 0.03028339, 0.02273193, 
    0.01091254, 0.006260678, 0.0122306, 0.01264593, 0.002560742, 
    -0.007111255, -0.0131867, -0.01035315, 0.006125636, 0.0485892, 
    0.09934958, 0.1516879, 0.167073, 0.1790219, 0.07658213, -0.1088234, 
    -0.148232, -0.1820948, -0.2036784, -0.2206169, -0.2334185, -0.2436307, 
    -0.2484079,
  -0.2448958, -0.2398185, -0.2311253, -0.2220462, -0.2088286, -0.1955992, 
    -0.1789737, -0.16232, -0.1424728, -0.1211122, -0.09741354, -0.07648739, 
    -0.05563086, -0.03625381, -0.01607198, 0.001437396, 0.01812109, 
    0.03114541, 0.04379759, 0.05421891, 0.06430314, 0.0717898, 0.07969426, 
    0.08494984, 0.09303603, 0.09783524, 0.1074897, 0.1009668, 0.06339105, 
    0.0754929, 0.1322253, 0.1567621, 0.1462054, 0.1289966, 0.1180302, 
    0.1328716, 0.1519564, 0.05555484, 0.01749353, 0.04928847, 0.08585401, 
    0.09156283, 0.07026337, 0.04725866, 0.02190004, -0.002491057, 
    -0.02759498, -0.05252964, -0.07635377, -0.09942813, -0.1229162, 
    -0.1473003, -0.1681462, -0.184804, -0.197242, -0.2059558, -0.21413, 
    -0.2158914, -0.2137634, -0.2012871, -0.1833465, -0.1588846, -0.1358051, 
    -0.1159865, -0.09843163, -0.07978505, -0.05566889, -0.03293693, 
    -0.01194599, 0.009964854, 0.03884232, 0.0653123, 0.09178764, 0.1207, 
    0.1408208, 0.1520912, 0.1621405, 0.1664277, 0.1707744, 0.1677075, 
    0.1602545, 0.1430426, 0.1238799, 0.1031932, 0.08191574, 0.05973652, 
    0.0404319, 0.01862988, 0.004405908, -0.006157093, -0.01062415, 
    -0.009638313, -0.01022557, -0.01178796, 0.002597237, 0.02897504, 
    0.05455896, 0.05310205, 0.02473541, -0.02483576, -0.06878913, -0.1086463, 
    -0.1317804, -0.1567928, -0.1716874, -0.190644, -0.2119576, -0.2120866, 
    -0.233533, -0.2360431, -0.2206586, -0.1956223, -0.1722226, -0.1354427, 
    -0.08491886, -0.02020107, 0.05945677, 0.1212703, 0.1311519, 0.1375846, 
    -0.04390371, -0.146049, -0.1642549, -0.2024552, -0.2199007, -0.2404617, 
    -0.2459816, -0.2497678,
  -0.246648, -0.2420876, -0.2321579, -0.2242641, -0.2113685, -0.1979187, 
    -0.1794492, -0.160365, -0.1380005, -0.1182055, -0.09687871, -0.07613644, 
    -0.05379924, -0.03403574, -0.01463112, 0.001354873, 0.01754448, 
    0.03132305, 0.04490231, 0.05506281, 0.06551188, 0.07365953, 0.08111391, 
    0.08725975, 0.09295972, 0.09508353, 0.09566487, 0.07092842, 0.06999796, 
    0.1283937, 0.1564875, 0.142301, 0.1337612, 0.128087, 0.1248001, 
    0.1105468, 0.1402803, 0.1217356, 0.1017131, 0.1454578, 0.1512397, 
    0.118597, 0.08726716, 0.06609088, 0.04664662, 0.02974491, 0.0134366, 
    -0.004286215, -0.02671276, -0.05125959, -0.07509516, -0.09417202, 
    -0.1103948, -0.1255558, -0.141368, -0.1576822, -0.1765315, -0.1949106, 
    -0.2140301, -0.2306975, -0.2402904, -0.2379252, -0.2190997, -0.1845582, 
    -0.1430137, -0.1101964, -0.08656366, -0.06574315, -0.03730479, 
    -0.004015148, 0.02423817, 0.05291438, 0.0854775, 0.1194791, 0.1349458, 
    0.1457009, 0.165307, 0.1778122, 0.1810166, 0.1778556, 0.1681467, 
    0.1501586, 0.1283122, 0.106883, 0.08347347, 0.06167831, 0.03868223, 
    0.02100136, 0.006473385, -0.0006712377, -0.006397642, -0.01281627, 
    -0.007777065, 0.02242221, 0.05446418, 0.05047355, -0.000342425, 
    -0.06628416, -0.1171018, -0.140867, -0.1524178, -0.1613177, -0.1742043, 
    -0.1893626, -0.2110353, -0.2318911, -0.2533062, -0.2646943, -0.2902281, 
    -0.2768915, -0.278068, -0.2806767, -0.2565385, -0.2046134, -0.1486844, 
    -0.08083535, -0.01353754, 0.05435215, 0.0775831, 0.1317156, 0.03612269, 
    -0.1374328, -0.1686831, -0.2051498, -0.2170578, -0.2334204, -0.2415253, 
    -0.2498067,
  -0.2438372, -0.237434, -0.2288517, -0.2182839, -0.2056273, -0.1917837, 
    -0.1755935, -0.158436, -0.1391604, -0.1175935, -0.09437779, -0.07321689, 
    -0.05290139, -0.03340012, -0.013724, 0.004062682, 0.02032924, 0.03348321, 
    0.04531638, 0.05585124, 0.06505474, 0.07217295, 0.0787724, 0.08532221, 
    0.09122835, 0.09946832, 0.09412478, 0.06183627, 0.09632219, 0.1554896, 
    0.1675133, 0.176091, 0.1696607, 0.1456316, 0.1381486, 0.1278189, 
    0.1222247, 0.1424233, 0.1667884, 0.2007779, 0.1939641, 0.151198, 
    0.118348, 0.1028314, 0.09170704, 0.08254701, 0.06954224, 0.05260146, 
    0.03169574, 0.01111275, -0.008638903, -0.02550867, -0.04072976, 
    -0.0560782, -0.07540208, -0.096692, -0.118597, -0.1391822, -0.1579597, 
    -0.1765997, -0.1980915, -0.2218227, -0.2446944, -0.2545963, -0.2410026, 
    -0.1983251, -0.1431248, -0.09437126, -0.06648663, -0.03535697, 
    0.0003221631, 0.03752974, 0.06716487, 0.1070288, 0.1370562, 0.1529168, 
    0.1682534, 0.1792212, 0.1827889, 0.1830112, 0.1732552, 0.1586346, 
    0.1354771, 0.1147136, 0.08853188, 0.06575703, 0.04273907, 0.02279857, 
    0.00925478, -0.001361609, -0.01213226, -0.003781185, 0.02667635, 
    0.05358705, 0.02181195, -0.05601782, -0.1247719, -0.1414071, -0.1381231, 
    -0.1414319, -0.1583515, -0.1737652, -0.1912244, -0.2108522, -0.234461, 
    -0.2513911, -0.2787622, -0.3051051, -0.3431784, -0.3572177, -0.3931509, 
    -0.3897721, -0.3458316, -0.2998231, -0.2385952, -0.1665367, -0.09893519, 
    -0.04334795, 0.01300254, 0.08879755, 0.07908262, -0.09992012, -0.1590937, 
    -0.195875, -0.2221211, -0.2390229, -0.2462851, -0.2470657,
  -0.2467426, -0.237446, -0.2310954, -0.2193999, -0.208646, -0.1923802, 
    -0.1763871, -0.1552812, -0.1350956, -0.1135594, -0.09441641, -0.07218987, 
    -0.05174318, -0.03033236, -0.01261297, 0.004911885, 0.01930494, 
    0.03449907, 0.04647386, 0.05761604, 0.06582062, 0.07592037, 0.08415937, 
    0.09477664, 0.1001386, 0.1074739, 0.1026695, 0.08095288, 0.1236925, 
    0.1771446, 0.1936271, 0.2028538, 0.202388, 0.1894216, 0.1585543, 
    0.1435399, 0.1390915, 0.1415114, 0.1477919, 0.1661193, 0.1739813, 
    0.1538039, 0.1317945, 0.1272734, 0.1214831, 0.1140279, 0.1000246, 
    0.0829141, 0.06160404, 0.04119615, 0.0199395, 0.001460999, -0.01984626, 
    -0.04298121, -0.07018192, -0.09680226, -0.1243381, -0.1469162, -0.165732, 
    -0.1772608, -0.1878261, -0.1962357, -0.2087584, -0.2235941, -0.2481465, 
    -0.2621415, -0.2516865, -0.1962993, -0.1329299, -0.07449299, -0.03621602, 
    0.004977748, 0.04637237, 0.09063689, 0.1296286, 0.1487732, 0.1645866, 
    0.1815268, 0.1866909, 0.1883792, 0.1805639, 0.1660294, 0.1435054, 
    0.1214132, 0.09561385, 0.06990082, 0.04635111, 0.02905517, 0.01293081, 
    -0.001642311, -0.004300203, 0.01856808, 0.04357067, 0.01492289, 
    -0.06271076, -0.1163889, -0.1234227, -0.1188427, -0.1308569, -0.1437037, 
    -0.1536514, -0.1573988, -0.1664648, -0.1778992, -0.1950731, -0.2166307, 
    -0.250131, -0.2865638, -0.3352616, -0.3763812, -0.4212013, -0.4204128, 
    -0.4018682, -0.3873102, -0.3200753, -0.2463525, -0.1600435, -0.07110574, 
    0.01373601, 0.05328654, 0.1030893, -0.0587132, -0.1654712, -0.1928136, 
    -0.2215104, -0.227461, -0.2433681, -0.2465866,
  -0.2427192, -0.2328288, -0.2263194, -0.2131879, -0.2029662, -0.1866356, 
    -0.1725713, -0.1535017, -0.1367028, -0.1135596, -0.09256443, -0.0697968, 
    -0.05158165, -0.03065485, -0.01294756, 0.006263265, 0.0206785, 
    0.03508351, 0.04470511, 0.05669524, 0.06658454, 0.07848648, 0.08524428, 
    0.08918826, 0.08685622, 0.08861415, 0.08048238, 0.07407831, 0.1314754, 
    0.1863889, 0.2018577, 0.22484, 0.2339505, 0.2318617, 0.2074981, 
    0.1658717, 0.1401216, 0.1472449, 0.1514823, 0.1432758, 0.1346913, 
    0.1376235, 0.1387156, 0.1397306, 0.1338819, 0.1269377, 0.1149654, 
    0.1025172, 0.08645444, 0.0689519, 0.04393606, 0.01655725, -0.0129932, 
    -0.03834265, -0.06415853, -0.08797929, -0.1156409, -0.1439936, 
    -0.1736504, -0.1955824, -0.2153503, -0.2297113, -0.2433763, -0.2443181, 
    -0.2460692, -0.2478611, -0.2663054, -0.2699969, -0.2479664, -0.1757588, 
    -0.09407823, -0.04062454, 0.002855472, 0.05192536, 0.1089119, 0.1467891, 
    0.1606103, 0.1820965, 0.1995316, 0.2011899, 0.1934636, 0.1764686, 
    0.1508818, 0.1269871, 0.1028533, 0.07726808, 0.05654427, 0.03452401, 
    0.01632092, 0.006274546, 0.01437987, 0.03652551, 0.01903476, -0.0628193, 
    -0.1387237, -0.1572822, -0.1428881, -0.1346841, -0.1267308, -0.1277345, 
    -0.1361468, -0.1411617, -0.1451098, -0.1512798, -0.1624319, -0.1772851, 
    -0.2048956, -0.2459876, -0.3058321, -0.3712365, -0.4371357, -0.4754556, 
    -0.502176, -0.4924546, -0.4242465, -0.3523575, -0.2461779, -0.1589735, 
    -0.05922641, -0.02789012, 0.07781921, -0.007435925, -0.1427691, 
    -0.1787167, -0.2245417, -0.2386475, -0.2468795, -0.2416069,
  -0.241943, -0.2346455, -0.2257191, -0.2149617, -0.202539, -0.1881092, 
    -0.1713358, -0.1517933, -0.1309279, -0.1107627, -0.09135327, -0.07024127, 
    -0.04944269, -0.02871285, -0.0107097, 0.006134942, 0.02064274, 
    0.03569001, 0.04911309, 0.06281134, 0.07338117, 0.08067939, 0.08241723, 
    0.08302638, 0.08166341, 0.08335219, 0.07866035, 0.07775424, 0.1335965, 
    0.1951066, 0.2161733, 0.233695, 0.2316, 0.2470491, 0.253878, 0.2224374, 
    0.1812949, 0.1493362, 0.1493421, 0.1682352, 0.1702843, 0.1692085, 
    0.1726795, 0.1695539, 0.1555014, 0.1407705, 0.1269272, 0.1173106, 
    0.1043918, 0.08584297, 0.05855861, 0.0305869, 0.0005245805, -0.0274021, 
    -0.05309339, -0.0767922, -0.1037321, -0.1300579, -0.1611918, -0.1918693, 
    -0.2207332, -0.2455767, -0.2696096, -0.2812312, -0.2867064, -0.282051, 
    -0.2814003, -0.2825111, -0.2912817, -0.2886392, -0.2282317, -0.1341291, 
    -0.05555513, 0.004675135, 0.0564678, 0.1155909, 0.1627222, 0.1850027, 
    0.1985825, 0.2074667, 0.206704, 0.1938633, 0.171526, 0.1416416, 
    0.1121624, 0.08635424, 0.06168241, 0.04180919, 0.01985503, 0.01275782, 
    0.02450929, 0.0261283, -0.02370416, -0.09442716, -0.1253876, -0.1244249, 
    -0.1104883, -0.1083407, -0.1186891, -0.1327364, -0.1307819, -0.1201262, 
    -0.1155962, -0.1125419, -0.1152128, -0.1245739, -0.1451936, -0.1763783, 
    -0.2313441, -0.308954, -0.391758, -0.4602851, -0.5129457, -0.5165736, 
    -0.4783963, -0.4064398, -0.3153177, -0.2097256, -0.1341808, -0.06504676, 
    0.08006363, 0.001972847, -0.1323209, -0.1732334, -0.203935, -0.2229246, 
    -0.2427439, -0.2482216,
  -0.248308, -0.2414196, -0.2319913, -0.2222353, -0.2092476, -0.1957103, 
    -0.1795022, -0.1636007, -0.1451689, -0.1250703, -0.1020525, -0.08199681, 
    -0.0619465, -0.04368465, -0.02386549, -0.006547213, 0.01109391, 
    0.02522574, 0.03895092, 0.04990537, 0.05836625, 0.06144483, 0.06671721, 
    0.06972186, 0.07024966, 0.06331715, 0.05445886, 0.06481743, 0.1236096, 
    0.1802292, 0.1988764, 0.2192032, 0.2369907, 0.2477252, 0.2403984, 
    0.2225416, 0.2294426, 0.2041533, 0.1503032, 0.1285029, 0.1486415, 
    0.1762166, 0.1880657, 0.1785197, 0.1671143, 0.1551477, 0.135934, 
    0.1191434, 0.1119597, 0.09862692, 0.07393961, 0.04382941, 0.01941985, 
    -0.005005687, -0.02921583, -0.05436918, -0.08218083, -0.1153406, 
    -0.1522789, -0.1945546, -0.232537, -0.2692107, -0.3044124, -0.3258291, 
    -0.3293979, -0.3247075, -0.3218255, -0.324919, -0.3165602, -0.3202641, 
    -0.3064468, -0.2810999, -0.2177276, -0.1211894, -0.03295393, 0.0345477, 
    0.1013023, 0.1566402, 0.1836904, 0.2032506, 0.2122341, 0.1995312, 
    0.1770072, 0.1486734, 0.1188388, 0.0893563, 0.06440336, 0.03798065, 
    0.01676271, 0.008503418, 0.01493223, 0.006434314, -0.06091013, 
    -0.1336768, -0.146503, -0.1446955, -0.1404369, -0.161593, -0.1617815, 
    -0.146966, -0.1435635, -0.1404335, -0.1338784, -0.1308517, -0.1276106, 
    -0.1203628, -0.1206121, -0.1382948, -0.1737147, -0.242112, -0.3326043, 
    -0.4222476, -0.5070776, -0.5638991, -0.5366979, -0.4994972, -0.4237877, 
    -0.308262, -0.1874184, -0.03947628, -0.00145144, -0.01370271, -0.1161277, 
    -0.1670982, -0.2088636, -0.2310225, -0.2372563, -0.2464547,
  -0.2687522, -0.2617192, -0.2598744, -0.2472263, -0.2411501, -0.2252873, 
    -0.2138871, -0.1928228, -0.1764401, -0.1547631, -0.1391671, -0.1165729, 
    -0.09830053, -0.0752344, -0.0581138, -0.03866863, -0.02475099, 
    -0.007888492, 0.00434123, 0.01811078, 0.02776494, 0.03948687, 0.04824976, 
    0.06457618, 0.07600547, 0.07229097, 0.0499503, 0.042889, 0.07425536, 
    0.1301776, 0.1663586, 0.1852827, 0.1927941, 0.2012497, 0.2003403, 
    0.1920771, 0.1944591, 0.1768112, 0.1364259, 0.1047127, 0.09632434, 
    0.1025011, 0.1175429, 0.1235508, 0.1350318, 0.1427523, 0.1294509, 
    0.1011614, 0.08765902, 0.08139436, 0.07169706, 0.05102765, 0.02733499, 
    -0.0007680357, -0.02961193, -0.06222074, -0.09684813, -0.1325748, 
    -0.1664787, -0.2125488, -0.2582929, -0.3018773, -0.3464777, -0.3807289, 
    -0.3969553, -0.3997538, -0.3974626, -0.402927, -0.4062014, -0.4046023, 
    -0.374008, -0.3658186, -0.3444706, -0.3004622, -0.2189498, -0.1212183, 
    -0.02714303, 0.05602945, 0.1224104, 0.1691554, 0.1974909, 0.1936504, 
    0.1768724, 0.1408072, 0.1002251, 0.06363723, 0.03675677, 0.009540883, 
    -0.0141961, -0.02647711, -0.01996068, -0.04894318, -0.1248063, 
    -0.1767879, -0.1769828, -0.1760513, -0.1717585, -0.1871467, -0.1736232, 
    -0.1811714, -0.1981892, -0.1938534, -0.1789772, -0.1712595, -0.1650746, 
    -0.1652959, -0.1524386, -0.1471755, -0.1532966, -0.1912641, -0.2642267, 
    -0.3657527, -0.4624313, -0.5827619, -0.6194216, -0.5752977, -0.4547083, 
    -0.3973645, -0.2745644, -0.190249, -0.1009791, -0.02039529, -0.159053, 
    -0.1851422, -0.2248071, -0.2415594, -0.2679482, -0.2642789,
  -0.2886809, -0.2766625, -0.2745605, -0.262129, -0.2559635, -0.2404911, 
    -0.2312542, -0.2137257, -0.202073, -0.1795374, -0.162235, -0.1386811, 
    -0.1235083, -0.1010077, -0.08529781, -0.06376503, -0.05096771, 
    -0.03426841, -0.02449601, -0.006322113, 0.00347887, 0.01425449, 
    0.01888739, 0.03537259, 0.05117082, 0.06746092, 0.06585696, 0.06500334, 
    0.06371535, 0.08692557, 0.1054735, 0.1286679, 0.1401202, 0.1460114, 
    0.1481913, 0.1484681, 0.1423701, 0.1153859, 0.07800721, 0.06187907, 
    0.06869207, 0.07511482, 0.08399272, 0.09802555, 0.1165684, 0.1300554, 
    0.1299168, 0.1134513, 0.09909937, 0.08860137, 0.08260584, 0.07096635, 
    0.05140817, 0.02000041, -0.0160144, -0.05161196, -0.08626965, -0.1261972, 
    -0.1617416, -0.2075209, -0.2641434, -0.3182741, -0.3793275, -0.4263052, 
    -0.4491984, -0.4550353, -0.4629098, -0.4791616, -0.4893886, -0.4985278, 
    -0.4978545, -0.4861819, -0.4577739, -0.4344099, -0.3950304, -0.333331, 
    -0.2393784, -0.1305461, -0.01862688, 0.07957941, 0.1564243, 0.186207, 
    0.1765653, 0.1484841, 0.1061567, 0.06331325, 0.03446109, 0.002190145, 
    -0.02831566, -0.04375045, -0.04448462, -0.07750203, -0.1570859, 
    -0.2029879, -0.2026134, -0.205969, -0.2012838, -0.2131536, -0.2147564, 
    -0.2174627, -0.207937, -0.2064714, -0.2082001, -0.2099641, -0.2068066, 
    -0.2105665, -0.2062973, -0.1954188, -0.181417, -0.1822273, -0.2077476, 
    -0.2871026, -0.3861459, -0.5004607, -0.6154474, -0.6077082, -0.5103356, 
    -0.4678077, -0.3137505, -0.265767, -0.0899442, -0.009940647, -0.1542852, 
    -0.191142, -0.2458302, -0.2577348, -0.278985, -0.2837887,
  -0.2941173, -0.2928752, -0.2874632, -0.2807429, -0.2737283, -0.2644065, 
    -0.2530779, -0.2378092, -0.2212387, -0.2045927, -0.1890163, -0.1694361, 
    -0.1502824, -0.1290293, -0.1118481, -0.0929721, -0.0783561, -0.06139418, 
    -0.04787375, -0.03281686, -0.02439564, -0.01260359, -0.0043009, 
    0.009243516, 0.01836705, 0.03090397, 0.04143776, 0.05619437, 0.06103215, 
    0.07035246, 0.07700152, 0.08304607, 0.08500513, 0.08576639, 0.078215, 
    0.07050467, 0.05468864, 0.04631987, 0.05441082, 0.06647189, 0.07560585, 
    0.08326852, 0.08845291, 0.09143973, 0.09553115, 0.1001844, 0.1043857, 
    0.1086038, 0.107152, 0.1008601, 0.09077152, 0.07851403, 0.06074986, 
    0.03357583, -0.001233459, -0.04358506, -0.08404113, -0.1184686, 
    -0.1506961, -0.1902869, -0.2498581, -0.3072217, -0.3756025, -0.4484921, 
    -0.4960913, -0.5143425, -0.5226943, -0.5423377, -0.5637279, -0.589375, 
    -0.6203667, -0.6413724, -0.6500661, -0.6301892, -0.5856156, -0.5334964, 
    -0.4685566, -0.3815867, -0.2691348, -0.1378258, 0.001354292, 0.1268917, 
    0.1903817, 0.1738309, 0.1318106, 0.09041724, 0.02860647, -0.01121531, 
    -0.03706193, -0.05818082, -0.06273738, -0.1028655, -0.1853438, 
    -0.2179022, -0.2117454, -0.2192813, -0.2188765, -0.2185682, -0.2224701, 
    -0.2154052, -0.2131165, -0.2124621, -0.2047029, -0.1983977, -0.1957654, 
    -0.2050858, -0.2226811, -0.2330435, -0.2231593, -0.2109414, -0.2015405, 
    -0.2182429, -0.2898432, -0.3925674, -0.5104688, -0.6237665, -0.6217533, 
    -0.5138288, -0.3955428, -0.2978752, -0.1469677, -0.09025151, -0.1426492, 
    -0.2074272, -0.2403159, -0.2698374, -0.2840472, -0.291196,
  -0.2990917, -0.2957527, -0.2895918, -0.2863516, -0.2773764, -0.2712967, 
    -0.2604336, -0.2527699, -0.2397067, -0.2258432, -0.2054088, -0.189259, 
    -0.1717152, -0.1570011, -0.1387355, -0.1242347, -0.110069, -0.1003471, 
    -0.09186065, -0.08654466, -0.08084865, -0.07667179, -0.06922502, 
    -0.06269403, -0.05570697, -0.04838748, -0.04089961, -0.03158901, 
    -0.01732237, -0.008106582, -0.001915876, 0.001336105, -0.006851289, 
    0.00150945, -0.00937219, -0.006942008, 0.002891995, 0.01245984, 
    0.01890488, 0.0277436, 0.03479904, 0.04290625, 0.0507648, 0.06131067, 
    0.07115662, 0.08179466, 0.09121078, 0.1001241, 0.1033523, 0.1023532, 
    0.09464423, 0.0835327, 0.06804498, 0.05361947, 0.02924655, -0.003360927, 
    -0.03905112, -0.07479538, -0.1056806, -0.1421991, -0.2058414, -0.2771139, 
    -0.3447598, -0.4314076, -0.5082512, -0.5464991, -0.564408, -0.5876874, 
    -0.618138, -0.6739718, -0.7319921, -0.7580942, -0.7742577, -0.7847545, 
    -0.7880238, -0.7680418, -0.723592, -0.6536511, -0.5605689, -0.4379442, 
    -0.2891915, -0.1180191, 0.05750789, 0.1758018, 0.1814101, 0.1214745, 
    0.05518555, 0.01690356, -0.02458149, -0.05663306, -0.06411539, 
    -0.09350162, -0.1713027, -0.2115415, -0.2131071, -0.2293681, -0.2291022, 
    -0.216639, -0.2248999, -0.2230881, -0.2150747, -0.1916757, -0.1854716, 
    -0.1967061, -0.2020203, -0.2041058, -0.2085192, -0.2325768, -0.2507363, 
    -0.2464491, -0.2378114, -0.2188333, -0.2251052, -0.2830968, -0.383268, 
    -0.4863066, -0.6073917, -0.6230357, -0.5531008, -0.3955292, -0.2510683, 
    -0.08639482, -0.02392322, -0.1832237, -0.2313824, -0.2742775, -0.2908578, 
    -0.3021634,
  -0.2940225, -0.2935326, -0.2904034, -0.2858093, -0.2837541, -0.2799169, 
    -0.2751323, -0.2648498, -0.2533696, -0.2439995, -0.2363943, -0.2233255, 
    -0.2057095, -0.18682, -0.1724711, -0.1598998, -0.1488403, -0.136703, 
    -0.125914, -0.1144525, -0.1043935, -0.09066014, -0.07888963, -0.06846163, 
    -0.06263336, -0.05776396, -0.05382333, -0.04887837, -0.04954316, 
    -0.04600389, -0.04599247, -0.03264384, -0.03777013, -0.03035903, 
    -0.02405316, -0.02274073, -0.02659746, -0.0281968, -0.02615819, 
    -0.02144937, -0.0170335, -0.009182241, -0.000440985, 0.00909498, 
    0.01790096, 0.02768422, 0.03576422, 0.04338805, 0.04852478, 0.05298467, 
    0.05452224, 0.05524897, 0.05155677, 0.04436037, 0.03072737, 0.01823507, 
    -0.007775813, -0.03406523, -0.05997093, -0.09752084, -0.1465912, 
    -0.2241488, -0.2903801, -0.3701888, -0.4773066, -0.5576888, -0.5870876, 
    -0.6094507, -0.64433, -0.7070472, -0.766269, -0.8083404, -0.8610203, 
    -0.9131097, -0.9403224, -0.9498314, -0.9447654, -0.9173822, -0.8615671, 
    -0.7697461, -0.634125, -0.4543102, -0.2461946, -0.02360993, 0.1565593, 
    0.2028307, 0.1401615, 0.06577259, 0.01044594, -0.02595652, -0.04644512, 
    -0.07308091, -0.1527495, -0.2017839, -0.2047183, -0.2113769, -0.2073167, 
    -0.1988588, -0.1984359, -0.1926203, -0.1855349, -0.1750023, -0.1886512, 
    -0.1756627, -0.1593512, -0.1904569, -0.1975576, -0.2095755, -0.2341606, 
    -0.2430899, -0.254153, -0.2424267, -0.2231171, -0.2192059, -0.2728879, 
    -0.3679072, -0.459182, -0.570828, -0.6421064, -0.5644453, -0.3826252, 
    -0.2450135, -0.09929521, -0.1417457, -0.2174235, -0.2363813, -0.2715353, 
    -0.2842214,
  -0.2655071, -0.2704367, -0.2714588, -0.2769065, -0.2750499, -0.2738368, 
    -0.2667791, -0.2635034, -0.2563803, -0.2481363, -0.2353515, -0.2283728, 
    -0.216388, -0.2021995, -0.1808186, -0.1625687, -0.1406276, -0.122566, 
    -0.1015512, -0.08315957, -0.06547562, -0.05649755, -0.05132917, 
    -0.0548743, -0.0562988, -0.05423066, -0.04715238, -0.04387063, 
    -0.03292152, -0.03077292, -0.02945526, -0.03910509, -0.04359052, 
    -0.05266091, -0.06908263, -0.07841118, -0.08138103, -0.0841312, 
    -0.08913981, -0.09436853, -0.09678237, -0.09844398, -0.09704585, 
    -0.09213046, -0.08265521, -0.07111634, -0.05759256, -0.04379765, 
    -0.02969238, -0.01680161, -0.004697185, 0.00560995, 0.01504634, 
    0.02403508, 0.03100265, 0.03231169, 0.02784641, 0.02007391, -0.008302465, 
    -0.03870954, -0.06784467, -0.1398488, -0.2169265, -0.2859908, -0.3810113, 
    -0.5028574, -0.5766793, -0.605888, -0.6330801, -0.6970913, -0.7594919, 
    -0.8117479, -0.8877179, -0.9644158, -1.006953, -1.036397, -1.051981, 
    -1.050339, -1.0407, -1.011558, -0.9468483, -0.8228271, -0.6241891, 
    -0.3708567, -0.09462267, 0.1455521, 0.2303135, 0.1496648, 0.0682248, 
    0.0208735, -0.01881914, -0.03128757, -0.09151566, -0.1647792, -0.1740745, 
    -0.1737441, -0.1758288, -0.1750447, -0.1643192, -0.1626408, -0.1674916, 
    -0.1566213, -0.1460852, -0.1411853, -0.1580825, -0.1744031, -0.1575467, 
    -0.1844635, -0.2154361, -0.2144788, -0.2430075, -0.2502979, -0.2292901, 
    -0.216671, -0.2044604, -0.2546919, -0.3464165, -0.4255802, -0.5151513, 
    -0.6000246, -0.5697781, -0.3646834, -0.2033442, -0.05479792, -0.1305642, 
    -0.2297633, -0.2446206, -0.2654867,
  -0.2404888, -0.2539006, -0.2485815, -0.2564065, -0.2554854, -0.2654096, 
    -0.2638999, -0.2656903, -0.2522278, -0.2467684, -0.2333381, -0.2248125, 
    -0.2069689, -0.1923512, -0.1680127, -0.1449619, -0.1144513, -0.08638239, 
    -0.05821758, -0.04717895, -0.04099668, -0.04391786, -0.039846, 
    -0.03983258, -0.02944854, -0.02083012, -0.01150401, -0.01406877, 
    -0.02360798, -0.03455185, -0.04883911, -0.0474563, -0.06111858, 
    -0.06096325, -0.06708637, -0.07570061, -0.09764439, -0.1188322, 
    -0.1397999, -0.1551733, -0.1721154, -0.1845848, -0.1963076, -0.2029517, 
    -0.2079684, -0.2067677, -0.2025327, -0.1927881, -0.181374, -0.1662077, 
    -0.1498044, -0.1296832, -0.1082634, -0.08492245, -0.06080537, 
    -0.03388335, -0.009620227, 0.006905641, 0.01391249, 0.01221695, 
    -0.01075827, -0.06067833, -0.1242977, -0.1936796, -0.2713715, -0.3872586, 
    -0.5081834, -0.5757713, -0.6058494, -0.6520103, -0.7121686, -0.7589825, 
    -0.8465171, -0.9303471, -0.981902, -1.036091, -1.089364, -1.112064, 
    -1.123574, -1.114323, -1.092112, -1.046897, -0.9511738, -0.7580493, 
    -0.4668566, -0.1313286, 0.165409, 0.2769703, 0.180327, 0.09665154, 
    0.04937905, 0.0226294, -0.005166373, -0.08221574, -0.1171695, -0.1175331, 
    -0.1275021, -0.1228493, -0.1133044, -0.1077197, -0.1070327, -0.1001809, 
    -0.1102207, -0.1141537, -0.1133277, -0.105477, -0.1322646, -0.1587526, 
    -0.1666455, -0.1684936, -0.2156418, -0.2236689, -0.2078416, -0.1965157, 
    -0.1873482, -0.173206, -0.2370271, -0.3173122, -0.4087315, -0.4610612, 
    -0.5856738, -0.5520955, -0.3229516, -0.037322, 0.07779481, -0.1226397, 
    -0.1869303, -0.2321594,
  -0.172401, -0.1838436, -0.1981402, -0.2094893, -0.2230787, -0.2352126, 
    -0.2429131, -0.2472768, -0.2499005, -0.2448469, -0.2288467, -0.2103249, 
    -0.1886977, -0.1705378, -0.1492769, -0.1175011, -0.08355182, -0.04982597, 
    -0.03037653, -0.01222165, -0.007421523, -0.0004288163, -0.001919936, 
    0.008525338, 0.009071399, 0.02123504, 0.01742518, 0.02120309, 
    0.009116061, 0.01203417, 0.0003677718, -0.007441022, -0.02299543, 
    -0.04411491, -0.07717439, -0.1112115, -0.1434704, -0.1698205, -0.1949219, 
    -0.2157679, -0.2335019, -0.2467503, -0.2583642, -0.2672845, -0.275229, 
    -0.2795179, -0.2807781, -0.2769626, -0.2698812, -0.2586308, -0.2455201, 
    -0.2291456, -0.2104628, -0.1867266, -0.1609237, -0.1328549, -0.103335, 
    -0.07034305, -0.04132443, -0.0199513, -0.01361045, -0.02318669, 
    -0.05313416, -0.09703495, -0.1560472, -0.2397333, -0.358072, -0.4674558, 
    -0.5391755, -0.5901339, -0.6459078, -0.6837103, -0.7534112, -0.841007, 
    -0.9022008, -0.9815893, -1.067909, -1.126417, -1.166836, -1.182125, 
    -1.180935, -1.161352, -1.112378, -1.019803, -0.8303154, -0.5036055, 
    -0.1111539, 0.2250787, 0.3302084, 0.2161129, 0.1405529, 0.1061631, 
    0.07867901, 0.01830262, -0.04799124, -0.05635455, -0.06356612, 
    -0.06406637, -0.05610824, -0.05119994, -0.05019193, -0.04496722, 
    -0.05107265, -0.0426352, -0.05624485, -0.07998699, -0.09427421, 
    -0.09392381, -0.1173115, -0.1519636, -0.178863, -0.1707774, -0.1585635, 
    -0.1593419, -0.1390939, -0.1136334, -0.1420428, -0.2132722, -0.2961434, 
    -0.3760932, -0.4265272, -0.5248926, -0.5001824, -0.2833309, -0.0199342, 
    -0.05424192, -0.1082586, -0.1392311,
  -0.1053744, -0.1345807, -0.1443199, -0.1654836, -0.1764276, -0.2012621, 
    -0.2172169, -0.2357152, -0.2291057, -0.2304083, -0.2215981, -0.2137253, 
    -0.2041877, -0.1816728, -0.1572285, -0.1166373, -0.09600732, -0.05760773, 
    -0.03306869, 0.002649819, 0.01691891, 0.035106, 0.04513979, 0.05738069, 
    0.06001985, 0.06285904, 0.05713057, 0.05228655, 0.04114113, 0.0224385, 
    -0.001749329, -0.03217191, -0.06841879, -0.1015242, -0.1290663, 
    -0.1547935, -0.1841381, -0.2155648, -0.2474521, -0.2787552, -0.3109345, 
    -0.3422149, -0.3730057, -0.4007839, -0.4239509, -0.4393376, -0.4467457, 
    -0.4454397, -0.43738, -0.4228514, -0.4033356, -0.3782631, -0.3479345, 
    -0.3114584, -0.2688664, -0.2211033, -0.1729708, -0.1276649, -0.08544356, 
    -0.04616771, -0.01242394, 0.01111919, 0.01734814, 0.0007655434, 
    -0.04321847, -0.1102496, -0.1948045, -0.2898335, -0.3943647, -0.4843189, 
    -0.5452872, -0.5905044, -0.6443385, -0.7249846, -0.7937201, -0.8815604, 
    -1.006349, -1.105438, -1.169995, -1.196338, -1.211373, -1.224988, 
    -1.220436, -1.165421, -1.043525, -0.82766, -0.4551513, -0.008562027, 
    0.3391513, 0.4049023, 0.2809129, 0.2155137, 0.1785053, 0.1501736, 
    0.08722907, 0.0400855, 0.0346485, 0.03489957, 0.02563249, 0.02445402, 
    0.02438779, 0.02959876, 0.0168469, 0.008162506, -0.001255468, 
    0.001235757, -0.01350807, -0.04403577, -0.07291311, -0.09376412, 
    -0.09723644, -0.09608103, -0.0940917, -0.08704914, -0.0555016, 
    -0.04264896, -0.07001273, -0.1422802, -0.2175128, -0.2958691, -0.3652934, 
    -0.4078618, -0.4512069, -0.4196134, -0.1149615, 0.1120835, 0.04376103, 
    -0.07709876,
  0.05232102, -0.01034555, -0.03150588, -0.06931265, -0.08602633, -0.1204447, 
    -0.1370551, -0.1712203, -0.1995761, -0.2143668, -0.2147087, -0.2023237, 
    -0.1907493, -0.1583431, -0.1543599, -0.1165398, -0.1036135, -0.0699524, 
    -0.0475822, -0.03210741, -0.01144096, 0.01137027, 0.02490951, 0.03613978, 
    0.0376087, 0.03626515, 0.02684305, 0.01414618, -0.002487388, -0.01752694, 
    -0.04184685, -0.07230245, -0.1077081, -0.1466578, -0.1946029, -0.2460911, 
    -0.3004512, -0.3536789, -0.4062364, -0.4529988, -0.4936166, -0.5258719, 
    -0.5521936, -0.572309, -0.5876836, -0.5965694, -0.6003275, -0.598186, 
    -0.59251, -0.5826078, -0.5693618, -0.5513107, -0.5286046, -0.4975054, 
    -0.456443, -0.4023887, -0.3356275, -0.2575699, -0.1775253, -0.1035542, 
    -0.04272362, 0.004601244, 0.03834323, 0.05541238, 0.04708592, 
    0.009222426, -0.04476051, -0.1035501, -0.2051763, -0.3371147, -0.4309804, 
    -0.4912577, -0.5272143, -0.5904939, -0.6721438, -0.7512149, -0.8969777, 
    -1.021513, -1.108018, -1.158814, -1.195771, -1.246022, -1.313571, 
    -1.32403, -1.222382, -1.022187, -0.7426656, -0.3164012, 0.1623886, 
    0.4804965, 0.479793, 0.3622414, 0.3079662, 0.2705291, 0.238818, 
    0.1800548, 0.1387476, 0.1329827, 0.1275408, 0.1233758, 0.1142874, 
    0.1162262, 0.1110199, 0.1065898, 0.08843565, 0.05804523, 0.0327078, 
    0.01528859, 0.003907677, -0.006696489, -0.007222753, -0.002593702, 
    0.01854005, 0.04648211, 0.06389758, 0.03996898, -0.01650084, -0.08811599, 
    -0.1646548, -0.2405436, -0.2977, -0.3504862, -0.3626538, -0.3913855, 
    -0.3026872, 0.1330547, 0.2822234, 0.07174995,
  0.1570651, 0.09393445, 0.02832346, -0.01820127, -0.06595713, -0.1106328, 
    -0.1447476, -0.1851186, -0.2168378, -0.2373874, -0.250727, -0.2560017, 
    -0.2542968, -0.1990208, -0.2008175, -0.1511158, -0.1223139, -0.1098441, 
    -0.07878084, -0.0383376, -0.02621364, -0.01641801, -0.01098782, 
    0.004647274, 0.01028765, 0.004844245, -0.0140273, -0.03246154, 
    -0.05656633, -0.08534086, -0.1251641, -0.1732391, -0.2338018, -0.2943821, 
    -0.3539964, -0.4077496, -0.4567481, -0.496384, -0.5319874, -0.5618564, 
    -0.589836, -0.6105942, -0.6278645, -0.6409643, -0.6526204, -0.6578055, 
    -0.659216, -0.6539812, -0.6463819, -0.6342149, -0.6197767, -0.5999717, 
    -0.577486, -0.5508571, -0.522325, -0.4873723, -0.4466213, -0.3935165, 
    -0.3230754, -0.2317027, -0.1308538, -0.0356074, 0.03667561, 0.08330254, 
    0.1037235, 0.1024442, 0.08084457, 0.03739186, -0.04622018, -0.1592464, 
    -0.2736201, -0.3559785, -0.3919135, -0.4572613, -0.5365431, -0.6060809, 
    -0.7617958, -0.9020321, -1.005864, -1.08117, -1.137247, -1.248513, 
    -1.409146, -1.468887, -1.399261, -1.206883, -0.9193351, -0.5646852, 
    -0.09584133, 0.3792572, 0.6272414, 0.5793186, 0.468998, 0.4224925, 
    0.3917059, 0.3580113, 0.3025337, 0.2663319, 0.2405433, 0.2385148, 
    0.2277258, 0.2229319, 0.2030852, 0.1793214, 0.1583348, 0.1471199, 
    0.1425638, 0.1294521, 0.1236839, 0.1277377, 0.1481485, 0.1732924, 
    0.197401, 0.1900235, 0.1511189, 0.08583715, 0.01238306, -0.07084823, 
    -0.1559057, -0.2345453, -0.301793, -0.3303006, -0.3365892, -0.2823174, 
    -0.2720743, -0.08118777, 0.33237, 0.2553886,
  0.3101113, 0.2370221, 0.132663, 0.05807521, -0.01200505, -0.08216919, 
    -0.1287074, -0.1567841, -0.1864984, -0.2137622, -0.2386346, -0.2689251, 
    -0.2662022, -0.2518673, -0.26686, -0.2410657, -0.2126785, -0.1957029, 
    -0.1868829, -0.1481624, -0.108335, -0.08834112, -0.09766835, -0.1047614, 
    -0.09648266, -0.09142805, -0.1082028, -0.1406291, -0.1884634, -0.2363495, 
    -0.2766241, -0.3126576, -0.3520627, -0.396847, -0.4464586, -0.4908616, 
    -0.5284756, -0.5649014, -0.6034399, -0.6389717, -0.6698231, -0.6945325, 
    -0.7138768, -0.7283424, -0.737492, -0.7404167, -0.7388688, -0.7332416, 
    -0.7240765, -0.7109014, -0.6929262, -0.6700613, -0.6419285, -0.6062156, 
    -0.5627786, -0.5127664, -0.4586621, -0.4041063, -0.3527489, -0.3002766, 
    -0.2347124, -0.1469663, -0.04351875, 0.05408528, 0.1264676, 0.1650051, 
    0.1713277, 0.1474821, 0.09037255, -0.01207372, -0.1291814, -0.2051896, 
    -0.2452654, -0.3169144, -0.3840943, -0.4592711, -0.6057307, -0.761731, 
    -0.8876423, -0.9781909, -1.047404, -1.239443, -1.457222, -1.500435, 
    -1.432507, -1.302926, -1.062725, -0.7237473, -0.3195994, 0.1690271, 
    0.5955429, 0.7796126, 0.7041393, 0.5984988, 0.5512003, 0.5221068, 
    0.4891881, 0.4487852, 0.406913, 0.3752303, 0.3514372, 0.3334455, 
    0.3237511, 0.3118008, 0.3088153, 0.2927569, 0.2862533, 0.2884843, 
    0.3124452, 0.3337909, 0.3525949, 0.3393216, 0.3023584, 0.2365369, 
    0.1614064, 0.06899385, -0.03087532, -0.1396236, -0.2347938, -0.3117077, 
    -0.3410023, -0.3469321, -0.3159842, -0.2833856, -0.1911539, -0.1059131, 
    0.2721876, 0.4873389,
  0.5449644, 0.3634583, 0.2470843, 0.1646805, 0.1076066, 0.07691174, 
    0.04273494, -0.008239873, -0.0426339, -0.07266725, -0.1088419, 
    -0.1421756, -0.1409632, -0.1859619, -0.1865419, -0.2001953, -0.1743914, 
    -0.1989837, -0.2052927, -0.1907427, -0.1606782, -0.1515437, -0.1535139, 
    -0.1669684, -0.1746093, -0.1822106, -0.1911055, -0.2225872, -0.2591141, 
    -0.2920359, -0.3212094, -0.364116, -0.4142643, -0.4693547, -0.5199004, 
    -0.5682432, -0.6124761, -0.6561954, -0.6903495, -0.718798, -0.7415812, 
    -0.7624482, -0.7787617, -0.7938684, -0.802761, -0.8073973, -0.8052931, 
    -0.7996947, -0.7885941, -0.7745082, -0.7543868, -0.7309008, -0.7010667, 
    -0.6674377, -0.6260188, -0.5768703, -0.5160165, -0.4453844, -0.3629598, 
    -0.2807611, -0.208368, -0.1507602, -0.09191979, -0.02124676, 0.05973164, 
    0.1304201, 0.1755904, 0.1802492, 0.1427377, 0.07474093, 0.008604519, 
    -0.04206073, -0.09360053, -0.1665897, -0.2338585, -0.3080676, -0.4503209, 
    -0.6239487, -0.7575228, -0.8468521, -0.9394693, -1.212232, -1.421476, 
    -1.399027, -1.314452, -1.217686, -1.090418, -0.8240066, -0.466944, 
    -0.04260536, 0.4300708, 0.7906148, 0.9287917, 0.863344, 0.7609121, 
    0.699973, 0.6713198, 0.6409541, 0.6157535, 0.5887527, 0.5656668, 
    0.5418558, 0.5179393, 0.4980839, 0.4880553, 0.4997101, 0.5190477, 
    0.5415744, 0.5403578, 0.5123156, 0.4512221, 0.3761806, 0.2840091, 
    0.1788347, 0.05335907, -0.07920377, -0.2087142, -0.319122, -0.4015259, 
    -0.4459177, -0.4566883, -0.4198663, -0.3345119, -0.2176081, -0.1078791, 
    -0.04339887, 0.2106755, 0.6430761,
  0.8101773, 0.5454631, 0.4130432, 0.316106, 0.2566937, 0.2434563, 0.2045604, 
    0.1708225, 0.1484069, 0.1273937, 0.108911, 0.06948498, 0.04451601, 
    -0.008529332, -0.04294071, -0.08687069, -0.1161336, -0.146696, 
    -0.1399538, -0.1536545, -0.1596154, -0.168047, -0.1687882, -0.1778384, 
    -0.185259, -0.1954849, -0.2187108, -0.257822, -0.2951701, -0.3377554, 
    -0.3902653, -0.4455236, -0.4932995, -0.5432612, -0.5918363, -0.6373541, 
    -0.6789432, -0.7214725, -0.7618409, -0.8004404, -0.8318655, -0.8580023, 
    -0.8768952, -0.8902246, -0.8954419, -0.8957313, -0.8897712, -0.8804685, 
    -0.866052, -0.848514, -0.8260642, -0.8007268, -0.7696919, -0.7318912, 
    -0.6844144, -0.6287641, -0.5639039, -0.4920309, -0.4128807, -0.3239611, 
    -0.2234723, -0.1226731, -0.03867438, 0.02237815, 0.07143086, 0.1169969, 
    0.1563928, 0.1806067, 0.184255, 0.1660993, 0.1337034, 0.09338694, 
    0.03888529, -0.02533431, -0.07840631, -0.1488249, -0.3101567, -0.481367, 
    -0.6141326, -0.7031679, -0.828956, -1.158372, -1.314198, -1.254869, 
    -1.182857, -1.065614, -0.9621629, -0.8346035, -0.5547069, -0.2003639, 
    0.2117615, 0.6423013, 0.9485461, 1.074243, 1.042278, 0.9608796, 
    0.8924923, 0.8446985, 0.8075458, 0.7799279, 0.7527761, 0.7404579, 
    0.7339633, 0.7502735, 0.7654779, 0.7747326, 0.7528985, 0.7027519, 
    0.6183986, 0.5214716, 0.407903, 0.2770997, 0.1217722, -0.03880421, 
    -0.1932876, -0.3240078, -0.4336084, -0.5116427, -0.5622383, -0.574958, 
    -0.5411654, -0.4663478, -0.366636, -0.2449366, -0.0618923, 0.1026915, 
    0.2203769, 0.6841056,
  1.020641, 0.75958, 0.6008103, 0.4920465, 0.4349056, 0.4397265, 0.4463219, 
    0.4164915, 0.397673, 0.4018155, 0.3952848, 0.3364766, 0.2673606, 
    0.2137456, 0.1317235, 0.0862768, 0.007300792, -0.02404824, -0.07000525, 
    -0.1014054, -0.1217899, -0.1348927, -0.15697, -0.1859301, -0.2135695, 
    -0.2369525, -0.268215, -0.2988466, -0.3336436, -0.3759953, -0.4267792, 
    -0.4801764, -0.5418636, -0.6008936, -0.6564232, -0.7094702, -0.7641277, 
    -0.8108625, -0.8472465, -0.8707212, -0.8883271, -0.9000476, -0.9097387, 
    -0.9138889, -0.9147052, -0.9085115, -0.8987963, -0.8829741, -0.864782, 
    -0.8419653, -0.8188771, -0.7916365, -0.7627105, -0.7295028, -0.6939695, 
    -0.6494628, -0.5958497, -0.5263075, -0.4426333, -0.3475547, -0.2507651, 
    -0.1480869, -0.04185568, 0.06080471, 0.140257, 0.1968796, 0.2331315, 
    0.2573575, 0.2645299, 0.2624545, 0.2458674, 0.2188293, 0.1751905, 
    0.1345092, 0.0836812, -0.01719235, -0.1894593, -0.3333023, -0.4706441, 
    -0.5502383, -0.7218593, -1.082335, -1.164952, -1.101666, -1.065633, 
    -0.9878742, -0.8335669, -0.7027214, -0.5744262, -0.2997108, 0.03168474, 
    0.4071915, 0.774294, 1.047328, 1.19094, 1.22468, 1.194996, 1.151574, 
    1.111169, 1.082946, 1.065671, 1.056945, 1.044346, 1.015952, 0.9652973, 
    0.8918536, 0.7942283, 0.6775501, 0.5412646, 0.379133, 0.1918509, 
    0.002422649, -0.1703559, -0.3161901, -0.4410845, -0.5449423, -0.6283999, 
    -0.6845011, -0.710394, -0.6917254, -0.6420544, -0.5332571, -0.3666728, 
    -0.1665234, -0.0273408, 0.1823815, 0.3232223, 0.6685188,
  1.144355, 1.042702, 0.8357803, 0.7717199, 0.739027, 0.7581834, 0.7230902, 
    0.6806233, 0.6490418, 0.6448808, 0.5924478, 0.5228627, 0.4200652, 
    0.3860085, 0.3000822, 0.2470646, 0.1727915, 0.1050595, 0.01443213, 
    -0.03044619, -0.08074103, -0.1052046, -0.1311257, -0.1545416, -0.1906366, 
    -0.2299257, -0.2805915, -0.3234522, -0.3704001, -0.4183693, -0.4803911, 
    -0.5422408, -0.6036956, -0.6580085, -0.7126333, -0.7553852, -0.7930175, 
    -0.822555, -0.8562895, -0.8884435, -0.9230767, -0.9489682, -0.9695084, 
    -0.9759689, -0.9751042, -0.9625949, -0.9475541, -0.9246556, -0.8999177, 
    -0.8675619, -0.8359262, -0.8003711, -0.7646278, -0.7193713, -0.6695998, 
    -0.6117888, -0.5542483, -0.4946813, -0.4364333, -0.363391, -0.2732531, 
    -0.1671847, -0.06133981, 0.04654637, 0.1490698, 0.2402251, 0.3049679, 
    0.3490725, 0.3717462, 0.380798, 0.37059, 0.3526174, 0.3207657, 0.2799239, 
    0.2060473, 0.08907199, -0.06199236, -0.1920474, -0.3367547, -0.3972711, 
    -0.6382475, -0.9822164, -0.9886014, -0.954945, -0.9017421, -0.830513, 
    -0.7692322, -0.6131681, -0.4642662, -0.3339467, -0.1016784, 0.1925986, 
    0.5162244, 0.8165786, 1.049642, 1.198482, 1.278136, 1.303328, 1.299095, 
    1.273025, 1.235532, 1.181166, 1.113518, 1.028235, 0.9262234, 0.797271, 
    0.6434931, 0.4582517, 0.254438, 0.0520317, -0.1237327, -0.2779651, 
    -0.4158969, -0.5448761, -0.6539385, -0.7384573, -0.7917892, -0.8133405, 
    -0.7997032, -0.75459, -0.658202, -0.5332476, -0.3913066, -0.1755899, 
    0.07850882, 0.2685235, 0.448976, 0.6913238,
  1.189276, 1.314899, 1.057596, 1.052498, 1.06925, 1.014737, 0.9527469, 
    0.9124994, 0.856768, 0.7942554, 0.6984789, 0.5920067, 0.5107944, 
    0.471435, 0.4006544, 0.3410525, 0.2836013, 0.2052433, 0.1270574, 
    0.064736, -0.005547205, -0.06140745, -0.1094015, -0.1457082, -0.1855033, 
    -0.2352672, -0.292193, -0.3456728, -0.397875, -0.4508686, -0.5057895, 
    -0.5584475, -0.6130712, -0.6630639, -0.7136701, -0.7725999, -0.8417636, 
    -0.9078914, -0.9642049, -1.003176, -1.024798, -1.026492, -1.015645, 
    -0.9938514, -0.9679705, -0.9373474, -0.9065472, -0.8721147, -0.838299, 
    -0.8033242, -0.7722815, -0.7420928, -0.7156515, -0.6898826, -0.6611591, 
    -0.6188834, -0.5586127, -0.4792269, -0.391843, -0.3112689, -0.2410981, 
    -0.1655467, -0.0739066, 0.02882404, 0.1313756, 0.23077, 0.3201567, 
    0.3915231, 0.4369433, 0.4625472, 0.4689195, 0.4591396, 0.4293489, 
    0.3811998, 0.2973084, 0.1782007, 0.04550759, -0.08368964, -0.2011138, 
    -0.2543599, -0.5812143, -0.8501574, -0.8125266, -0.7992585, -0.7270397, 
    -0.6612874, -0.60482, -0.5622365, -0.4193513, -0.2604009, -0.1313428, 
    0.03444453, 0.2613558, 0.5155928, 0.7572045, 0.9447113, 1.07216, 
    1.141554, 1.167599, 1.154833, 1.11437, 1.044391, 0.9491031, 0.8209926, 
    0.66637, 0.4870817, 0.2984802, 0.1151403, -0.04637168, -0.1989297, 
    -0.3508863, -0.5013742, -0.6284129, -0.7217909, -0.773174, -0.7951926, 
    -0.7893055, -0.7743745, -0.7455537, -0.7046025, -0.6404331, -0.5058971, 
    -0.2971107, -0.1116318, 0.1291673, 0.3739087, 0.5639969, 0.7512036,
  1.182325, 1.50642, 1.346518, 1.263252, 1.322338, 1.285483, 1.232398, 
    1.120267, 0.981786, 0.860056, 0.7735049, 0.699029, 0.6513325, 0.5718952, 
    0.4632837, 0.3902267, 0.3356447, 0.2714171, 0.2172059, 0.1545556, 
    0.07750165, -0.004206553, -0.06936499, -0.1188982, -0.1684372, 
    -0.2263809, -0.2856857, -0.3394293, -0.3894422, -0.4416411, -0.4994979, 
    -0.5621724, -0.6318128, -0.7186854, -0.8153989, -0.8970901, -0.9398239, 
    -0.9425199, -0.9150145, -0.8718066, -0.8203499, -0.7683316, -0.7163638, 
    -0.6686984, -0.6251789, -0.5872234, -0.552986, -0.5225642, -0.4934482, 
    -0.4670231, -0.442877, -0.4245972, -0.4137969, -0.4093767, -0.4134009, 
    -0.4238334, -0.4335386, -0.4265226, -0.3887037, -0.3113611, -0.2129218, 
    -0.1188749, -0.04007632, 0.03787711, 0.123168, 0.2131449, 0.2993107, 
    0.3785839, 0.4445147, 0.4900366, 0.5114807, 0.5110883, 0.4876204, 
    0.4342259, 0.3503372, 0.2479936, 0.142215, 0.02028663, -0.05156504, 
    -0.1559346, -0.5443575, -0.6850188, -0.6452377, -0.6369568, -0.5932164, 
    -0.6016687, -0.5388913, -0.4584317, -0.3908866, -0.2826606, -0.1262568, 
    0.004936058, 0.1265617, 0.2630423, 0.4206862, 0.5742801, 0.7018886, 
    0.7842447, 0.821135, 0.8119902, 0.7641647, 0.680601, 0.5708305, 
    0.4422247, 0.3052932, 0.1649753, 0.02690898, -0.1197249, -0.2785624, 
    -0.4358237, -0.5615755, -0.6440494, -0.6817275, -0.6873289, -0.6699136, 
    -0.6426684, -0.6133534, -0.5810597, -0.5454239, -0.5105839, -0.4491693, 
    -0.3992031, -0.2487095, -0.01829772, 0.2100696, 0.4648862, 0.6878635, 
    0.8345501,
  1.144064, 1.53431, 1.647951, 1.542931, 1.534704, 1.511692, 1.408937, 
    1.226601, 1.036877, 0.8908454, 0.7942334, 0.7377355, 0.6932752, 
    0.6184404, 0.535209, 0.4540635, 0.3927751, 0.344502, 0.2960011, 
    0.2306771, 0.1502216, 0.0563273, -0.02123127, -0.07919546, -0.1327828, 
    -0.1981706, -0.2574938, -0.3174114, -0.3794893, -0.4541585, -0.5399667, 
    -0.6419687, -0.7460176, -0.8142262, -0.8183612, -0.7741349, -0.7016636, 
    -0.6237806, -0.5443166, -0.4780996, -0.4201822, -0.3752936, -0.335247, 
    -0.3065226, -0.2799822, -0.2577792, -0.2338724, -0.2123016, -0.1877469, 
    -0.1661531, -0.1429919, -0.1242577, -0.1072364, -0.1000429, -0.09844732, 
    -0.107049, -0.1254772, -0.1582982, -0.1926788, -0.2148678, -0.1952904, 
    -0.1253693, -0.02397889, 0.0718751, 0.1523161, 0.2239909, 0.2977105, 
    0.3660758, 0.4266668, 0.4735014, 0.5070431, 0.5145268, 0.4992695, 
    0.4553508, 0.3975432, 0.3139866, 0.2209584, 0.1173714, 0.09227002, 
    -0.1271053, -0.4851753, -0.503855, -0.4939132, -0.4805472, -0.4909029, 
    -0.4781919, -0.4445194, -0.4139744, -0.3312573, -0.2670601, -0.1917577, 
    -0.07858445, 0.04674701, 0.1526734, 0.2428693, 0.3204058, 0.3860903, 
    0.4317853, 0.4523588, 0.4442033, 0.4096482, 0.3505428, 0.2710066, 
    0.1715555, 0.0550049, -0.07834445, -0.2228131, -0.357688, -0.4570387, 
    -0.5161923, -0.5442585, -0.548757, -0.533682, -0.5063098, -0.4724514, 
    -0.435813, -0.3879982, -0.3472274, -0.3274345, -0.3329098, -0.2938095, 
    -0.1988757, -0.1043276, 0.0943473, 0.3140613, 0.540199, 0.7824517, 
    0.9324728,
  1.143755, 1.402145, 1.690734, 1.769906, 1.740628, 1.672063, 1.523281, 
    1.310816, 1.118928, 0.9782242, 0.8624638, 0.7619611, 0.6891671, 
    0.6544738, 0.5915456, 0.5245397, 0.4779502, 0.4204228, 0.3604498, 
    0.2993546, 0.2104273, 0.1148359, 0.03844005, -0.02941411, -0.103294, 
    -0.1840734, -0.2629672, -0.34829, -0.4491425, -0.5588123, -0.6581352, 
    -0.7118312, -0.6852433, -0.5971808, -0.5007116, -0.4172249, -0.3526284, 
    -0.3022743, -0.2666159, -0.2460713, -0.2346816, -0.233035, -0.2331731, 
    -0.2321284, -0.2257001, -0.2163043, -0.2005081, -0.1825932, -0.1582674, 
    -0.1313749, -0.09825272, -0.06421353, -0.02526125, 0.01367306, 
    0.05193283, 0.07768694, 0.09248997, 0.09077461, 0.07366679, 0.03915885, 
    -0.0001625568, -0.03176576, -0.01773161, 0.05021062, 0.1510934, 
    0.2437448, 0.3189065, 0.3800755, 0.4367962, 0.4798502, 0.5097109, 
    0.5216488, 0.5181369, 0.4906145, 0.4439228, 0.3739336, 0.2980006, 
    0.2425172, 0.188114, -0.1595632, -0.3750902, -0.3409089, -0.3467853, 
    -0.3537758, -0.3725607, -0.3696485, -0.3792938, -0.3492252, -0.3253496, 
    -0.2638197, -0.1984227, -0.1428441, -0.08252114, -0.00419235, 0.07283043, 
    0.1396151, 0.1860974, 0.2132295, 0.2161335, 0.196941, 0.1522044, 
    0.08684903, 0.001096327, -0.09525337, -0.1964768, -0.2851682, -0.3493184, 
    -0.389268, -0.4211209, -0.4402103, -0.4359289, -0.4086245, -0.3713026, 
    -0.3298792, -0.3002365, -0.2720169, -0.2185076, -0.1088607, -0.03118072, 
    -0.06336814, -0.1045231, -0.02794364, 0.0524448, 0.195393, 0.421324, 
    0.6237363, 0.8477758, 1.022116,
  1.174149, 1.28593, 1.476978, 1.649552, 1.700899, 1.638384, 1.497038, 
    1.337128, 1.22295, 1.111223, 0.9691868, 0.845512, 0.7753125, 0.7342544, 
    0.6834958, 0.6394941, 0.5655518, 0.4852444, 0.4201152, 0.3527016, 
    0.2544586, 0.1608419, 0.0662568, -0.02859373, -0.1254185, -0.2331127, 
    -0.3486559, -0.4695077, -0.5676793, -0.6093646, -0.5706296, -0.466904, 
    -0.3603055, -0.285576, -0.2371956, -0.2046507, -0.191963, -0.1866663, 
    -0.1912445, -0.195712, -0.1985013, -0.1891015, -0.175532, -0.1569337, 
    -0.1443081, -0.1286386, -0.1190009, -0.1055349, -0.09568331, -0.08145486, 
    -0.06871459, -0.04720322, -0.02124352, 0.01582298, 0.06171148, 0.1175482, 
    0.1663147, 0.1991757, 0.2099756, 0.2081642, 0.1955793, 0.1757314, 
    0.1439332, 0.1183945, 0.1363278, 0.2108664, 0.3096335, 0.3963939, 
    0.4573915, 0.5052749, 0.5390728, 0.5584005, 0.5539932, 0.5366968, 
    0.4936344, 0.4446974, 0.3785964, 0.3615328, 0.1715733, -0.1747997, 
    -0.2199183, -0.2069599, -0.2189272, -0.2408289, -0.2563221, -0.2819304, 
    -0.2833308, -0.2836876, -0.2723338, -0.2572377, -0.238365, -0.1902231, 
    -0.1424464, -0.1036606, -0.07183541, -0.04273532, -0.02256688, 
    -0.01413858, -0.02094168, -0.04218056, -0.07603003, -0.1196665, 
    -0.1677364, -0.2156655, -0.2565447, -0.2908479, -0.3215965, -0.3432557, 
    -0.3346204, -0.29539, -0.2440701, -0.1933123, -0.1408091, -0.09273911, 
    -0.06763773, -0.0662514, -0.04022101, 0.02410109, 0.1112088, 0.1133618, 
    0.06420761, 0.1470206, 0.2450381, 0.3378141, 0.5134244, 0.6956112, 
    0.8779533, 1.061222,
  1.178163, 1.260812, 1.335715, 1.415991, 1.473614, 1.47451, 1.435667, 
    1.37959, 1.311671, 1.192413, 1.084837, 1.006443, 0.9271758, 0.869617, 
    0.8173153, 0.731792, 0.6244036, 0.5454536, 0.4722788, 0.3859332, 
    0.2733185, 0.1547791, 0.04248001, -0.08285886, -0.2295115, -0.3710102, 
    -0.4845552, -0.5235404, -0.4797377, -0.3752414, -0.2601839, -0.1870798, 
    -0.1500905, -0.1306603, -0.1196345, -0.1229064, -0.1225831, -0.1193514, 
    -0.1096797, -0.08901481, -0.05918996, -0.03693631, -0.02024653, 
    -0.01192726, -0.004077367, 0.002189643, 0.01165824, 0.02292513, 
    0.03463369, 0.04490894, 0.05167091, 0.05481086, 0.05596452, 0.06516875, 
    0.08569583, 0.126379, 0.1834636, 0.2416736, 0.2747748, 0.2814269, 
    0.2698669, 0.2611239, 0.2638447, 0.2649438, 0.2450493, 0.2369972, 
    0.2800149, 0.3712874, 0.4650491, 0.5302983, 0.5675431, 0.5880005, 
    0.5926712, 0.5750155, 0.5447499, 0.5013039, 0.4740387, 0.4070861, 
    0.07780106, -0.1114514, -0.08318145, -0.08364379, -0.1160826, -0.1355358, 
    -0.1602633, -0.1868358, -0.196252, -0.2119376, -0.2241392, -0.2294275, 
    -0.2175664, -0.2154754, -0.2030378, -0.1819464, -0.1550896, -0.1370699, 
    -0.1250824, -0.123465, -0.1278468, -0.1408018, -0.1586812, -0.1815811, 
    -0.2067515, -0.2308771, -0.248047, -0.2461118, -0.2186756, -0.1747475, 
    -0.1322318, -0.1028666, -0.07278043, -0.03767312, 0.01636522, 0.07876354, 
    0.138879, 0.177859, 0.2134824, 0.2576311, 0.2951544, 0.2815251, 
    0.2486036, 0.3043353, 0.3954557, 0.4470963, 0.5755411, 0.7474803, 
    0.8987012, 1.046523,
  1.111239, 1.197859, 1.261228, 1.305207, 1.334924, 1.347625, 1.345515, 
    1.324728, 1.2882, 1.241142, 1.206115, 1.140995, 1.066298, 1.000286, 
    0.9052911, 0.79933, 0.6838809, 0.6021186, 0.5067559, 0.374981, 0.2317485, 
    0.09618604, -0.06854068, -0.2529495, -0.3862762, -0.4376757, -0.3988767, 
    -0.309357, -0.2093723, -0.1237767, -0.07957694, -0.06107825, -0.05210014, 
    -0.05183497, -0.05186044, -0.03910563, -0.02106064, 0.0002096286, 
    0.02953041, 0.05308317, 0.06326316, 0.06745652, 0.06764311, 0.06689987, 
    0.06653422, 0.06659979, 0.07095484, 0.08045502, 0.09821469, 0.116766, 
    0.13472, 0.145104, 0.1534971, 0.1536724, 0.1563112, 0.1677013, 0.209331, 
    0.2695186, 0.3282108, 0.3517615, 0.3429853, 0.315203, 0.3003556, 
    0.3054442, 0.3264689, 0.3261634, 0.3272309, 0.3683073, 0.4580415, 
    0.5452393, 0.6057172, 0.6268849, 0.6296669, 0.6149666, 0.5975593, 
    0.5621409, 0.5417908, 0.295083, 0.03082324, 0.002266273, 0.02226877, 
    0.01817253, -0.02607829, -0.04664361, -0.07623813, -0.0977146, 
    -0.1218545, -0.1383065, -0.1593966, -0.1720523, -0.1855018, -0.1759422, 
    -0.1684185, -0.1656613, -0.1651126, -0.1596266, -0.1556744, -0.156012, 
    -0.1587978, -0.1590682, -0.1563156, -0.1552913, -0.145101, -0.124487, 
    -0.0936167, -0.05703961, -0.03410939, -0.009036534, 0.0324484, 
    0.09700195, 0.1524137, 0.2084367, 0.2404472, 0.2760526, 0.30716, 
    0.3405692, 0.3686951, 0.3917067, 0.4281373, 0.4269623, 0.3934181, 
    0.4318437, 0.5443849, 0.6022785, 0.6349139, 0.7371903, 0.881699, 1.003214,
  1.017553, 1.103922, 1.168746, 1.209521, 1.231153, 1.238684, 1.242505, 
    1.240974, 1.236951, 1.218684, 1.188556, 1.139302, 1.093056, 1.035431, 
    0.931748, 0.8218119, 0.7153151, 0.6305221, 0.4784464, 0.2973937, 
    0.133003, -0.07075366, -0.2672052, -0.35593, -0.3409108, -0.2576681, 
    -0.1734034, -0.1139214, -0.05348, -0.01293221, 0.002828006, 0.006552991, 
    0.008717049, 0.02199647, 0.0399102, 0.05713938, 0.08138072, 0.1174586, 
    0.1385165, 0.151869, 0.1645428, 0.1685578, 0.1640219, 0.1602589, 
    0.1530595, 0.1450897, 0.1340428, 0.1367806, 0.1478887, 0.1699302, 
    0.1868545, 0.2018233, 0.2094538, 0.2213957, 0.2290979, 0.2472157, 
    0.2807021, 0.3344683, 0.3643856, 0.3555765, 0.334296, 0.342986, 
    0.3543952, 0.350181, 0.351069, 0.3678585, 0.3788115, 0.4113798, 
    0.4861558, 0.5726532, 0.6342279, 0.6681607, 0.6715429, 0.6590856, 
    0.6299078, 0.6178862, 0.4461397, 0.1576191, 0.07973078, 0.09682645, 
    0.1036688, 0.07959118, 0.06117788, 0.02091716, -0.0007314608, 
    -0.03020634, -0.05092222, -0.07228988, -0.09666249, -0.1171888, 
    -0.1186811, -0.1289007, -0.13323, -0.1221905, -0.1119465, -0.1043711, 
    -0.09158385, -0.0743487, -0.06184604, -0.0535512, -0.04226509, 
    -0.02301099, -0.001369301, 0.01387141, 0.02335148, 0.04351082, 0.10362, 
    0.1809781, 0.2523248, 0.2792236, 0.2750971, 0.3041756, 0.3361134, 
    0.379421, 0.4296235, 0.4786682, 0.5194606, 0.5543891, 0.5795884, 
    0.6079098, 0.6021891, 0.5609265, 0.5735688, 0.6471161, 0.7042942, 
    0.7387122, 0.8119953, 0.9114046,
  0.8507268, 0.9181553, 0.9885946, 1.057192, 1.109517, 1.137354, 1.154877, 
    1.156471, 1.150944, 1.138028, 1.120958, 1.081257, 1.043613, 0.9810388, 
    0.8797482, 0.8012827, 0.7348664, 0.5984103, 0.3724887, 0.1628678, 
    -0.07022095, -0.2578348, -0.297511, -0.243973, -0.1302515, -0.05124795, 
    -0.0206891, 0.02147152, 0.04808692, 0.05299788, 0.05581656, 0.06987767, 
    0.08968943, 0.1010539, 0.1075405, 0.1313191, 0.1748095, 0.1996974, 
    0.2140915, 0.2390039, 0.2447285, 0.2286335, 0.2111268, 0.2024689, 
    0.1993227, 0.1870738, 0.1769128, 0.1838182, 0.2045534, 0.2243302, 
    0.2407054, 0.2553157, 0.261252, 0.2609294, 0.2795483, 0.3333474, 
    0.3871723, 0.4093376, 0.4050609, 0.3948976, 0.3699422, 0.3667673, 
    0.3872675, 0.3874479, 0.3808838, 0.4030471, 0.4278329, 0.4699284, 
    0.5404012, 0.6192091, 0.668245, 0.6881149, 0.6866915, 0.6800546, 
    0.6668042, 0.5394945, 0.264775, 0.1506466, 0.128821, 0.1655774, 
    0.1748563, 0.1373558, 0.1155133, 0.0876067, 0.05055839, 0.03187323, 
    0.008926284, -0.02220236, -0.03393608, -0.06116102, -0.08586569, 
    -0.0709824, -0.04280868, -0.03311843, -0.02527144, -0.02083004, 
    -0.004749017, 0.008129844, 0.01592437, 0.01958473, 0.03357124, 
    0.04831904, 0.063913, 0.09142724, 0.1593828, 0.2395149, 0.2659433, 
    0.2178298, 0.163894, 0.1169822, 0.107488, 0.1215563, 0.1517478, 
    0.1875964, 0.2392836, 0.2946755, 0.3550722, 0.4056145, 0.4645711, 
    0.5201532, 0.5889676, 0.6514505, 0.6791078, 0.6886846, 0.7242241, 
    0.7582368, 0.7842818, 0.8011796,
  0.7900581, 0.8084292, 0.8238093, 0.8484813, 0.8889092, 0.9279262, 
    0.9708736, 1.001394, 1.01463, 1.008085, 0.9848435, 0.9543989, 0.924743, 
    0.8604701, 0.8092273, 0.7854221, 0.6959071, 0.4661518, 0.1988755, 
    -0.06454195, -0.2384323, -0.2221583, -0.1666116, -0.08938807, 
    0.006324265, 0.03929025, 0.06960882, 0.07665416, 0.07694427, 0.09521617, 
    0.1165667, 0.1311359, 0.1368359, 0.1442504, 0.1603764, 0.1977082, 
    0.2338888, 0.2485396, 0.2768878, 0.3008575, 0.2941, 0.2735331, 0.2506393, 
    0.2414064, 0.2348686, 0.2189973, 0.2132803, 0.2300911, 0.2476738, 
    0.2616123, 0.278072, 0.2817009, 0.284122, 0.3384856, 0.4053046, 
    0.4308593, 0.4157012, 0.3939644, 0.4066104, 0.4247609, 0.4151069, 
    0.4161955, 0.4230436, 0.4170319, 0.427714, 0.4561929, 0.4941428, 
    0.546682, 0.6082039, 0.6557703, 0.6838214, 0.7004904, 0.704607, 
    0.6861134, 0.5738268, 0.3318301, 0.2135027, 0.1975439, 0.1799923, 
    0.1831774, 0.1898111, 0.1848502, 0.1550327, 0.1337613, 0.1033913, 
    0.0640958, 0.05082692, 0.03580365, -0.002627008, -0.0165442, -0.03130506, 
    -0.03502968, -0.004773237, 0.03846195, 0.06464709, 0.08948192, 
    0.09832481, 0.09648812, 0.08987041, 0.09933083, 0.1122563, 0.137156, 
    0.185352, 0.24773, 0.2582684, 0.1957915, 0.09923913, 0.06516879, 
    0.07560574, 0.1048474, 0.1304785, 0.1529303, 0.1705939, 0.1952777, 
    0.2152265, 0.2355269, 0.2463253, 0.2682545, 0.2793376, 0.3018758, 
    0.3296355, 0.3614486, 0.434321, 0.5116303, 0.5848232, 0.641884, 
    0.7107612, 0.7590392,
  0.5152077, 0.6040794, 0.6778327, 0.7379924, 0.7745769, 0.7965783, 
    0.8155993, 0.839618, 0.8525574, 0.8652869, 0.8579808, 0.8442948, 
    0.8088231, 0.7797671, 0.7738459, 0.7461811, 0.5618078, 0.2621517, 
    -0.04362962, -0.2122925, -0.177566, -0.07923188, -0.04606106, 
    -0.0005453266, 0.04433578, 0.06854434, 0.08086046, 0.09387016, 0.1243037, 
    0.1422743, 0.1543844, 0.159168, 0.1686914, 0.1748127, 0.1895411, 
    0.2257032, 0.2647741, 0.2877181, 0.3155309, 0.3255606, 0.3221704, 
    0.3016667, 0.2722976, 0.2595892, 0.2559637, 0.24192, 0.2439929, 0.261141, 
    0.2745209, 0.2859111, 0.2911331, 0.3091021, 0.3661456, 0.4198115, 
    0.4434589, 0.4570256, 0.4685328, 0.4685029, 0.462338, 0.4562731, 
    0.4546819, 0.4576938, 0.456041, 0.4700655, 0.5010825, 0.5390086, 
    0.572458, 0.6103325, 0.6396022, 0.675271, 0.6958197, 0.7118614, 
    0.6771243, 0.5687677, 0.352871, 0.2413966, 0.2156516, 0.1945839, 
    0.2449268, 0.2251432, 0.2164285, 0.196746, 0.1795433, 0.1509579, 
    0.1349017, 0.108868, 0.07084184, 0.0536691, 0.05143587, 0.01162781, 
    -0.01231562, -0.006442413, 0.02699184, 0.05688405, 0.08437694, 
    0.09955468, 0.112872, 0.1175844, 0.1360785, 0.1591079, 0.1964403, 
    0.2352383, 0.2503255, 0.1874332, 0.1041417, 0.07027857, 0.1017201, 
    0.1399922, 0.1525986, 0.1520766, 0.1624601, 0.183136, 0.2155349, 
    0.2475908, 0.2774065, 0.3051288, 0.327371, 0.3346903, 0.3301563, 
    0.321417, 0.3017924, 0.2962103, 0.2675443, 0.2650073, 0.2791196, 
    0.3240353, 0.3729558, 0.43754,
  0.1914086, 0.2250055, 0.2855359, 0.3817019, 0.500865, 0.6128474, 0.6911485, 
    0.7341688, 0.7549649, 0.7583165, 0.7541096, 0.7415905, 0.7216096, 
    0.7288054, 0.7312318, 0.6218674, 0.3253646, -0.01467669, -0.2034977, 
    -0.1544494, -0.07926797, -0.009533968, 0.02873441, 0.06814834, 
    0.08265539, 0.0949039, 0.1118208, 0.1374807, 0.1499313, 0.1622012, 
    0.1697372, 0.1763384, 0.1790205, 0.1858283, 0.1973656, 0.2337039, 
    0.2762409, 0.3049356, 0.3217711, 0.331461, 0.3431066, 0.3292133, 
    0.290108, 0.2683869, 0.2664185, 0.2606817, 0.256675, 0.271499, 0.2812422, 
    0.2864056, 0.2967843, 0.3641621, 0.4382513, 0.4588728, 0.4700504, 
    0.4813631, 0.4933154, 0.4922259, 0.4916302, 0.489462, 0.4874808, 
    0.4893706, 0.506922, 0.5340262, 0.565731, 0.5862436, 0.6121719, 
    0.6371281, 0.6711473, 0.6946778, 0.6901038, 0.640739, 0.5316725, 
    0.3467425, 0.2306531, 0.2241403, 0.1971521, 0.2099207, 0.2281371, 
    0.2303422, 0.2274303, 0.2118948, 0.1940391, 0.16785, 0.1394446, 
    0.1165879, 0.102112, 0.06700006, 0.04522515, 0.047131, 0.02516819, 
    -0.008220926, -0.004851155, 0.03155912, 0.07815214, 0.1186084, 0.1492329, 
    0.1718107, 0.189231, 0.2019547, 0.1996696, 0.1538767, 0.08968951, 
    0.04685941, 0.07018679, 0.1072666, 0.123826, 0.11694, 0.1210883, 
    0.1311486, 0.1536569, 0.1771766, 0.2104881, 0.2359755, 0.268729, 
    0.2931263, 0.3143921, 0.2978375, 0.2775531, 0.2495696, 0.2291811, 
    0.2021774, 0.2091964, 0.1984931, 0.1833945, 0.1661421, 0.1623578, 
    0.1790841,
  0.09236242, 0.1098514, 0.1152555, 0.1245586, 0.1636004, 0.2780254, 
    0.4378129, 0.5697287, 0.6426785, 0.6784388, 0.6871518, 0.6802066, 
    0.6830403, 0.6881156, 0.6290543, 0.3734106, 0.001606049, -0.2033809, 
    -0.1432805, -0.08131574, -0.05261199, 0.01488826, 0.03948649, 0.06079439, 
    0.07064018, 0.1014853, 0.1201762, 0.1397278, 0.1547405, 0.1699694, 
    0.1704804, 0.1729963, 0.1760792, 0.1862531, 0.1903885, 0.2126769, 
    0.2512506, 0.2952962, 0.3180526, 0.333537, 0.351701, 0.3447487, 
    0.3046449, 0.2647062, 0.2541527, 0.2629782, 0.2552225, 0.2687604, 
    0.2771208, 0.2750407, 0.3217978, 0.4146742, 0.4483606, 0.4703414, 
    0.4878213, 0.5063152, 0.5138409, 0.5136243, 0.5112002, 0.5119212, 
    0.5172589, 0.5324304, 0.5481969, 0.5718602, 0.5849, 0.6132765, 0.6376657, 
    0.6647981, 0.6677291, 0.6464806, 0.5785547, 0.467192, 0.3235507, 
    0.2263556, 0.2570639, 0.1770907, 0.1970265, 0.2428443, 0.2406116, 
    0.2390616, 0.2210074, 0.2029894, 0.1815496, 0.1657393, 0.1466147, 
    0.1212614, 0.09306138, 0.08046449, 0.05903134, 0.03210431, 0.02915655, 
    0.02635427, 0.005195074, -0.0105637, -0.004007276, 0.01738565, 
    0.04264061, 0.06404021, 0.06597136, 0.05662684, 0.03401019, 0.02358674, 
    0.04317089, 0.08208108, 0.107323, 0.1162355, 0.1240657, 0.1289343, 
    0.1286186, 0.129473, 0.1391946, 0.1553524, 0.1761923, 0.2002763, 0.23046, 
    0.2672445, 0.2919075, 0.2875124, 0.2734215, 0.2565305, 0.2311247, 
    0.2025311, 0.190573, 0.1562817, 0.1268644, 0.09334129, 0.0878592, 
    0.0758439,
  0.03432147, 0.03722867, 0.08452092, 0.08802414, 0.07261627, 0.08541571, 
    0.2042792, 0.3789468, 0.5199835, 0.5842059, 0.6138576, 0.6267008, 
    0.6197091, 0.5860719, 0.3842402, -0.009437488, -0.2548849, -0.2037564, 
    -0.084077, -0.05563217, -0.01328799, 0.02911931, 0.03976034, 0.0628805, 
    0.08991417, 0.1128993, 0.1251916, 0.1424704, 0.15219, 0.1590709, 
    0.1594808, 0.1615097, 0.1604988, 0.1671926, 0.1743494, 0.1861102, 
    0.2078985, 0.2477535, 0.2874329, 0.3165449, 0.3384029, 0.3434653, 
    0.3188593, 0.2653344, 0.2205867, 0.2370512, 0.2453528, 0.2421239, 
    0.2447427, 0.2534562, 0.3275931, 0.4073576, 0.4370556, 0.4684998, 
    0.4798652, 0.493618, 0.4913924, 0.4995584, 0.512876, 0.5280619, 
    0.5362502, 0.5472797, 0.5634032, 0.5784633, 0.5996059, 0.629542, 
    0.6276159, 0.6226178, 0.5714393, 0.5082494, 0.3999766, 0.2963071, 
    0.1983491, 0.2185932, 0.1990633, 0.1464834, 0.2176293, 0.2273065, 
    0.2326326, 0.2278382, 0.2216247, 0.2048937, 0.1791303, 0.147806, 
    0.1237656, 0.1068497, 0.09204192, 0.06498362, 0.04834034, 0.03932458, 
    0.0200735, 0.007480744, 0.008717731, 0.004584074, -0.005154625, 
    -0.01254934, -0.01250315, -0.01184937, -0.007658664, 0.002993986, 
    0.02422312, 0.04851505, 0.06514052, 0.07423495, 0.08765274, 0.1007245, 
    0.1004283, 0.09442823, 0.09321402, 0.09652254, 0.1014362, 0.1078293, 
    0.117452, 0.1304476, 0.149317, 0.1804786, 0.2298094, 0.2615277, 
    0.2471168, 0.2365124, 0.2310547, 0.2126267, 0.2063003, 0.2054453, 
    0.1795354, 0.1364816, 0.09824634, 0.05517224,
  0.1101033, 0.09240182, 0.07127133, 0.05411284, 0.0491352, 0.03342883, 
    0.1188673, 0.2663758, 0.4224266, 0.5157281, 0.5624834, 0.5483675, 
    0.5348929, 0.3692448, -0.01424251, -0.3043782, -0.2388418, -0.1323307, 
    -0.1029386, -0.05451555, -0.01419253, 0.008953858, 0.03304618, 
    0.06484295, 0.08168179, 0.09629832, 0.1085984, 0.1227019, 0.1341731, 
    0.1404504, 0.1371301, 0.1347673, 0.1359717, 0.1405905, 0.1462934, 
    0.1541417, 0.1638736, 0.1845448, 0.2196723, 0.2607595, 0.296546, 
    0.314727, 0.3129774, 0.2724981, 0.1919771, 0.1763068, 0.2163432, 
    0.2278826, 0.226163, 0.2291837, 0.2974305, 0.3832925, 0.4127056, 
    0.4362019, 0.4533837, 0.4623716, 0.4687396, 0.4886791, 0.5035042, 
    0.5128605, 0.5179238, 0.5355034, 0.5537919, 0.5638182, 0.5823988, 
    0.5759688, 0.5457362, 0.4986804, 0.426616, 0.3442786, 0.2537023, 
    0.1648102, 0.1672767, 0.2046305, 0.1123248, 0.1463913, 0.2024499, 
    0.1984928, 0.1954976, 0.1852913, 0.1764397, 0.1636372, 0.1513123, 
    0.1352369, 0.1102842, 0.08160235, 0.05961763, 0.05193711, 0.03619798, 
    0.01570098, 0.008325059, 0.002994802, -0.007474221, -0.01249544, 
    -0.01326584, -0.01257358, -0.01163334, -0.006389551, -0.001406297, 
    0.005036287, 0.01201492, 0.02283654, 0.04145329, 0.06511159, 0.08132248, 
    0.08947632, 0.09533804, 0.09682053, 0.0886208, 0.07837111, 0.06985156, 
    0.06537884, 0.06414029, 0.06745297, 0.07341562, 0.08709268, 0.1137819, 
    0.1662642, 0.2140396, 0.2244252, 0.2228555, 0.2154734, 0.2008102, 
    0.1859285, 0.1812769, 0.1763423, 0.1531624, 0.1333573,
  0.05781904, 0.04224314, 0.02829993, 0.02837569, 0.01086294, 0.04536325, 
    0.1322088, 0.2608857, 0.3945675, 0.448904, 0.4628505, 0.4508957, 
    0.3172901, -0.04758248, -0.3148947, -0.3047414, -0.161486, -0.1270468, 
    -0.08632034, -0.044239, -0.02101439, 0.006859273, 0.03760229, 0.05604956, 
    0.07127585, 0.0833243, 0.09456442, 0.1039589, 0.1102104, 0.1095209, 
    0.1065092, 0.1048075, 0.1038215, 0.1038003, 0.1078458, 0.1155866, 
    0.1254192, 0.1324408, 0.1469692, 0.1808216, 0.2278731, 0.267122, 
    0.2870942, 0.2779356, 0.1954037, 0.118364, 0.1456151, 0.1906203, 
    0.203365, 0.2013437, 0.2286034, 0.3169172, 0.3776312, 0.3969488, 
    0.4143133, 0.420191, 0.4269671, 0.4446266, 0.4605279, 0.474842, 
    0.4840078, 0.5007799, 0.5158951, 0.5088803, 0.4993587, 0.4729885, 
    0.4321996, 0.3745618, 0.3062145, 0.2297837, 0.1602183, 0.1181449, 
    0.1744543, 0.1624769, 0.08992707, 0.1589305, 0.1734793, 0.1625121, 
    0.1718004, 0.1755846, 0.1663382, 0.1459189, 0.1160279, 0.09109342, 
    0.07309707, 0.0571801, 0.03494233, 0.01033872, -0.0006041601, 
    -0.001420077, -0.01485003, -0.02429371, -0.02746476, -0.02904178, 
    -0.03316443, -0.03335369, -0.03316645, -0.02925782, -0.02480116, 
    -0.01244117, 0.004246138, 0.02385202, 0.03507842, 0.04237334, 0.04995218, 
    0.05963606, 0.05951878, 0.05758151, 0.05396179, 0.0493384, 0.03570873, 
    0.01967873, 0.004215062, -0.002014697, -0.00509122, -0.007429004, 
    -0.007481113, 0.01715335, 0.06615859, 0.1273162, 0.1603651, 0.1745849, 
    0.1807303, 0.1817484, 0.1673124, 0.1556627, 0.1304558, 0.0928499,
  0.1291198, 0.08429128, 0.06017457, 0.05638866, 0.08282843, 0.1429691, 
    0.1996106, 0.300348, 0.3686164, 0.40072, 0.3757226, 0.2099334, 
    -0.1198241, -0.3207348, -0.2775343, -0.1947762, -0.1514026, -0.1148691, 
    -0.0638334, -0.03956301, -0.006300043, 0.02122727, 0.04280787, 
    0.05561386, 0.06703503, 0.07299466, 0.08088642, 0.08692402, 0.09569998, 
    0.0959602, 0.09165631, 0.08609165, 0.08758159, 0.08825816, 0.09010942, 
    0.09205429, 0.09893482, 0.1068984, 0.1165027, 0.1312989, 0.1684321, 
    0.2150347, 0.2505725, 0.2751252, 0.2381668, 0.1302615, 0.098748, 
    0.1509861, 0.1792915, 0.1791523, 0.176964, 0.2415001, 0.3414791, 
    0.3755085, 0.3897328, 0.4007292, 0.4090836, 0.4304206, 0.4456538, 
    0.4539147, 0.4603035, 0.4576178, 0.4567327, 0.4401892, 0.4146708, 
    0.3746467, 0.3235754, 0.2622037, 0.2030744, 0.1543252, 0.1133133, 
    0.1209923, 0.1798041, 0.1303606, 0.0953472, 0.1519373, 0.1544997, 
    0.1710326, 0.1780528, 0.1647354, 0.1499754, 0.1341934, 0.1162607, 
    0.09107956, 0.06086663, 0.03549295, 0.01848333, 0.007895472, -0.0112292, 
    -0.02840652, -0.0284562, -0.02656982, -0.03008161, -0.03247139, 
    -0.03189726, -0.03111254, -0.02905114, -0.02233661, -0.01326445, 
    -0.003854245, 0.003679007, 0.01113401, 0.02230963, 0.03694475, 0.0474082, 
    0.05287874, 0.05834334, 0.06086567, 0.05537935, 0.0456543, 0.03136763, 
    0.009183183, -0.01717582, -0.03702578, -0.04796204, -0.05384406, 
    -0.06238778, -0.06517386, -0.05469348, -0.01775597, 0.04679324, 
    0.1031656, 0.1279384, 0.1397352, 0.1517139, 0.1560078, 0.1583705, 
    0.1601985,
  0.2055164, 0.2096774, 0.20207, 0.2120676, 0.2435898, 0.2648657, 0.2940944, 
    0.3286796, 0.3164814, 0.2180487, -0.001380943, -0.2612516, -0.3676959, 
    -0.2696253, -0.1803689, -0.1473879, -0.1123001, -0.06620398, -0.03405029, 
    -0.002830642, 0.0254508, 0.04410968, 0.05697496, 0.06511427, 0.07237747, 
    0.07909623, 0.08756203, 0.09677494, 0.1015508, 0.09645543, 0.0909711, 
    0.08947718, 0.087437, 0.08657044, 0.0893369, 0.09158581, 0.09139143, 
    0.09222731, 0.09735914, 0.1057281, 0.1246892, 0.1632249, 0.2120301, 
    0.2575563, 0.2790511, 0.211574, 0.1050491, 0.1068968, 0.1568288, 
    0.1711487, 0.165531, 0.1845587, 0.2787061, 0.3609058, 0.379333, 
    0.3812653, 0.3837081, 0.3950965, 0.4074799, 0.4132788, 0.4176602, 
    0.4008119, 0.3811885, 0.347927, 0.3060494, 0.2603252, 0.2175551, 
    0.1769399, 0.1414579, 0.1098812, 0.1037791, 0.1467284, 0.1735525, 
    0.1032229, 0.101243, 0.1572042, 0.1688714, 0.1773727, 0.1601762, 
    0.1514502, 0.1408848, 0.124155, 0.1024826, 0.08450455, 0.06739095, 
    0.04560509, 0.02124327, -5.339272e-05, -0.008903482, -0.01394372, 
    -0.02781986, -0.03453166, -0.03154228, -0.0271591, -0.02422385, 
    -0.02045277, -0.01619825, -0.01021706, -0.003324158, 0.006232269, 
    0.01830305, 0.0306779, 0.03824554, 0.04078945, 0.04403786, 0.04805358, 
    0.04717633, 0.04447851, 0.04367185, 0.04227635, 0.03533973, 0.01841675, 
    -0.00986664, -0.04013923, -0.06091976, -0.07603237, -0.08994398, 
    -0.1031802, -0.1158729, -0.1176097, -0.1112511, -0.080739, -0.02531657, 
    0.02449193, 0.07059681, 0.1065943, 0.1381154, 0.1698469,
  0.04750147, 0.09909357, 0.1455319, 0.1731147, 0.1860112, 0.1790199, 
    0.1375131, 0.05075717, -0.08897798, -0.2576299, -0.3753313, -0.3651022, 
    -0.2670869, -0.1861992, -0.1517175, -0.1162135, -0.07629824, -0.04256986, 
    -0.01227157, 0.01608171, 0.03393813, 0.04550323, 0.05330538, 0.06178056, 
    0.06834272, 0.07609692, 0.08324713, 0.09018454, 0.09380766, 0.09193534, 
    0.08768762, 0.08466775, 0.08405823, 0.08460616, 0.08437208, 0.08299046, 
    0.08030703, 0.08081189, 0.08334592, 0.08510689, 0.08980452, 0.1093007, 
    0.1459447, 0.188822, 0.2344515, 0.2612574, 0.1842023, 0.08746602, 
    0.1044362, 0.1504545, 0.16225, 0.1673373, 0.1985588, 0.2785404, 
    0.3538902, 0.3751674, 0.3677391, 0.3623673, 0.3608983, 0.3533922, 
    0.3454682, 0.3190477, 0.2909951, 0.2556459, 0.224115, 0.1907008, 
    0.1567403, 0.1235768, 0.102791, 0.09414372, 0.1148551, 0.155563, 
    0.1716046, 0.1040111, 0.1033853, 0.1633855, 0.1611466, 0.156339, 
    0.1563857, 0.1585298, 0.1474986, 0.1326278, 0.1101056, 0.0842458, 
    0.05752712, 0.0381192, 0.02134638, 0.007704332, -0.01263617, -0.02773505, 
    -0.02855586, -0.02812835, -0.03170276, -0.03235382, -0.02988161, 
    -0.02560363, -0.0197669, -0.01107553, -0.003586896, 0.003394775, 
    0.009039849, 0.0146262, 0.02269941, 0.03487664, 0.04513115, 0.05161795, 
    0.05698785, 0.05848415, 0.05218197, 0.04296704, 0.03427465, 0.02299257, 
    0.002759382, -0.02928659, -0.06132463, -0.07961556, -0.09338847, 
    -0.1097424, -0.1258853, -0.1417432, -0.1538532, -0.1651704, -0.1788167, 
    -0.1823474, -0.1608119, -0.1203695, -0.06619675, -0.007475957,
  -0.2332115, -0.213312, -0.1991279, -0.1933929, -0.2023183, -0.2341923, 
    -0.284049, -0.3396934, -0.3760887, -0.3689469, -0.3120174, -0.2437929, 
    -0.1983827, -0.1602515, -0.1198024, -0.08041486, -0.04673836, 
    -0.01538276, 0.01175483, 0.02963176, 0.03895947, 0.0473756, 0.05643281, 
    0.06413125, 0.0720029, 0.07944046, 0.08680488, 0.09523938, 0.09978689, 
    0.09488892, 0.08933236, 0.08668184, 0.08315545, 0.08190113, 0.08235796, 
    0.08133517, 0.07738785, 0.07336891, 0.07105312, 0.07145761, 0.07236765, 
    0.07685879, 0.09001762, 0.1176838, 0.1529021, 0.2085564, 0.2421349, 
    0.1631827, 0.07515598, 0.09424806, 0.1333425, 0.1392166, 0.1421244, 
    0.1823322, 0.262831, 0.3259445, 0.3536628, 0.3489476, 0.3325272, 
    0.3160756, 0.3039436, 0.2823042, 0.2647061, 0.2343651, 0.1980411, 
    0.1514286, 0.1151932, 0.09180319, 0.0808748, 0.08386174, 0.1197971, 
    0.1522602, 0.162609, 0.09176019, 0.09760135, 0.1582872, 0.1498142, 
    0.1685187, 0.171426, 0.1628169, 0.1473504, 0.1299747, 0.1076959, 
    0.08877058, 0.06686857, 0.04261762, 0.01868794, 0.0008384436, 
    -0.00786647, -0.01452398, -0.02964171, -0.03597177, -0.03399016, 
    -0.02991827, -0.02736585, -0.022728, -0.01834852, -0.01249525, 
    -0.006728739, 0.003367752, 0.01547746, 0.02824212, 0.03728919, 
    0.04311086, 0.04741225, 0.0515185, 0.04998108, 0.04710385, 0.04454324, 
    0.04115075, 0.03267637, 0.02197734, 0.00821346, -0.01233356, -0.04513176, 
    -0.08006041, -0.1018083, -0.11435, -0.1321497, -0.1498417, -0.1699801, 
    -0.1818478, -0.1932606, -0.2084982, -0.2324442, -0.2547219, -0.2606117, 
    -0.2526736,
  -0.3069582, -0.3118211, -0.3156021, -0.3227136, -0.3281765, -0.3315449, 
    -0.3297813, -0.3177615, -0.2980615, -0.2716941, -0.2384211, -0.204601, 
    -0.1685098, -0.1301185, -0.09411243, -0.05848645, -0.02694898, 
    -0.0005851313, 0.01510452, 0.02541386, 0.03491904, 0.04581101, 
    0.05503454, 0.06384405, 0.07055376, 0.07749339, 0.08501648, 0.09280452, 
    0.09411829, 0.08823935, 0.08342751, 0.08084203, 0.08150807, 0.08270541, 
    0.08080719, 0.07596102, 0.07061008, 0.06846987, 0.06584679, 0.05945836, 
    0.05461705, 0.05437075, 0.05550112, 0.06395547, 0.08331193, 0.1149935, 
    0.1772386, 0.2200177, 0.1529387, 0.06507902, 0.06960954, 0.1084385, 
    0.1170481, 0.1208348, 0.1568076, 0.2129361, 0.2772941, 0.313874, 
    0.3270938, 0.3176665, 0.301354, 0.2782567, 0.2521229, 0.2125703, 
    0.1724502, 0.127481, 0.09272557, 0.06906745, 0.06697288, 0.07884607, 
    0.1181268, 0.1373213, 0.1558099, 0.09612748, 0.09680533, 0.1593961, 
    0.1656474, 0.1776376, 0.1590241, 0.1524033, 0.1405023, 0.1267375, 
    0.1054204, 0.08296844, 0.05931492, 0.04195434, 0.02300156, 0.006994508, 
    -0.013979, -0.02663958, -0.02723504, -0.02710417, -0.03155032, 
    -0.03240399, -0.03110506, -0.02708226, -0.02199499, -0.01302029, 
    -0.004985817, 0.003513485, 0.009422407, 0.01556696, 0.02308843, 
    0.03441844, 0.04396184, 0.05165658, 0.05796199, 0.06067161, 0.05487427, 
    0.04593268, 0.03520907, 0.02231558, 0.006756052, -0.01009139, 
    -0.03126275, -0.0589028, -0.09368709, -0.1201925, -0.134823, -0.1476176, 
    -0.1600869, -0.177817, -0.2044451, -0.2277364, -0.246444, -0.2596838, 
    -0.2788257, -0.2954655,
  -0.2996732, -0.304483, -0.3095209, -0.3115653, -0.3134682, -0.3104224, 
    -0.3019831, -0.2910228, -0.2733704, -0.2386674, -0.1995756, -0.1678568, 
    -0.1375551, -0.1025369, -0.06556229, -0.03332257, -0.009985849, 
    0.005529769, 0.01670544, 0.0285188, 0.03935754, 0.04921605, 0.05805465, 
    0.06561179, 0.07345713, 0.08124176, 0.08869611, 0.09495196, 0.09658416, 
    0.09200097, 0.08930923, 0.08743577, 0.08407542, 0.08235604, 0.08140779, 
    0.07808734, 0.07180469, 0.06574486, 0.06048929, 0.05376261, 0.04609716, 
    0.04168932, 0.04025517, 0.04104715, 0.04630091, 0.05712663, 0.07631445, 
    0.1339777, 0.1930542, 0.1564838, 0.06883138, 0.03978468, 0.06624166, 
    0.09343438, 0.09800944, 0.0981003, 0.1406782, 0.1825076, 0.2179318, 
    0.2403081, 0.2496736, 0.2413551, 0.2247371, 0.1949213, 0.1620351, 
    0.1213245, 0.08769731, 0.06500363, 0.06809172, 0.07923758, 0.1088887, 
    0.1199602, 0.1426919, 0.08241218, 0.08880255, 0.167167, 0.1590396, 
    0.1565906, 0.1554463, 0.1579863, 0.1453384, 0.1307271, 0.1075975, 
    0.08774057, 0.06360716, 0.04001626, 0.01789027, 0.002867274, 
    -0.006153286, -0.01443565, -0.03052703, -0.0359716, -0.03385738, 
    -0.02914709, -0.02662993, -0.02204656, -0.01837394, -0.01237474, 
    -0.006765157, 0.003379352, 0.01522831, 0.02885026, 0.03886204, 0.0464755, 
    0.05187061, 0.05663051, 0.0547848, 0.05167869, 0.04876596, 0.04593397, 
    0.03777625, 0.02626243, 0.01011266, -0.008444242, -0.03047091, 
    -0.0532308, -0.07782049, -0.1075425, -0.1397362, -0.1604977, -0.1773605, 
    -0.1865963, -0.1957349, -0.2104321, -0.2346965, -0.2602846, -0.2790432, 
    -0.2898267,
  -0.2851675, -0.2921293, -0.2984048, -0.2989536, -0.2940744, -0.2814318, 
    -0.2684074, -0.2510195, -0.2269556, -0.1968844, -0.1716902, -0.1422552, 
    -0.1089509, -0.07449171, -0.04787689, -0.02682344, -0.0121795, 
    0.001917273, 0.01486813, 0.02752027, 0.03786691, 0.04826146, 0.05773147, 
    0.06684145, 0.07312384, 0.0795442, 0.08608875, 0.09389231, 0.09502882, 
    0.08903335, 0.08388007, 0.08008623, 0.08014908, 0.08092927, 0.078168, 
    0.07270753, 0.0671653, 0.06471404, 0.0596494, 0.04833713, 0.03802212, 
    0.03166556, 0.02723391, 0.02474886, 0.02354573, 0.0268136, 0.02970184, 
    0.03657271, 0.07976443, 0.1489137, 0.1621782, 0.1028397, 0.0383267, 
    0.02051152, 0.03286376, 0.05454604, 0.0754655, 0.07727148, 0.1005078, 
    0.1208045, 0.1364006, 0.1418801, 0.1398285, 0.1260941, 0.1137964, 
    0.0965014, 0.07443598, 0.05061775, 0.05262342, 0.0642885, 0.09575596, 
    0.1043884, 0.1266131, 0.06525689, 0.08879861, 0.1625674, 0.1508426, 
    0.1695489, 0.1675763, 0.159345, 0.1438516, 0.1286464, 0.1061871, 
    0.08472997, 0.06197542, 0.04456314, 0.02346417, 0.005530253, -0.01502776, 
    -0.02515548, -0.0250223, -0.02554321, -0.03093749, -0.03207105, 
    -0.03094714, -0.02646601, -0.02097686, -0.01150151, -0.003304567, 
    0.005854689, 0.01244509, 0.01899523, 0.02579935, 0.03621909, 0.04495918, 
    0.05274832, 0.05972452, 0.0636802, 0.05863918, 0.05013482, 0.03990709, 
    0.02805298, 0.01268084, -0.005964167, -0.02840792, -0.05085723, 
    -0.07446115, -0.09527974, -0.1177925, -0.1459505, -0.1719895, -0.1979016, 
    -0.2245501, -0.2420345, -0.2504844, -0.2550817, -0.2650511, -0.2753447,
  -0.2703786, -0.2740381, -0.2787501, -0.2784916, -0.2716182, -0.2580551, 
    -0.2444759, -0.2283428, -0.2074077, -0.1794967, -0.1497014, -0.117076, 
    -0.08858047, -0.06265585, -0.04272447, -0.02428164, -0.009490401, 
    0.006238908, 0.01892478, 0.03136878, 0.04149833, 0.05234534, 0.06008431, 
    0.06669945, 0.07361765, 0.08253658, 0.09043863, 0.09649276, 0.09435804, 
    0.08865312, 0.08618896, 0.08558745, 0.08321338, 0.08277566, 0.0817085, 
    0.07842407, 0.07105491, 0.06461319, 0.05736595, 0.04812586, 0.03761187, 
    0.03020617, 0.02380542, 0.01928993, 0.01288378, 0.00734736, 0.003698468, 
    0.002868131, -0.002173007, 0.01299864, 0.06062345, 0.115462, 0.1242488, 
    0.08863406, 0.04152361, 0.0173844, 0.005011663, 0.0109514, 0.02719887, 
    0.03114127, 0.04869481, 0.06214749, 0.07880081, 0.08623952, 0.09656619, 
    0.09659515, 0.07783067, 0.05345051, 0.0462586, 0.05294612, 0.08061588, 
    0.08882794, 0.1036148, 0.04863217, 0.1053563, 0.1607606, 0.1571269, 
    0.1696463, 0.1554387, 0.1531783, 0.1409789, 0.1276315, 0.1060209, 
    0.08637792, 0.06186652, 0.03902668, 0.01913386, 0.005708277, 
    -0.004138812, -0.01473445, -0.03117607, -0.03537595, -0.03219338, 
    -0.02697599, -0.02434211, -0.02003579, -0.01667759, -0.01075236, 
    -0.005143177, 0.004949059, 0.01640161, 0.03009357, 0.04107261, 
    0.05042981, 0.0572801, 0.06308961, 0.06150361, 0.0580983, 0.05484023, 
    0.05194122, 0.04352781, 0.03181822, 0.01605788, -0.001911841, 
    -0.02512437, -0.05088694, -0.0753824, -0.09758398, -0.1191483, 
    -0.1360601, -0.1581406, -0.1773318, -0.1942818, -0.2120507, -0.2328623, 
    -0.2486207, -0.2574944, -0.2643331,
  -0.242878, -0.2432954, -0.2456371, -0.2484859, -0.246711, -0.2356653, 
    -0.2188942, -0.1971849, -0.1748047, -0.1509389, -0.1266001, -0.1006486, 
    -0.07961553, -0.05946203, -0.04335558, -0.02576862, -0.01072463, 
    0.00548546, 0.01795508, 0.03147414, 0.04159647, 0.05174687, 0.05980271, 
    0.07020059, 0.07642132, 0.08303048, 0.08744278, 0.09412728, 0.09381769, 
    0.09012906, 0.08609121, 0.08380342, 0.08335783, 0.08396182, 0.07919189, 
    0.07342222, 0.06718788, 0.06545076, 0.05878308, 0.04630405, 0.03419991, 
    0.02710448, 0.01961072, 0.01391637, 0.007004872, 0.0001507849, 
    -0.01083602, -0.01842642, -0.02468623, -0.03130272, -0.04600386, 
    -0.03945367, -0.004812449, 0.04677442, 0.07119467, 0.07707117, 
    0.05672957, 0.05068462, 0.02700494, 0.01551126, 0.02542634, 0.009864196, 
    0.01425382, 0.0355641, 0.05173864, 0.05795661, 0.0483937, 0.03662974, 
    0.02634078, 0.03406377, 0.05286391, 0.06695324, 0.07734853, 0.03568792, 
    0.1198956, 0.1579804, 0.1566737, 0.1604327, 0.157091, 0.155894, 
    0.1430632, 0.1280777, 0.1065456, 0.08495188, 0.0638735, 0.04520851, 
    0.0229768, 0.003173565, -0.01512593, -0.0231936, -0.02187508, 
    -0.02424207, -0.03013486, -0.0320598, -0.03015676, -0.02550441, 
    -0.01888207, -0.009394851, -0.0005474817, 0.008666852, 0.01625053, 
    0.02316435, 0.0300911, 0.03934889, 0.04720897, 0.05426628, 0.06181527, 
    0.06705713, 0.0636059, 0.0558332, 0.04614645, 0.03417978, 0.01861827, 
    -0.0002066307, -0.02202447, -0.04518019, -0.07188839, -0.0962236, 
    -0.1169079, -0.1371394, -0.1530512, -0.1723848, -0.1964168, -0.2135817, 
    -0.2225379, -0.2285196, -0.2358452, -0.2403804,
  -0.2412046, -0.2338702, -0.2262463, -0.2188575, -0.2119946, -0.2041207, 
    -0.1923768, -0.1779403, -0.1593175, -0.1380354, -0.1165751, -0.09826659, 
    -0.0802108, -0.0608165, -0.04148354, -0.02231558, -0.005784489, 
    0.01002957, 0.02290723, 0.03470793, 0.04367176, 0.05449195, 0.06311578, 
    0.0694203, 0.0748465, 0.08359896, 0.0918639, 0.09847495, 0.09473731, 
    0.08877335, 0.08592775, 0.08500658, 0.08198053, 0.08186601, 0.08087175, 
    0.07864016, 0.07143015, 0.06539883, 0.057971, 0.04868349, 0.03730169, 
    0.0292768, 0.02142617, 0.01456633, 0.00498423, -0.003897607, -0.01478827, 
    -0.02565992, -0.039386, -0.04904991, -0.05777943, -0.06967025, 
    -0.09049389, -0.09936452, -0.09441677, -0.06447262, -0.04521224, 
    -0.007901743, -0.002257399, 0.01098823, 0.03214752, 0.02690712, 
    0.02625864, 0.04337574, 0.04929261, 0.04701626, 0.03069849, 0.02030004, 
    0.01134213, 0.02927718, 0.03512017, 0.0575794, 0.04362236, 0.03033713, 
    0.140477, 0.1513034, 0.1546403, 0.1630426, 0.1641177, 0.1556113, 
    0.1443275, 0.1271966, 0.1071773, 0.0847376, 0.06165832, 0.03843516, 
    0.02258301, 0.008365706, -0.001961067, -0.01642253, -0.03126873, 
    -0.03476782, -0.02891791, -0.0245428, -0.02087201, -0.01809815, 
    -0.01388477, -0.009063542, -0.002286196, 0.006910726, 0.01924177, 
    0.03187155, 0.04407697, 0.05368875, 0.06284651, 0.06942903, 0.06936923, 
    0.06501988, 0.06186511, 0.05829902, 0.05050664, 0.03819123, 0.02274035, 
    0.00386155, -0.01936213, -0.04572915, -0.06994218, -0.09470642, 
    -0.1192371, -0.1388523, -0.1583892, -0.1716903, -0.1834458, -0.2011016, 
    -0.2215887, -0.2383804, -0.245553, -0.2461771,
  -0.243798, -0.2394235, -0.232523, -0.225227, -0.214505, -0.2022953, 
    -0.1874897, -0.1712262, -0.1537491, -0.1379698, -0.1199314, -0.100143, 
    -0.07877148, -0.05900517, -0.03958981, -0.02212755, -0.005513322, 
    0.009024676, 0.02174622, 0.03381965, 0.04562879, 0.05516242, 0.06262143, 
    0.07115465, 0.07919027, 0.08605273, 0.09036745, 0.09391402, 0.09221247, 
    0.08877502, 0.0861662, 0.08409591, 0.08511398, 0.08619856, 0.08248749, 
    0.07623109, 0.07016127, 0.06762058, 0.06087112, 0.04735917, 0.03558612, 
    0.02773154, 0.02047509, 0.01335642, 0.005191594, -0.004914105, 
    -0.01681781, -0.02862135, -0.04030439, -0.05419564, -0.07153335, 
    -0.08535308, -0.09285265, -0.1025028, -0.1199715, -0.1426238, -0.1632937, 
    -0.1672707, -0.1757786, -0.1691232, -0.1622899, -0.1348622, -0.1020647, 
    -0.05466643, -0.01043718, 0.03170437, 0.05679647, 0.06458701, 0.02033871, 
    -0.006117046, 0.004364908, 0.043457, 0.002435058, 0.05287012, 0.1515685, 
    0.1408897, 0.1624804, 0.1599457, 0.1560904, 0.1475285, 0.1401204, 
    0.1238067, 0.1068678, 0.0848484, 0.06627643, 0.04442054, 0.02182415, 
    0.0006969869, -0.01355927, -0.02032776, -0.01811877, -0.02360368, 
    -0.02945919, -0.03235051, -0.02865374, -0.02419278, -0.01583189, 
    -0.0070149, 0.003074542, 0.01154172, 0.02056779, 0.02703933, 0.03525836, 
    0.04325696, 0.05121157, 0.0563602, 0.06464231, 0.07037055, 0.0694076, 
    0.0618161, 0.05320906, 0.04053521, 0.02544695, 0.005716585, -0.01563787, 
    -0.04002304, -0.06711291, -0.09293172, -0.1142186, -0.1368014, -0.154433, 
    -0.1752915, -0.1965052, -0.2125403, -0.2218282, -0.2307497, -0.2399774, 
    -0.2451427,
  -0.2444127, -0.2396758, -0.2328822, -0.2248032, -0.2151943, -0.2049578, 
    -0.1918793, -0.1779274, -0.1602566, -0.140038, -0.1175891, -0.09789708, 
    -0.07720796, -0.05726181, -0.0362607, -0.01847998, -0.00135228, 
    0.01293264, 0.02728212, 0.0384244, 0.04785632, 0.05608385, 0.06573433, 
    0.07165736, 0.07770908, 0.08394309, 0.09267595, 0.09858358, 0.09622225, 
    0.08993906, 0.08882115, 0.08758517, 0.08537182, 0.08324328, 0.0819578, 
    0.07842998, 0.07253163, 0.06603473, 0.06035754, 0.05058944, 0.03985652, 
    0.0304696, 0.02314574, 0.01481959, 0.00590989, -0.00503087, -0.01649556, 
    -0.02985546, -0.04286766, -0.05634373, -0.06796923, -0.08348188, 
    -0.1017539, -0.1195111, -0.1266072, -0.1289971, -0.1328509, -0.1520287, 
    -0.1774936, -0.210407, -0.2361294, -0.2497406, -0.2510481, -0.239274, 
    -0.2172206, -0.1677275, -0.08685258, -0.005449966, 0.02285049, 
    0.004089735, 0.01217604, 0.009134002, -0.02343513, 0.09858347, 0.1487421, 
    0.1433815, 0.1578827, 0.1540689, 0.1614128, 0.1557029, 0.1461866, 
    0.1277212, 0.1069574, 0.08327979, 0.06088501, 0.04006273, 0.02628249, 
    0.01136249, -0.00196217, -0.01825362, -0.03176713, -0.03238434, 
    -0.02527028, -0.02098355, -0.01798901, -0.0156956, -0.01164989, 
    -0.006676883, 0.0003428459, 0.009632975, 0.02210206, 0.03467767, 
    0.04724689, 0.05726136, 0.06781486, 0.07587108, 0.0774402, 0.07285018, 
    0.06945375, 0.0655089, 0.05804482, 0.0452809, 0.02960464, 0.009927906, 
    -0.0136058, -0.04031473, -0.06461078, -0.09071905, -0.1164997, 
    -0.1371752, -0.1572537, -0.1717574, -0.1847667, -0.2026619, -0.2216636, 
    -0.2364625, -0.2429706, -0.2460706,
  -0.244288, -0.2406188, -0.2351528, -0.2282628, -0.2191091, -0.2066283, 
    -0.1919059, -0.1739489, -0.1556007, -0.1371617, -0.1181935, -0.09650253, 
    -0.07490122, -0.05423315, -0.03530396, -0.01777388, -0.001191862, 
    0.013349, 0.02538539, 0.03598215, 0.04732757, 0.05774986, 0.06610884, 
    0.07361138, 0.08168787, 0.08899858, 0.09399629, 0.09540898, 0.0919911, 
    0.08843543, 0.08666415, 0.083901, 0.08494468, 0.08628316, 0.08422007, 
    0.07860452, 0.07326815, 0.07002181, 0.06333244, 0.04947749, 0.03808048, 
    0.02974439, 0.02268073, 0.01495007, 0.006634474, -0.004181445, 
    -0.01613662, -0.02911702, -0.04169774, -0.05604917, -0.07214099, 
    -0.08622921, -0.09556615, -0.1075935, -0.1223248, -0.1296149, -0.123936, 
    -0.1249759, -0.1544833, -0.2073907, -0.2517191, -0.2741424, -0.270357, 
    -0.2636373, -0.2653179, -0.2754118, -0.2386662, -0.1197222, -0.002327733, 
    0.01500629, 0.0005403832, -0.05291775, 0.01426581, 0.139998, 0.1337246, 
    0.1449172, 0.1558963, 0.1618166, 0.1575158, 0.1483064, 0.1380149, 
    0.1241969, 0.1069083, 0.087376, 0.06638896, 0.04367167, 0.01878887, 
    0.0009395182, -0.01122092, -0.01524331, -0.01594096, -0.0227744, 
    -0.03035611, -0.03130856, -0.02746242, -0.02101362, -0.01308134, 
    -0.003127456, 0.00618273, 0.01581615, 0.02424034, 0.03194332, 0.03968257, 
    0.04858454, 0.05545136, 0.06032208, 0.06730756, 0.07448852, 0.0747177, 
    0.06890446, 0.06036124, 0.04826468, 0.03241432, 0.0125451, -0.009837728, 
    -0.03442875, -0.06252378, -0.08849616, -0.1113501, -0.1347443, 
    -0.1536434, -0.1748048, -0.1965039, -0.2122121, -0.2226509, -0.2314301, 
    -0.2403085, -0.2443949,
  -0.2458596, -0.2403259, -0.2336327, -0.225385, -0.2162865, -0.2053751, 
    -0.192055, -0.1767912, -0.1588025, -0.1371804, -0.1144938, -0.09310007, 
    -0.07283725, -0.05217971, -0.03229129, -0.01399034, 0.001786806, 
    0.01595978, 0.02938209, 0.04206863, 0.05188265, 0.05997556, 0.06743934, 
    0.07364805, 0.07981576, 0.08590314, 0.0927615, 0.09817905, 0.09591365, 
    0.09094383, 0.08977461, 0.08961554, 0.08781962, 0.08615017, 0.08398196, 
    0.08006904, 0.07354495, 0.06738222, 0.06197363, 0.05293205, 0.04155207, 
    0.03221166, 0.02435637, 0.01625919, 0.006809443, -0.004057884, 
    -0.01635551, -0.02936307, -0.04281902, -0.05602878, -0.06891298, 
    -0.08323085, -0.09876877, -0.1115779, -0.1220338, -0.1278329, -0.1166585, 
    -0.09184331, -0.08610485, -0.1209277, -0.1834247, -0.2520379, -0.2998728, 
    -0.3045812, -0.2902858, -0.2984114, -0.3083416, -0.2295054, -0.09132567, 
    -0.02037908, -0.06541967, -0.05046435, 0.09614872, 0.1357757, 0.1300858, 
    0.1503199, 0.1528628, 0.1553054, 0.1549674, 0.1535752, 0.1433348, 
    0.1268268, 0.1046964, 0.08271575, 0.06137925, 0.04396093, 0.02979729, 
    0.01299465, -0.003913373, -0.02002102, -0.03116222, -0.0282107, 
    -0.02090627, -0.01708615, -0.01551318, -0.0132826, -0.009605139, 
    -0.003851891, 0.003073037, 0.01297969, 0.02508515, 0.03834537, 
    0.05076018, 0.06170577, 0.07263231, 0.08280513, 0.08564442, 0.0820117, 
    0.07761914, 0.07369876, 0.06571175, 0.05310671, 0.03656714, 0.016553, 
    -0.008092746, -0.03487244, -0.05957383, -0.08609021, -0.113303, 
    -0.1346506, -0.1556493, -0.1704299, -0.1848188, -0.2031496, -0.2226197, 
    -0.2373285, -0.2444937, -0.247509,
  -0.244412, -0.2406856, -0.2349517, -0.2280661, -0.218557, -0.2058602, 
    -0.1904801, -0.1720421, -0.1525138, -0.1332503, -0.1135219, -0.09200723, 
    -0.07070215, -0.05025221, -0.03161675, -0.01414781, 0.002302298, 
    0.01744283, 0.02961341, 0.0396587, 0.04907923, 0.05892505, 0.06774777, 
    0.07607954, 0.08360518, 0.09096707, 0.09632049, 0.09768347, 0.09315039, 
    0.09000419, 0.0887783, 0.08647138, 0.08640888, 0.087185, 0.08478093, 
    0.07981083, 0.07491651, 0.07188603, 0.06479433, 0.05137938, 0.03983703, 
    0.0313732, 0.02382216, 0.01616082, 0.007444531, -0.003420889, 
    -0.01591814, -0.02910325, -0.04224813, -0.05618054, -0.07159099, 
    -0.08503455, -0.09528556, -0.1045332, -0.11424, -0.1277861, -0.1397062, 
    -0.1286064, -0.09547633, -0.07279614, -0.07902638, -0.1224388, 
    -0.2009089, -0.274629, -0.2995771, -0.289987, -0.2684109, -0.2027344, 
    -0.1133183, -0.100083, -0.08126349, 0.0564671, 0.1285084, 0.12046, 
    0.1363447, 0.1437018, 0.1528145, 0.1597852, 0.1584521, 0.1504486, 
    0.1398053, 0.1259625, 0.10891, 0.0882681, 0.06552422, 0.04099226, 
    0.01763058, 0.002962589, -0.006270856, -0.01096725, -0.014471, 
    -0.02379997, -0.03064182, -0.03015453, -0.02464199, -0.0175364, 
    -0.009019256, 0.0007097125, 0.01038212, 0.02005541, 0.02892601, 
    0.03664476, 0.04486063, 0.0539127, 0.06096715, 0.06509769, 0.07133535, 
    0.07858798, 0.08025098, 0.07582565, 0.06821062, 0.05631551, 0.04023213, 
    0.01958014, -0.003719434, -0.02945065, -0.05810565, -0.08406848, 
    -0.107638, -0.1325478, -0.1522276, -0.1740721, -0.1957248, -0.2113318, 
    -0.2220295, -0.2314582, -0.2405072, -0.2447402 ;
}
