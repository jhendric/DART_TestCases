netcdf sampling_error_correction_table {
dimensions:
	bins = 200 ;
	ens_sizes = UNLIMITED ; // (40 currently)
variables:
	int count(ens_sizes, bins) ;
		count:description = "number of samples in each bin" ;
	double true_corr_mean(ens_sizes, bins) ;
	double alpha(ens_sizes, bins) ;
		alpha:description = "sampling error correction factors" ;
	int ens_sizes(ens_sizes) ;
		ens_sizes:description = "ensemble size used for calculation" ;

// global attributes:
		:num_samples = 100000000 ;
		:title = "Sampling Error Corrections for fixed ensemble sizes." ;
		:reference = "Anderson, J., 2012: Localization and Sampling Error Correction in Ensemble Kalman Filter Data Assimilation. Mon. Wea. Rev., 140, 2359-2371, doi: 10.1175/MWR-D-11-00013.1." ;
		:version = "$Id: gen_sampling_err_table.f90 10966 2017-01-27 21:14:27Z nancy@ucar.edu $" ;
data:

 count =
  1597443, 1336022, 1200480, 1106023, 1030861, 972969, 922597, 880032, 
    840077, 810628, 780319, 755222, 728582, 707971, 688830, 670002, 651611, 
    637303, 622960, 608345, 595763, 583701, 573152, 561961, 551450, 541395, 
    533883, 523983, 517067, 507927, 501521, 493281, 486655, 480179, 474162, 
    469790, 462548, 457518, 451755, 447751, 442642, 438724, 434552, 429324, 
    426324, 422144, 418222, 413142, 410063, 406672, 404270, 401244, 399292, 
    396085, 392425, 389736, 387118, 384062, 382936, 380106, 377839, 375125, 
    373430, 370618, 371437, 366872, 366386, 364311, 362291, 361218, 360412, 
    357323, 357354, 355078, 354541, 353334, 352844, 350874, 349810, 348949, 
    348504, 347104, 346817, 344990, 344833, 345203, 343921, 344281, 341320, 
    342485, 339724, 340870, 340190, 340410, 340089, 340126, 339594, 339141, 
    340196, 339001, 339465, 339191, 340676, 339825, 339206, 339123, 340907, 
    340090, 340478, 340995, 342060, 342267, 342485, 343850, 344335, 344205, 
    345677, 347167, 347476, 347809, 347715, 349572, 352065, 351654, 352651, 
    355535, 355156, 357330, 358644, 359525, 361634, 362512, 364634, 365521, 
    368528, 369845, 371752, 373509, 375850, 378495, 380853, 382195, 384280, 
    387926, 389814, 392269, 395760, 397738, 401415, 404167, 407958, 411061, 
    414237, 417695, 422107, 425929, 429880, 433992, 436494, 442025, 446567, 
    452891, 458344, 462808, 469911, 473802, 480376, 486682, 493448, 500560, 
    508337, 516375, 523210, 533415, 541889, 551070, 562490, 572515, 583785, 
    593864, 608883, 622486, 636488, 652805, 669958, 689178, 708027, 730840, 
    752414, 779125, 809445, 841651, 880976, 921879, 973631, 1030331, 1106657, 
    1201415, 1335930, 1596685,
  1165953, 1066496, 997563, 944768, 901188, 864915, 831589, 803190, 779830, 
    755067, 734672, 714786, 695829, 680723, 668120, 651272, 638022, 625890, 
    614042, 601486, 593161, 581888, 575212, 563624, 556144, 550696, 539817, 
    534110, 526243, 518643, 513616, 507553, 502015, 497580, 491026, 484979, 
    480294, 475832, 471163, 467551, 463284, 459198, 455438, 451819, 448516, 
    445126, 440184, 437960, 434734, 432249, 430020, 424676, 422704, 418608, 
    418427, 415328, 411951, 411080, 409603, 406541, 403956, 404009, 399164, 
    398160, 396003, 394378, 392864, 389606, 390333, 388602, 386404, 386458, 
    383796, 383882, 382120, 380732, 378480, 378846, 378284, 377107, 376805, 
    376349, 373766, 374300, 374299, 372143, 372545, 370858, 369163, 370601, 
    370101, 369185, 368602, 367970, 368996, 368706, 369043, 367289, 368483, 
    368477, 367978, 368634, 368388, 368660, 368077, 367897, 370563, 368564, 
    369972, 370340, 370532, 371428, 370944, 372630, 372586, 372468, 374058, 
    374044, 376029, 375128, 377009, 378117, 378917, 379939, 381515, 382202, 
    383947, 384283, 385820, 387221, 388558, 390109, 391823, 392261, 394114, 
    395987, 397914, 399735, 403553, 404311, 406149, 407777, 409842, 412764, 
    415059, 417115, 419790, 422599, 425408, 428198, 431808, 434900, 438079, 
    441043, 443664, 448000, 453878, 454838, 460172, 461636, 466804, 471047, 
    477080, 481999, 486902, 492529, 496207, 501438, 506328, 514012, 518979, 
    527086, 533834, 540614, 549171, 556078, 564576, 574055, 583711, 592497, 
    603331, 613389, 626785, 639106, 652694, 665332, 682935, 697202, 716283, 
    733288, 756341, 778418, 803572, 831206, 865276, 901263, 945364, 998632, 
    1064811, 1165991,
  967723, 918106, 876435, 845427, 816014, 794005, 769038, 748140, 731341, 
    712928, 699097, 683540, 669946, 657031, 645014, 633600, 623505, 612497, 
    604825, 594953, 586190, 578597, 569807, 562139, 555413, 549195, 542381, 
    537003, 531757, 524902, 519551, 515353, 508821, 504200, 500361, 493918, 
    490155, 486394, 482471, 478310, 473477, 470421, 466511, 463271, 460457, 
    456104, 455834, 451604, 449219, 445519, 443285, 440985, 438862, 435213, 
    435364, 431447, 429655, 426519, 424590, 423280, 422777, 420329, 417924, 
    415676, 413726, 414592, 411196, 409261, 408134, 406997, 405573, 405068, 
    402654, 402368, 400427, 399839, 398988, 397760, 397931, 397020, 395117, 
    394617, 393988, 392629, 393945, 391744, 393064, 389989, 390737, 390052, 
    390024, 389434, 389308, 388287, 389250, 388760, 388966, 388074, 387252, 
    387525, 387442, 388799, 387488, 388299, 388398, 388397, 389286, 389628, 
    389850, 388965, 389648, 390265, 391376, 391445, 391847, 391415, 392847, 
    393952, 394825, 394399, 396605, 397608, 398835, 398429, 399635, 399818, 
    402914, 403239, 405602, 406272, 406338, 408322, 411099, 412485, 412410, 
    415072, 415736, 417208, 419029, 420607, 424240, 426937, 427047, 429771, 
    430855, 434362, 436362, 438484, 440605, 442929, 445655, 449199, 451313, 
    455014, 456210, 460707, 464416, 467086, 470997, 473326, 479573, 482466, 
    486642, 489566, 495927, 498562, 503447, 509197, 513992, 519269, 524282, 
    530189, 536582, 543030, 549910, 557003, 561242, 569316, 577939, 586329, 
    594133, 603748, 613038, 623383, 634425, 645658, 657437, 670543, 683995, 
    696961, 714426, 730516, 749359, 770002, 792333, 815929, 843828, 877575, 
    916878, 967318,
  856761, 827670, 802682, 780170, 758634, 740229, 725510, 709890, 696829, 
    681445, 669200, 657450, 647133, 636418, 626975, 618543, 609757, 601669, 
    593580, 585662, 578455, 572011, 564845, 557320, 552973, 546479, 542945, 
    535939, 530828, 526841, 521988, 516901, 512851, 507334, 504546, 498813, 
    496000, 493059, 488407, 486046, 482736, 479449, 474013, 472829, 470381, 
    466822, 462920, 460522, 458595, 455962, 453563, 452700, 449441, 446526, 
    444236, 443032, 439801, 438687, 437596, 435568, 433636, 431517, 431121, 
    428127, 427143, 426295, 423234, 422570, 422104, 419961, 419798, 418665, 
    418047, 416608, 416220, 413194, 412266, 411722, 411533, 409401, 409076, 
    409620, 409004, 406875, 407889, 406312, 406313, 404640, 404396, 403846, 
    404048, 404076, 404122, 404161, 402807, 402760, 403130, 402703, 401776, 
    403365, 403170, 402211, 402699, 403365, 403349, 403890, 403970, 403824, 
    404492, 404805, 405193, 404510, 405272, 405243, 407030, 407528, 406990, 
    408198, 407946, 409144, 410201, 413724, 411346, 413362, 414153, 414994, 
    414578, 416168, 418416, 418844, 421136, 420848, 422040, 424298, 425453, 
    427490, 427863, 431119, 432778, 434292, 435732, 436325, 438976, 439414, 
    443473, 444495, 446768, 449720, 450993, 453091, 455769, 458338, 461156, 
    464906, 467155, 469626, 472132, 475804, 479347, 483044, 484908, 489048, 
    491014, 496826, 500433, 503808, 506797, 512564, 516569, 521870, 526343, 
    530426, 536473, 541724, 546472, 552266, 558709, 566575, 571926, 578510, 
    586142, 592276, 600324, 607646, 618121, 627152, 639068, 646849, 657488, 
    670310, 680147, 696212, 709650, 724640, 742573, 759888, 779902, 802376, 
    826393, 857137,
  789523, 768914, 749938, 734097, 718713, 703170, 692502, 679764, 669227, 
    658509, 648772, 638263, 628898, 621346, 613645, 604632, 598842, 590909, 
    583334, 577789, 570981, 564215, 560587, 554936, 550223, 544501, 539700, 
    535306, 531113, 524577, 521856, 518073, 511971, 511099, 506078, 501553, 
    497482, 496392, 492348, 489317, 487814, 483247, 480356, 478208, 474058, 
    472274, 469357, 468328, 465411, 463505, 460874, 458506, 457148, 454168, 
    452450, 451043, 449383, 447853, 445283, 444457, 443984, 440889, 439446, 
    437570, 436963, 436348, 434637, 434024, 431724, 430576, 428652, 426956, 
    428015, 426209, 424493, 424709, 423245, 422137, 422165, 421824, 420827, 
    419689, 418948, 418860, 417935, 417031, 416935, 417703, 415988, 415699, 
    414618, 415589, 413834, 412972, 415539, 413498, 414456, 414634, 413734, 
    413579, 413971, 414779, 415306, 413033, 415087, 413851, 414290, 415083, 
    414530, 415649, 416202, 417353, 416924, 417362, 417763, 418858, 418405, 
    419368, 420361, 420003, 420813, 421970, 422830, 424003, 424410, 426586, 
    426290, 427746, 428708, 429402, 430276, 431464, 433536, 434265, 434009, 
    436443, 438017, 439203, 440946, 443172, 444149, 446035, 447684, 449302, 
    452291, 453178, 455208, 457260, 458885, 461225, 462351, 465189, 468111, 
    470289, 473183, 475217, 478197, 480578, 483263, 486251, 489309, 492919, 
    497153, 497891, 501864, 506569, 510737, 513848, 517354, 521251, 525624, 
    530145, 535476, 538672, 544310, 549328, 554374, 560117, 564787, 572982, 
    578529, 584750, 590399, 599317, 606547, 612571, 621063, 628479, 640104, 
    647986, 657741, 668533, 678956, 691462, 703855, 718888, 734671, 750949, 
    769479, 787445,
  741991, 725632, 713981, 700494, 688140, 677144, 667459, 657416, 647834, 
    639298, 630919, 623151, 613996, 608614, 601622, 594678, 588848, 582287, 
    575722, 572552, 566399, 560544, 555397, 551401, 546223, 541712, 537705, 
    533724, 529671, 526505, 521273, 517331, 513796, 511684, 508106, 503982, 
    501381, 498683, 494946, 491836, 489316, 487121, 483990, 482054, 479929, 
    477335, 475849, 471174, 470821, 468917, 466835, 464661, 462804, 461507, 
    459240, 457668, 455601, 452925, 451319, 451842, 449120, 447904, 445624, 
    445791, 443661, 442359, 441679, 438942, 440463, 438115, 437851, 436490, 
    435939, 434248, 432788, 433368, 430566, 432177, 429802, 429330, 428849, 
    429356, 427897, 427120, 426461, 425254, 426008, 424570, 426021, 424174, 
    424500, 424360, 423478, 423357, 424930, 423922, 422816, 422184, 422928, 
    422823, 422460, 421458, 423409, 422494, 423657, 422798, 424680, 422885, 
    425470, 424766, 424466, 423746, 425746, 426860, 426190, 427546, 426837, 
    427301, 428762, 428642, 429290, 431245, 431181, 431862, 432066, 433090, 
    433961, 434960, 436921, 437697, 437272, 439550, 440180, 441991, 442338, 
    443215, 443793, 447339, 447940, 449366, 451166, 453559, 453802, 454660, 
    457002, 459213, 460788, 462895, 463271, 466263, 468126, 470413, 472395, 
    474649, 476870, 479577, 481773, 484918, 486603, 489963, 492775, 495093, 
    498819, 501277, 504494, 507899, 510426, 515213, 517530, 521174, 524688, 
    529303, 533607, 538546, 542313, 544652, 549801, 555551, 560749, 565278, 
    571808, 576291, 583884, 588699, 595781, 601752, 608298, 616259, 623779, 
    630343, 637616, 648515, 658090, 667314, 676393, 688303, 700235, 713465, 
    726888, 741552,
  683225, 672087, 662605, 655640, 647252, 638872, 633003, 625288, 618534, 
    610570, 605555, 600098, 594612, 589860, 582335, 578986, 573996, 570018, 
    564055, 559303, 555168, 551679, 547013, 543713, 540602, 537449, 533403, 
    530627, 526944, 522898, 519702, 517947, 513989, 511370, 509615, 506200, 
    503622, 501610, 496585, 496289, 493825, 491423, 490098, 486315, 484995, 
    482803, 481200, 478882, 478730, 475679, 474219, 472366, 469130, 469002, 
    467351, 466842, 465103, 462385, 462268, 460366, 459782, 457871, 457612, 
    456261, 454118, 453453, 453401, 451232, 449059, 450123, 449356, 447300, 
    447717, 446872, 446145, 443979, 443590, 442988, 442549, 441057, 441154, 
    440987, 440763, 438616, 440311, 438035, 439228, 440109, 438255, 437261, 
    436590, 437672, 436644, 438156, 437105, 435863, 435265, 435695, 436149, 
    435384, 434897, 436188, 433594, 437143, 436735, 437038, 436431, 437023, 
    437239, 438841, 437522, 437712, 437918, 438810, 438724, 440046, 440021, 
    440058, 440885, 440558, 442728, 442485, 442682, 443991, 444127, 444557, 
    446135, 446303, 447777, 447931, 449860, 450564, 451689, 452295, 453599, 
    453638, 456494, 458548, 457545, 458290, 461491, 462659, 462474, 463686, 
    465671, 470040, 470611, 470801, 471674, 474366, 474506, 477063, 478991, 
    481814, 483019, 486790, 486307, 488868, 491690, 493214, 497060, 497049, 
    501499, 502663, 506598, 508943, 510861, 515427, 518301, 520420, 523986, 
    527222, 529624, 532977, 536788, 540300, 545062, 547920, 552241, 557742, 
    559846, 565905, 569463, 573069, 579245, 582907, 588613, 593911, 599958, 
    604886, 611442, 618163, 623648, 631056, 640071, 647492, 655981, 662833, 
    672425, 683038,
  646514, 639812, 632502, 627221, 619617, 614082, 609391, 603873, 599077, 
    593006, 588342, 584959, 580683, 574972, 570093, 565898, 563505, 560087, 
    555471, 551741, 548872, 544347, 541384, 537552, 536290, 532723, 529778, 
    527355, 522131, 522166, 517831, 516376, 512609, 511899, 507790, 507470, 
    503299, 502782, 500832, 499037, 495512, 493637, 492011, 491058, 488731, 
    486613, 484509, 482594, 482219, 480284, 479873, 477528, 476653, 475271, 
    473881, 471335, 471057, 469147, 467702, 467217, 464782, 464794, 463433, 
    461873, 461465, 460832, 460296, 459602, 458442, 458861, 456324, 456079, 
    453938, 453095, 454092, 453389, 453846, 451405, 452284, 449775, 450813, 
    450101, 448724, 448905, 448598, 447614, 449318, 446519, 447319, 447933, 
    446532, 446381, 446292, 446107, 445715, 445080, 444940, 445761, 445217, 
    445098, 446300, 447281, 445232, 445863, 444509, 445659, 445459, 445386, 
    446603, 447247, 446116, 445700, 446761, 446859, 448090, 448426, 449150, 
    449646, 449207, 449855, 450852, 451011, 451525, 452677, 453086, 453008, 
    453582, 454630, 455255, 457036, 458005, 458758, 458723, 461028, 460670, 
    461689, 462782, 464184, 464665, 466128, 466711, 467660, 469982, 469792, 
    473006, 473899, 474408, 474606, 477434, 479453, 479890, 481862, 482275, 
    485075, 487700, 488434, 491240, 491851, 494632, 497158, 497884, 499639, 
    501767, 504285, 506848, 508681, 511664, 513285, 515233, 519751, 521709, 
    524225, 527265, 529738, 532004, 536564, 538732, 541129, 545203, 548162, 
    552035, 554916, 557872, 563283, 566526, 570727, 574626, 579708, 584064, 
    591109, 593911, 597751, 602700, 608019, 614770, 621891, 626422, 631935, 
    640366, 646114,
  632668, 627224, 622887, 615207, 609180, 605958, 601045, 594191, 591117, 
    584910, 582184, 578347, 573188, 570014, 566206, 561801, 557814, 556544, 
    552772, 547978, 545189, 539817, 540440, 536684, 533788, 530195, 527638, 
    525235, 522897, 520792, 517624, 514500, 512011, 510730, 508516, 506774, 
    504816, 502180, 500580, 498041, 496839, 495455, 493104, 492014, 489298, 
    487873, 486210, 484120, 483854, 482012, 480520, 479766, 478507, 477730, 
    476219, 475043, 472317, 471184, 470089, 470198, 469602, 467061, 466199, 
    465758, 464237, 464479, 463099, 462485, 460305, 460478, 459930, 459596, 
    458553, 459398, 457115, 457271, 456435, 454693, 454296, 454216, 453929, 
    452645, 452734, 451610, 451623, 451524, 451004, 450267, 449359, 450669, 
    450414, 450717, 449828, 449351, 449920, 449722, 449044, 449229, 449336, 
    448553, 449395, 451185, 449906, 448630, 450292, 448811, 449689, 449715, 
    450565, 449881, 450028, 450187, 451102, 451812, 452140, 452158, 452463, 
    451579, 453621, 454206, 453641, 454754, 454980, 456258, 457054, 456997, 
    458721, 457970, 458759, 458905, 458849, 461477, 461991, 461987, 464359, 
    463569, 465126, 466868, 467638, 469444, 469785, 470282, 472146, 471573, 
    474745, 476057, 476400, 478662, 479730, 479996, 482417, 483422, 485369, 
    488026, 487695, 489547, 490680, 494150, 495291, 496038, 499718, 500782, 
    502758, 505451, 505489, 508618, 510681, 513246, 513703, 517622, 520115, 
    522192, 524525, 527855, 530687, 533241, 537271, 540224, 541396, 545796, 
    547936, 551576, 555422, 558086, 562815, 565950, 570579, 573125, 578193, 
    582581, 586651, 590760, 593954, 599223, 605465, 610175, 616193, 622461, 
    626851, 633192,
  622679, 617351, 611071, 606555, 599639, 597920, 592894, 588208, 585945, 
    580024, 575313, 572338, 568413, 565152, 561632, 557978, 554189, 550548, 
    547547, 546049, 543729, 540255, 536960, 534764, 532683, 528020, 525598, 
    523860, 522193, 520154, 517280, 514999, 512144, 510356, 508109, 506304, 
    505245, 501886, 500314, 499825, 497670, 495398, 494721, 491991, 491368, 
    489125, 487840, 487384, 484398, 483815, 482296, 480175, 479524, 478854, 
    476498, 476674, 474996, 475092, 471642, 472356, 470895, 468831, 468302, 
    467199, 468128, 465758, 465984, 464828, 463912, 461609, 462355, 461435, 
    461294, 459945, 460550, 458956, 459205, 457746, 458819, 457316, 456867, 
    455866, 454896, 455187, 455378, 455512, 453756, 455395, 453424, 453095, 
    452909, 453466, 453160, 452587, 453333, 452406, 451503, 452616, 452748, 
    453485, 452056, 451786, 452010, 452729, 452491, 452518, 452377, 453345, 
    452232, 453332, 453537, 455221, 454161, 453219, 455306, 455600, 455349, 
    455659, 456556, 456456, 457486, 457509, 456724, 459672, 458857, 460257, 
    460901, 461085, 460939, 463282, 463173, 463518, 464599, 465231, 467708, 
    468048, 468739, 468360, 469943, 472187, 471538, 472382, 473363, 473831, 
    476486, 477471, 479110, 480213, 479753, 482288, 484043, 485156, 485683, 
    487514, 489994, 490556, 493519, 494419, 496656, 496569, 498957, 500177, 
    504355, 504492, 507261, 509247, 511074, 512410, 515384, 516632, 518252, 
    521588, 523113, 526298, 528310, 531259, 533101, 536926, 539108, 542859, 
    545512, 548601, 551527, 555224, 557493, 561603, 564952, 568801, 571421, 
    577235, 580285, 584363, 589481, 592396, 597669, 602895, 606244, 610898, 
    616288, 623010,
  604581, 600439, 597175, 591752, 588221, 584675, 579843, 576246, 574564, 
    569076, 565825, 563143, 559994, 556284, 553432, 551109, 548585, 545667, 
    543218, 540768, 538886, 535743, 531932, 531123, 528893, 526987, 525313, 
    521257, 519122, 517752, 515691, 512851, 510994, 508753, 508219, 506130, 
    504704, 505065, 500957, 499584, 498420, 497198, 495187, 494504, 492923, 
    491758, 489914, 488048, 487011, 485995, 485701, 483047, 481978, 481709, 
    481217, 478317, 478368, 477032, 475639, 475042, 475997, 474885, 472325, 
    471070, 471614, 470153, 470442, 468728, 468134, 467738, 467112, 465980, 
    465253, 465199, 464108, 463117, 464105, 463823, 461590, 461843, 462438, 
    461265, 459921, 460128, 459038, 459888, 459006, 459828, 457755, 458023, 
    458623, 459368, 458116, 458131, 458181, 457801, 457488, 457920, 459547, 
    458015, 457808, 457035, 457058, 457438, 458473, 459517, 458347, 458635, 
    458414, 458102, 458453, 459705, 458161, 460062, 459910, 461324, 459633, 
    462620, 460946, 460618, 461022, 461929, 462857, 463856, 464163, 465121, 
    464854, 466043, 466532, 466486, 467599, 467756, 469421, 469608, 469892, 
    472209, 472053, 473272, 473557, 475462, 476157, 475453, 477560, 477952, 
    479283, 481430, 481700, 483341, 483264, 485396, 484669, 486718, 487943, 
    489798, 491564, 493702, 494433, 495530, 495950, 498032, 499708, 502181, 
    503493, 503811, 507723, 508163, 509520, 512182, 512906, 516001, 518265, 
    518956, 521051, 524749, 527340, 528930, 530401, 534065, 534915, 537383, 
    539986, 542544, 545846, 548309, 551029, 553765, 556928, 559367, 562742, 
    566571, 569805, 573503, 577846, 579924, 584973, 588833, 592355, 595958, 
    600641, 604248,
  592031, 587597, 585681, 580684, 578638, 573660, 571259, 568807, 565233, 
    562243, 559078, 556346, 552795, 551387, 549001, 545050, 543485, 541398, 
    538882, 535602, 534002, 531903, 529361, 527987, 525891, 524163, 522329, 
    520196, 517762, 516464, 513997, 513016, 510361, 509109, 507962, 505786, 
    504269, 502938, 501524, 500915, 498402, 498660, 495866, 495534, 493086, 
    493889, 491446, 489646, 488537, 487892, 487056, 485204, 483718, 483836, 
    482767, 482146, 480172, 479973, 480241, 477823, 477452, 476909, 475919, 
    474752, 474129, 472221, 472830, 472382, 471555, 470976, 469458, 469183, 
    469123, 468845, 468887, 467185, 468338, 466804, 467477, 465847, 465370, 
    464958, 464105, 464652, 464375, 463440, 464208, 463336, 463360, 463289, 
    462629, 463407, 461715, 461351, 463338, 462727, 461846, 461482, 460785, 
    462325, 462300, 462137, 462815, 462752, 462293, 463466, 462635, 462446, 
    463114, 463123, 463370, 463840, 463124, 464698, 465025, 464144, 462794, 
    464470, 465508, 466635, 465384, 467209, 466479, 466852, 467322, 468786, 
    470180, 469474, 470080, 470172, 470334, 471721, 470515, 472932, 473259, 
    473635, 474721, 475755, 476778, 477491, 478189, 479823, 479601, 481599, 
    481924, 483274, 482132, 484090, 485504, 487276, 487143, 487750, 490057, 
    491700, 493016, 492013, 493601, 496441, 497946, 497736, 499784, 502482, 
    502996, 505712, 506531, 508312, 508517, 511010, 512811, 514386, 515938, 
    518557, 519561, 522162, 524814, 525762, 527993, 529821, 532216, 535427, 
    536551, 538342, 541505, 545046, 545495, 547293, 550980, 553644, 555133, 
    558980, 560583, 563990, 568817, 570128, 575828, 578760, 581432, 584073, 
    588907, 591481,
  581951, 579670, 575338, 571880, 568474, 566734, 562165, 560789, 558385, 
    556659, 554821, 550596, 548325, 547114, 544213, 542090, 538646, 536719, 
    533906, 532506, 532092, 528826, 527250, 525662, 522994, 522026, 519688, 
    518561, 515974, 515549, 513412, 511356, 511539, 508745, 506618, 505014, 
    504101, 502967, 502797, 501032, 500020, 498211, 497019, 495541, 494960, 
    493436, 491778, 490415, 490593, 488947, 487975, 485985, 486099, 484284, 
    484177, 484873, 482643, 481722, 481238, 479479, 480457, 478146, 478840, 
    478385, 477176, 475688, 475085, 474085, 474399, 473714, 472963, 472942, 
    471261, 471724, 473184, 471011, 470564, 469404, 469479, 469575, 468214, 
    469078, 468025, 468093, 467285, 467716, 467730, 466068, 466150, 466664, 
    466562, 464563, 464814, 465302, 465126, 465674, 465146, 465566, 465530, 
    466915, 466098, 465692, 466603, 465200, 466186, 466691, 465660, 465930, 
    466849, 466651, 467744, 466965, 466744, 467292, 466509, 469439, 467482, 
    469216, 468462, 467944, 470359, 469998, 469925, 470498, 470572, 471532, 
    470303, 471363, 472347, 474324, 473956, 474548, 474507, 475142, 475834, 
    477894, 477184, 477170, 479878, 479315, 481614, 481743, 481311, 481281, 
    482872, 484322, 484709, 485303, 487641, 487471, 490261, 491838, 491443, 
    492850, 493453, 494243, 495657, 496504, 499029, 500224, 501022, 501399, 
    504305, 505062, 506321, 508072, 508449, 510386, 510629, 513126, 513379, 
    516778, 517017, 520608, 521173, 524586, 526505, 526534, 529776, 531288, 
    532736, 534336, 537955, 539362, 541841, 542664, 546192, 548216, 550333, 
    551509, 555272, 559315, 560587, 564091, 565543, 568627, 573535, 575945, 
    578702, 582166,
  573945, 571005, 567505, 565250, 562951, 559466, 557334, 555284, 552154, 
    550774, 548875, 545555, 544534, 543687, 539948, 537288, 536550, 533172, 
    532194, 529311, 528034, 525632, 524211, 524103, 520183, 520700, 517749, 
    517515, 516192, 515421, 513283, 512171, 510653, 508081, 505552, 506614, 
    504097, 503385, 501693, 501693, 499099, 497792, 498573, 496458, 493250, 
    493314, 493373, 492500, 491568, 489780, 489378, 489662, 487093, 485556, 
    487640, 485502, 482927, 484200, 483220, 482368, 480891, 480376, 480201, 
    480364, 479892, 478339, 478913, 477559, 477240, 476129, 475156, 474256, 
    473731, 474089, 473354, 472575, 472696, 473351, 473490, 470916, 471458, 
    471737, 469867, 470751, 469310, 471307, 469509, 471061, 467896, 470445, 
    471004, 469223, 468031, 468328, 467967, 468339, 467613, 469253, 469759, 
    467674, 469600, 468155, 467828, 468066, 468638, 469283, 468005, 470303, 
    467907, 469623, 468756, 468935, 468981, 468898, 470423, 472187, 470045, 
    470935, 470820, 471495, 470826, 471637, 472536, 473387, 472624, 474010, 
    473681, 475592, 474623, 475079, 476609, 477846, 475900, 478037, 479838, 
    478854, 480599, 480458, 481465, 481733, 482278, 482634, 484325, 484966, 
    485027, 485375, 487965, 487218, 488233, 489232, 489941, 491239, 491841, 
    491852, 493685, 494702, 497335, 496318, 498660, 500027, 499954, 502782, 
    502215, 505073, 505930, 508240, 507892, 509401, 511360, 511687, 514850, 
    515382, 517421, 517811, 519780, 521307, 523296, 525457, 527234, 528457, 
    530063, 531898, 532660, 535583, 537455, 539618, 541696, 543621, 546766, 
    548857, 551072, 553569, 555329, 557690, 559559, 563486, 564329, 568338, 
    571597, 573167,
  561955, 558187, 557562, 554594, 551969, 551328, 548104, 546239, 544788, 
    542060, 540610, 539195, 537526, 535803, 535320, 532742, 529238, 527207, 
    527541, 526958, 524651, 523303, 522405, 518585, 519319, 517775, 515333, 
    515998, 512888, 511317, 512030, 509507, 509012, 507283, 506551, 505537, 
    503383, 503087, 502700, 501327, 499782, 499513, 496929, 497532, 494688, 
    495197, 494189, 493700, 493551, 492128, 491942, 490837, 488928, 487340, 
    488679, 487657, 487140, 486982, 486108, 484349, 484023, 484127, 483815, 
    482560, 482198, 482631, 481347, 480693, 479162, 479140, 478815, 478916, 
    479250, 477558, 477176, 477548, 476517, 477991, 474743, 475390, 474434, 
    476029, 475605, 474562, 474302, 474263, 475305, 473911, 473742, 474028, 
    474634, 473315, 472714, 473699, 473961, 473690, 472903, 473103, 472504, 
    474949, 473442, 472118, 472750, 473126, 472327, 473024, 472745, 473517, 
    473681, 473297, 473515, 472879, 474827, 474163, 474595, 474459, 475389, 
    474127, 475283, 476215, 477148, 475741, 477202, 477142, 476912, 478683, 
    478092, 478575, 478709, 478869, 478893, 480915, 481419, 480947, 480578, 
    480984, 483320, 481335, 483649, 484773, 484464, 485129, 486025, 485785, 
    487727, 488284, 489545, 489139, 490549, 491569, 493489, 490450, 495056, 
    495270, 495797, 496108, 497019, 497659, 498644, 499995, 500848, 501943, 
    503277, 503195, 505395, 506115, 507136, 509069, 509705, 511053, 512622, 
    513901, 514884, 516490, 516721, 518767, 519868, 522239, 522326, 524129, 
    526050, 526692, 529494, 530468, 531877, 534266, 534625, 537847, 539641, 
    540704, 543036, 544099, 547221, 548708, 551124, 551939, 555079, 556181, 
    559411, 561445,
  556494, 555071, 552254, 549130, 549617, 547303, 544456, 543819, 541679, 
    539957, 537946, 537102, 534996, 532559, 531215, 529307, 528596, 526676, 
    525561, 524268, 523758, 520716, 520167, 518539, 516640, 515172, 515964, 
    513290, 512286, 510418, 509900, 510127, 509017, 506077, 505909, 504590, 
    505272, 503302, 502144, 501669, 501197, 499080, 498366, 498403, 498314, 
    495367, 494155, 494691, 493788, 491812, 492490, 491494, 488557, 488720, 
    489155, 488280, 487993, 487878, 486867, 485015, 485132, 485344, 483925, 
    483783, 482795, 483074, 482814, 481669, 480523, 480362, 481776, 480707, 
    481430, 478977, 479571, 478295, 478191, 478372, 477603, 477808, 477018, 
    478351, 475731, 476997, 476577, 475766, 477157, 476214, 475376, 476403, 
    475108, 475817, 475460, 475210, 473978, 473368, 475854, 474413, 474768, 
    474144, 474615, 475581, 475785, 474480, 475661, 475286, 472914, 475028, 
    474544, 475267, 475283, 475085, 474337, 475616, 476374, 475832, 476279, 
    476045, 478369, 477818, 479066, 477911, 478611, 479201, 478916, 478291, 
    479554, 479763, 479993, 482262, 480963, 481292, 481998, 482071, 483594, 
    482176, 483213, 483873, 485197, 485706, 485975, 487222, 488156, 487345, 
    489078, 488681, 489653, 491431, 490340, 491638, 494358, 493895, 493912, 
    494268, 495765, 496279, 497289, 499178, 499438, 499975, 502214, 500752, 
    503842, 504231, 504384, 507029, 507483, 506802, 509804, 509889, 510912, 
    513843, 512983, 515371, 515537, 516921, 519352, 520220, 520796, 521953, 
    524632, 525489, 526133, 528982, 529842, 530457, 533318, 535295, 535587, 
    537064, 539394, 541923, 543916, 545472, 546226, 549888, 551496, 551461, 
    554866, 556068,
  553098, 550697, 548681, 548178, 544131, 543135, 542207, 540966, 539536, 
    536831, 536117, 533747, 531630, 530634, 529685, 528065, 525999, 524908, 
    524256, 522953, 522064, 520503, 519192, 516529, 516497, 515545, 513793, 
    512771, 511377, 510784, 509398, 507031, 507069, 506013, 505027, 504911, 
    504589, 502388, 503427, 499931, 500451, 498690, 498273, 497647, 497659, 
    495730, 495590, 496361, 493550, 493339, 492989, 492561, 490773, 491474, 
    488690, 488414, 489250, 488165, 485854, 486591, 486123, 485471, 485913, 
    484711, 483994, 484271, 484071, 483174, 481962, 482563, 483220, 482027, 
    480880, 480952, 481092, 480280, 479357, 480387, 480078, 478509, 478019, 
    479245, 477584, 478939, 478097, 477444, 477401, 478332, 477263, 477631, 
    477519, 477199, 476752, 476909, 475800, 477951, 477524, 475371, 476181, 
    476889, 476457, 476909, 475849, 476824, 476466, 477585, 475948, 475810, 
    477032, 477648, 476404, 477096, 477603, 477706, 478566, 477499, 478628, 
    478055, 478442, 478208, 478979, 480183, 479517, 479541, 479901, 479716, 
    480108, 480627, 480187, 481503, 483289, 481928, 482838, 484184, 484787, 
    483886, 485242, 486674, 486185, 487861, 486491, 487190, 488710, 489182, 
    489422, 491369, 489631, 491004, 492546, 494270, 491791, 492790, 494286, 
    496147, 495988, 496596, 497798, 498066, 498131, 499668, 500905, 501429, 
    501918, 503561, 504820, 505305, 505951, 507652, 508527, 508827, 510737, 
    510789, 514146, 513690, 516666, 515333, 517262, 519408, 519901, 521753, 
    521825, 524846, 525331, 526571, 528376, 530077, 531694, 531178, 534449, 
    535492, 536684, 538695, 539458, 541165, 542536, 545950, 547851, 549434, 
    551333, 552098,
  546074, 544632, 543351, 540632, 540021, 538553, 536180, 534766, 534766, 
    532099, 530196, 530391, 528903, 527872, 525917, 526032, 522750, 521186, 
    521027, 519374, 519693, 519160, 517000, 516011, 514137, 513908, 512063, 
    512457, 510531, 510556, 508875, 507453, 505693, 505124, 505231, 505190, 
    503446, 502313, 502381, 500291, 500329, 498559, 499004, 497433, 497715, 
    497220, 495624, 495069, 495304, 494100, 492542, 492562, 492438, 492279, 
    490158, 490580, 490881, 489604, 488562, 490254, 487279, 488721, 486587, 
    484854, 486843, 485976, 485513, 486359, 485334, 483615, 483322, 483339, 
    483554, 483152, 482754, 482657, 484289, 482200, 482165, 480645, 479342, 
    480022, 481644, 479885, 480128, 481893, 480451, 479456, 480538, 479442, 
    480236, 478715, 478836, 479560, 479798, 479584, 477849, 479447, 478198, 
    478156, 479749, 479045, 479119, 478220, 478160, 480386, 478914, 478714, 
    479755, 480017, 480084, 480072, 479360, 480921, 480033, 480306, 480746, 
    480140, 480313, 480230, 481045, 481190, 482982, 481596, 481265, 483670, 
    484169, 483861, 482755, 483895, 484317, 484607, 485684, 486283, 486256, 
    485685, 486877, 487201, 487455, 488189, 489793, 488827, 489369, 489740, 
    489480, 490237, 492721, 492544, 493850, 493751, 493669, 495658, 494403, 
    495086, 496250, 497319, 497664, 498734, 498984, 500320, 500845, 501561, 
    503143, 504518, 504686, 505165, 505461, 507480, 508938, 508090, 509669, 
    511287, 511566, 512007, 514174, 514098, 516197, 516265, 518410, 519340, 
    520557, 521364, 522755, 524451, 524633, 525146, 527972, 529198, 529713, 
    530737, 531754, 534326, 535642, 535514, 538513, 539667, 541210, 542687, 
    544551, 546254,
  540533, 540302, 537725, 536590, 536346, 534317, 532761, 530715, 530081, 
    529110, 527934, 528196, 525548, 523342, 523682, 522612, 521237, 521957, 
    518893, 519527, 517405, 516269, 513919, 513410, 512375, 513103, 512458, 
    509344, 510257, 507859, 507498, 506443, 506562, 505484, 504457, 503659, 
    504787, 501653, 502612, 500977, 500318, 501228, 497899, 498719, 497240, 
    496363, 496058, 495658, 494367, 494485, 494100, 494074, 493455, 492274, 
    492464, 491596, 491647, 491276, 490091, 489039, 490057, 487604, 488543, 
    488656, 487712, 488648, 485936, 485134, 486540, 485276, 486078, 485554, 
    484855, 484439, 483949, 484173, 483849, 482717, 483427, 482789, 484700, 
    483536, 482279, 482636, 482714, 482405, 483142, 481452, 482766, 481421, 
    481663, 480803, 481230, 481457, 481955, 480483, 481289, 479505, 481502, 
    481232, 480969, 482569, 481220, 480649, 483111, 480313, 480888, 481002, 
    482675, 482522, 482189, 481784, 484060, 481956, 481061, 481497, 484014, 
    482662, 482636, 482100, 483291, 483018, 483193, 483525, 484592, 484835, 
    484079, 485470, 484081, 485192, 486139, 485564, 487637, 487332, 487645, 
    488808, 487973, 488801, 489001, 487461, 490045, 490648, 490280, 489972, 
    491460, 492386, 492459, 493160, 493675, 493601, 494449, 495860, 496767, 
    496500, 497050, 498012, 498767, 498293, 498684, 500014, 502564, 501930, 
    502400, 504196, 504984, 507055, 505640, 506045, 505968, 507518, 509044, 
    509452, 510362, 511199, 511419, 513178, 514128, 513936, 516471, 517261, 
    518885, 518898, 520380, 520617, 522305, 522397, 524596, 524012, 525850, 
    528382, 529278, 530071, 532940, 533437, 533945, 535820, 536793, 538675, 
    539071, 540905,
  537300, 534563, 535465, 532258, 532831, 531264, 530570, 528542, 527112, 
    525869, 524301, 524915, 522706, 521920, 521366, 520184, 518425, 518438, 
    516045, 517256, 515507, 514540, 513733, 512320, 510668, 511501, 511024, 
    508944, 508418, 507565, 507721, 506036, 506382, 505448, 504358, 503845, 
    503409, 502501, 501741, 500882, 501622, 499612, 499949, 498419, 497088, 
    497513, 495894, 496127, 495140, 496850, 494222, 494636, 492859, 493545, 
    493361, 492155, 492289, 491813, 492704, 490527, 491023, 490158, 489616, 
    489211, 488962, 487795, 487797, 487248, 486943, 486645, 487144, 486886, 
    486060, 485835, 485052, 486326, 485276, 485401, 484656, 485531, 485725, 
    482716, 484698, 484253, 483991, 483854, 485102, 483847, 482767, 483489, 
    482031, 484647, 483819, 483288, 483662, 483584, 482647, 482712, 483572, 
    481645, 483309, 483697, 483761, 482936, 482328, 482613, 484181, 483341, 
    483473, 483005, 481790, 483224, 483489, 484006, 482255, 483353, 484322, 
    484698, 483523, 484106, 485596, 483787, 485314, 484634, 487235, 486361, 
    486743, 486740, 486799, 487134, 487146, 486946, 486307, 489184, 489003, 
    488831, 490605, 489592, 489942, 491034, 491491, 491285, 491123, 492526, 
    492278, 492869, 492791, 493736, 494908, 493574, 496126, 496157, 495378, 
    497116, 497345, 497989, 497980, 499110, 499984, 500036, 501346, 501080, 
    504193, 502743, 503428, 504267, 504889, 505691, 507449, 507089, 507801, 
    508164, 509628, 509989, 510921, 512503, 512552, 514807, 513897, 515509, 
    517511, 517882, 517621, 520303, 519972, 521226, 521785, 523128, 523748, 
    525145, 525019, 527099, 528116, 530198, 531244, 532191, 532895, 534294, 
    535882, 536837,
  533381, 532139, 531363, 531135, 528498, 528463, 527351, 525095, 524949, 
    524570, 523656, 521699, 520838, 520817, 519498, 519318, 517056, 515651, 
    515785, 514626, 514233, 514265, 513038, 510628, 511139, 509887, 509241, 
    508121, 508784, 508417, 506501, 505250, 505262, 504545, 504534, 504282, 
    503708, 501335, 501738, 500826, 500177, 500338, 500026, 498279, 497217, 
    497246, 496358, 496427, 496628, 495323, 495961, 495357, 494696, 494162, 
    492736, 492854, 493426, 491833, 492937, 492413, 491214, 491043, 490276, 
    490149, 490428, 488734, 489389, 489193, 488931, 488290, 487019, 488115, 
    487611, 488086, 485688, 487654, 486153, 486713, 487401, 486939, 485900, 
    485288, 484885, 485931, 485607, 485531, 484594, 484742, 483539, 486067, 
    484063, 484450, 484191, 484991, 484511, 484115, 483052, 484083, 483687, 
    484554, 484432, 484743, 484979, 484744, 484089, 484695, 484055, 484235, 
    484575, 483921, 484863, 486084, 484862, 486413, 484796, 484767, 485133, 
    485770, 485831, 486533, 486075, 486449, 485807, 485942, 488218, 487076, 
    486611, 487378, 487509, 487776, 488749, 488232, 488191, 488634, 489792, 
    489475, 489393, 491110, 491451, 490773, 492086, 492778, 493169, 492757, 
    492644, 492703, 493901, 495275, 495238, 495666, 496368, 495755, 497048, 
    496905, 497355, 498445, 498900, 499338, 499361, 500658, 501951, 501836, 
    501676, 503739, 504698, 503469, 505429, 505788, 505969, 506172, 507917, 
    507954, 508318, 509069, 509698, 511483, 512104, 510936, 513079, 513283, 
    514189, 516916, 518209, 518012, 518713, 518794, 521693, 520421, 521008, 
    522434, 524438, 523921, 526729, 525569, 528012, 529327, 530747, 530769, 
    532820, 533376,
  532388, 532193, 531065, 529030, 527858, 527110, 525759, 525042, 524888, 
    525342, 522886, 521494, 520040, 519813, 519588, 517655, 516924, 516080, 
    515593, 514109, 514336, 513022, 511674, 511172, 510536, 511355, 509263, 
    509220, 508413, 505680, 506591, 506632, 504375, 505531, 505038, 503270, 
    503031, 501824, 501305, 500935, 501417, 499959, 499094, 497484, 498779, 
    496493, 496801, 495922, 497093, 496024, 495646, 495162, 494210, 494418, 
    494035, 492653, 492717, 492318, 492604, 492057, 491451, 490579, 490893, 
    490449, 489523, 491189, 489650, 489186, 488968, 490429, 489427, 488636, 
    487198, 487271, 486641, 486393, 486111, 485990, 486309, 486171, 487417, 
    487200, 486322, 486491, 484667, 484456, 485329, 486300, 485155, 484638, 
    485048, 483765, 485185, 485266, 485017, 485153, 485247, 484464, 483776, 
    484607, 486015, 483881, 485123, 483531, 483752, 484532, 485040, 485139, 
    485254, 485633, 484016, 485614, 485070, 485072, 484505, 485065, 485534, 
    485282, 485512, 486949, 486217, 486409, 486721, 487657, 487746, 487994, 
    488725, 488068, 488546, 488634, 488553, 488392, 490161, 489609, 488873, 
    490591, 488986, 489503, 490226, 491407, 491773, 492096, 492349, 493526, 
    494406, 493934, 493894, 492874, 495231, 496799, 495016, 496001, 497217, 
    497277, 498632, 498005, 498849, 499388, 500215, 500007, 500796, 501606, 
    501373, 502939, 503063, 503811, 505245, 504983, 505224, 506705, 507494, 
    507939, 508751, 510175, 510026, 510815, 511924, 511735, 512314, 514095, 
    515208, 515517, 516514, 516667, 519552, 519549, 519815, 520711, 520900, 
    521335, 523212, 526239, 525743, 525154, 527636, 529200, 528637, 531245, 
    531298, 532915,
  532119, 530993, 530881, 528873, 526962, 526282, 525913, 525567, 524593, 
    523641, 521766, 521559, 520771, 518568, 517172, 518348, 516153, 515429, 
    515014, 515006, 513117, 512406, 512027, 511759, 511270, 509220, 509665, 
    508887, 508404, 507875, 506132, 506438, 503995, 504509, 503489, 503053, 
    502473, 502897, 502656, 500371, 499621, 500612, 499685, 498192, 498633, 
    497384, 497784, 497356, 495707, 496322, 496039, 495830, 493182, 493445, 
    493710, 493777, 491868, 492170, 494228, 491859, 491818, 489784, 490924, 
    489572, 490243, 490367, 489562, 489849, 489170, 488629, 489841, 488156, 
    488144, 487194, 488307, 487437, 487444, 488408, 487081, 486298, 486361, 
    485792, 486210, 486839, 485487, 485970, 484739, 486204, 485562, 486098, 
    484563, 484741, 486872, 484701, 484216, 485542, 483408, 485397, 484689, 
    485236, 484504, 484516, 485197, 484459, 486409, 484390, 486115, 484432, 
    485291, 486046, 486814, 484622, 485805, 485721, 485687, 485314, 486073, 
    487613, 486436, 485675, 486515, 486393, 486611, 487367, 487166, 487189, 
    489160, 488503, 487714, 488309, 488073, 488938, 488555, 489570, 489809, 
    489588, 489913, 489927, 491314, 492123, 491820, 492229, 492995, 493476, 
    494452, 493892, 493486, 494600, 495264, 496098, 495678, 496382, 496369, 
    497556, 498320, 498456, 497370, 498999, 501306, 501618, 500792, 500849, 
    502427, 502520, 503965, 504049, 503198, 505241, 506195, 505955, 508067, 
    507797, 508437, 509960, 509814, 510628, 512417, 511090, 512433, 513370, 
    514761, 514922, 516599, 515621, 517256, 518820, 519543, 520648, 521097, 
    523161, 521875, 523589, 524620, 526284, 527907, 527123, 529244, 529734, 
    531198, 532059,
  530695, 529787, 529052, 527969, 524658, 526432, 525098, 523273, 524247, 
    521750, 520523, 520858, 519524, 518505, 517161, 517971, 516952, 515896, 
    514375, 514228, 512593, 511490, 510901, 510578, 510790, 510909, 509496, 
    508720, 507748, 506816, 506851, 506371, 504367, 503471, 502982, 501982, 
    500669, 502999, 500481, 500117, 499736, 499688, 498273, 499727, 498622, 
    498902, 498029, 497173, 495636, 496442, 495578, 494575, 494855, 494267, 
    494645, 495067, 492934, 492555, 493577, 492590, 492063, 491013, 492189, 
    489799, 489480, 490819, 489244, 489735, 489618, 489574, 489242, 489482, 
    489513, 488392, 487892, 487961, 488499, 488088, 488237, 486760, 486978, 
    486889, 487977, 486456, 485722, 486336, 484748, 486388, 485767, 485524, 
    485398, 485931, 484607, 484962, 485258, 486071, 486431, 486836, 484936, 
    484716, 485252, 486040, 485334, 486435, 485025, 486537, 485766, 486615, 
    486226, 484755, 487148, 485247, 485163, 485596, 485930, 486785, 487039, 
    486470, 487042, 487291, 487444, 487475, 487724, 488495, 488356, 487154, 
    489106, 487787, 488431, 489437, 490459, 489416, 490084, 489631, 491209, 
    489772, 489909, 491002, 491613, 492348, 492601, 493826, 492050, 494027, 
    493781, 494256, 495406, 494438, 494614, 496654, 496480, 496038, 497321, 
    496728, 498290, 498419, 499815, 499418, 499526, 501057, 500132, 500369, 
    502121, 502412, 502341, 502380, 504350, 505085, 505787, 506367, 507020, 
    506962, 509386, 509329, 509241, 511587, 511351, 510525, 512350, 512233, 
    514783, 514444, 515422, 516316, 517955, 517154, 517202, 519409, 520060, 
    520582, 522835, 522650, 524037, 525364, 525952, 526421, 527965, 527756, 
    530741, 530643,
  528656, 527246, 525981, 526014, 523636, 523538, 523067, 521504, 521225, 
    521012, 520230, 519521, 517858, 516827, 516682, 515303, 514701, 514523, 
    512776, 513971, 512435, 511657, 510511, 510720, 510085, 509302, 508291, 
    506219, 506810, 505928, 504915, 505428, 504377, 503302, 504327, 503297, 
    503243, 500663, 501417, 501765, 500797, 498390, 499108, 499375, 498476, 
    498504, 497336, 496975, 497017, 497620, 496205, 494700, 494188, 495027, 
    494768, 493517, 493787, 493616, 493409, 493659, 493104, 491803, 491670, 
    491187, 491216, 490362, 490215, 491196, 489947, 491296, 490527, 490721, 
    490037, 489634, 487592, 488609, 488212, 489074, 489112, 488587, 488436, 
    488528, 487850, 488230, 487526, 487405, 486744, 487260, 486772, 488002, 
    485891, 487270, 486180, 486419, 485951, 488220, 486146, 488059, 487813, 
    485977, 485884, 486997, 486561, 484733, 486987, 486802, 487188, 486230, 
    486610, 485790, 486853, 487293, 486819, 486856, 487628, 486972, 486157, 
    487645, 490630, 488098, 488185, 487077, 489064, 487263, 487422, 489210, 
    489766, 489515, 490156, 490158, 489338, 489986, 491168, 490674, 491616, 
    491156, 491358, 491106, 493682, 493267, 492290, 492614, 494710, 495032, 
    494782, 493609, 494274, 495937, 496167, 495400, 495794, 496196, 496519, 
    497464, 498392, 497856, 498476, 500539, 499720, 500786, 500604, 501665, 
    502419, 502425, 502332, 502952, 504278, 504546, 504725, 504810, 506322, 
    507624, 507427, 506576, 508662, 510951, 510564, 510465, 511272, 510918, 
    512644, 513884, 514049, 515635, 516270, 516070, 518185, 518951, 519079, 
    519401, 520007, 521282, 523330, 523416, 522884, 525110, 525800, 526194, 
    527150, 528447,
  526007, 525830, 524212, 523842, 523612, 522720, 519307, 520726, 520786, 
    518138, 519513, 517322, 517291, 514654, 515572, 514022, 515394, 511941, 
    512602, 511343, 511612, 510330, 510786, 508908, 509024, 508994, 507119, 
    507930, 506577, 505955, 505590, 506466, 504526, 503878, 503032, 502609, 
    502025, 501363, 502276, 499344, 500387, 499862, 499617, 498005, 498517, 
    498764, 499569, 497386, 497576, 497105, 496321, 495302, 495743, 495562, 
    494769, 493496, 495269, 494444, 492791, 494120, 493280, 491430, 492093, 
    491826, 491281, 490988, 491046, 491835, 491225, 491684, 490584, 490428, 
    490588, 490132, 488984, 488929, 489389, 489070, 489792, 488658, 488721, 
    488489, 489530, 488582, 487871, 488446, 488034, 488566, 488714, 488614, 
    488659, 487415, 488164, 486780, 487577, 488325, 488139, 487203, 486972, 
    486600, 487562, 487153, 487917, 487161, 486662, 487606, 487172, 487449, 
    486085, 487687, 489138, 487857, 487696, 488603, 488983, 487292, 488831, 
    487562, 489845, 488312, 489389, 488862, 489546, 489325, 489631, 490860, 
    489928, 491110, 490105, 490655, 490065, 489193, 491750, 492150, 491196, 
    492927, 491919, 492102, 491793, 493672, 492997, 493887, 493817, 495404, 
    494412, 494182, 495324, 495510, 495054, 496742, 496829, 497772, 497588, 
    497509, 498479, 497285, 499304, 499536, 499344, 500352, 500815, 502216, 
    501494, 503708, 503442, 502321, 505244, 504699, 504158, 506124, 505080, 
    506006, 506055, 506479, 509172, 509916, 509903, 509549, 511250, 512070, 
    510611, 512838, 512968, 513287, 514165, 514974, 516098, 517218, 517334, 
    517651, 520113, 518672, 521640, 521062, 522450, 522420, 523845, 524531, 
    524532, 527385,
  524247, 523976, 522949, 523268, 521420, 520057, 520730, 519475, 519300, 
    516518, 515594, 515991, 515437, 516680, 514629, 513876, 512426, 512541, 
    512437, 511924, 510808, 508902, 509105, 508273, 508412, 506769, 508205, 
    505735, 505828, 506414, 505466, 504706, 503390, 502523, 502180, 502367, 
    502974, 501496, 501502, 501584, 501176, 499918, 499145, 499550, 499404, 
    497762, 499205, 497624, 497694, 496872, 497524, 496281, 495596, 494666, 
    495374, 494949, 495348, 493908, 495440, 495343, 493688, 492189, 493498, 
    492648, 490842, 494031, 491695, 491337, 491326, 490823, 490382, 490329, 
    491090, 490990, 491744, 490130, 490046, 489320, 489564, 488926, 489323, 
    488444, 488766, 488830, 489526, 488752, 488076, 489125, 488663, 488274, 
    489321, 488445, 488350, 487250, 488721, 487822, 488876, 487924, 488634, 
    488004, 488352, 489139, 488376, 487770, 489131, 487724, 489018, 488242, 
    487519, 487242, 488444, 488466, 488241, 489060, 488573, 488415, 490203, 
    488698, 490266, 488908, 490303, 490440, 490233, 490268, 491640, 490292, 
    490057, 491075, 490706, 491335, 492338, 491415, 492785, 491034, 490618, 
    492143, 492389, 494530, 492815, 492804, 493582, 493766, 494535, 495317, 
    494646, 494800, 495731, 495366, 496356, 496831, 496460, 498358, 498171, 
    496849, 499716, 498763, 499724, 498931, 499684, 499882, 500615, 501228, 
    502275, 502648, 503039, 504635, 502988, 505144, 504097, 504209, 504554, 
    506510, 506220, 507636, 508064, 508298, 509052, 508116, 509703, 510034, 
    512499, 512405, 511832, 513378, 514205, 513772, 516036, 514352, 516296, 
    518265, 517219, 519311, 518206, 520280, 521174, 521142, 522407, 522883, 
    523149, 525031,
  522018, 521588, 520793, 520032, 520088, 518216, 519372, 517519, 517312, 
    515871, 515612, 514158, 514575, 513436, 513366, 511574, 511096, 511935, 
    511211, 509509, 510490, 509865, 507630, 507766, 508083, 507064, 506561, 
    505499, 505960, 504462, 505129, 505577, 502838, 504237, 501691, 502359, 
    501844, 502239, 501398, 500075, 501346, 500731, 499354, 498305, 499116, 
    498788, 498532, 499144, 496695, 497476, 496683, 496780, 496975, 497034, 
    495404, 495828, 494646, 494660, 494135, 493386, 493282, 492102, 493718, 
    493717, 493835, 493610, 493584, 492393, 492896, 492056, 491450, 492041, 
    491122, 491588, 490620, 491172, 491774, 492716, 490528, 491521, 489991, 
    490173, 491125, 489854, 489031, 489635, 489909, 490207, 489967, 487632, 
    489436, 489886, 489224, 489414, 490055, 489546, 489426, 488526, 489437, 
    489031, 488804, 489673, 487888, 489497, 487359, 489179, 489390, 488626, 
    489534, 489898, 489836, 489465, 490392, 491486, 488951, 490395, 490157, 
    489140, 489708, 490753, 490791, 490039, 491086, 490741, 492290, 490319, 
    491265, 491412, 492561, 492033, 492435, 492696, 491925, 492271, 492851, 
    492917, 493153, 493325, 494431, 493670, 494413, 495064, 495118, 494300, 
    496515, 495407, 496354, 497453, 495450, 497717, 497332, 497414, 497603, 
    498066, 498618, 499769, 499273, 498754, 500373, 501184, 500073, 501371, 
    501781, 501937, 501780, 502827, 503669, 503666, 503559, 506135, 504622, 
    504937, 505943, 505476, 507056, 507654, 507552, 509480, 508839, 510816, 
    509693, 511077, 511302, 511763, 512189, 512826, 513459, 514111, 514868, 
    515399, 516699, 517438, 517323, 518480, 518268, 519997, 519218, 522061, 
    521247, 522593,
  521575, 520706, 520829, 519767, 518782, 517430, 518329, 516593, 516479, 
    515598, 515061, 515146, 512950, 513391, 512620, 512474, 511821, 511058, 
    510074, 509743, 510520, 508476, 509279, 507179, 508732, 507524, 506108, 
    503614, 505291, 505252, 504554, 506039, 503754, 503707, 503322, 501972, 
    501824, 500365, 500226, 500146, 501142, 499866, 499310, 499414, 499552, 
    498762, 497757, 496831, 497194, 496242, 498267, 497274, 495070, 496103, 
    497551, 496894, 495859, 495381, 495368, 494804, 493670, 495327, 494155, 
    492929, 492711, 493201, 492458, 493368, 492731, 491765, 492939, 492412, 
    491338, 489993, 490420, 491610, 489639, 491193, 491670, 491737, 490411, 
    491533, 489801, 490886, 490720, 490246, 489694, 489044, 490029, 490282, 
    491106, 489266, 489026, 488796, 490103, 489104, 489879, 490496, 488908, 
    489513, 489317, 489029, 489336, 489707, 489249, 489633, 490807, 489236, 
    489069, 490936, 490398, 489466, 491469, 489866, 489431, 490004, 490514, 
    490752, 490727, 490115, 490294, 491591, 490801, 492006, 489993, 492455, 
    491971, 491197, 491827, 491933, 491793, 492391, 491465, 492686, 492189, 
    493556, 493100, 492942, 494650, 494392, 493773, 495245, 495538, 495414, 
    495265, 496164, 496844, 495685, 497742, 496815, 497240, 497564, 497648, 
    498188, 498480, 499002, 498424, 500606, 500767, 499672, 501865, 501738, 
    502019, 502109, 502187, 503527, 503710, 502230, 502594, 504580, 504899, 
    505582, 505681, 507398, 508101, 507434, 508625, 507196, 508941, 509492, 
    509603, 509368, 511874, 511132, 511327, 512427, 513780, 513950, 515356, 
    515390, 515105, 516223, 517646, 517706, 517863, 519622, 519219, 520391, 
    520710, 521970,
  519653, 518984, 517914, 516576, 518436, 516921, 515395, 515047, 514078, 
    515200, 513244, 512729, 513006, 510839, 511465, 509470, 511878, 510071, 
    509784, 509056, 508741, 507677, 507302, 505638, 506620, 506569, 506498, 
    506408, 503920, 503656, 504064, 504107, 503630, 501784, 502311, 502166, 
    502377, 501296, 500103, 500103, 499345, 500283, 500758, 499024, 499044, 
    498792, 497993, 499425, 498983, 497718, 498487, 498292, 497011, 495918, 
    497460, 496143, 496946, 495372, 494062, 495581, 494641, 493851, 493287, 
    493528, 494384, 493164, 493242, 492859, 492909, 493712, 493045, 492955, 
    493859, 492534, 491992, 491363, 492259, 493040, 492071, 491512, 491191, 
    492526, 490498, 490821, 490926, 491710, 490707, 490585, 491562, 491860, 
    490568, 490797, 491012, 490106, 490601, 490469, 490982, 490551, 490670, 
    490489, 491779, 490520, 490869, 489951, 490220, 491122, 489724, 490997, 
    490789, 490685, 490051, 491251, 491695, 490987, 491130, 490991, 490500, 
    491039, 491083, 491524, 491742, 492598, 491635, 492729, 492873, 491846, 
    491692, 492932, 493934, 492860, 492069, 493992, 493734, 494591, 493563, 
    494996, 494386, 494265, 495644, 494684, 494472, 495215, 495870, 495045, 
    496266, 496403, 495324, 496338, 497438, 496661, 497415, 498132, 498014, 
    499243, 498605, 499052, 499138, 499149, 500345, 499609, 500098, 501409, 
    502276, 501830, 502840, 501058, 503453, 503723, 503492, 504785, 502746, 
    506240, 504937, 506044, 507846, 507478, 507213, 506117, 507883, 508979, 
    508883, 509621, 509161, 510921, 510235, 511523, 512106, 512739, 512638, 
    513635, 514547, 513287, 516415, 514750, 515931, 517501, 517718, 518346, 
    518467, 519531,
  518420, 518330, 517003, 516086, 516174, 516700, 514023, 514396, 514298, 
    512904, 512533, 512645, 513165, 511382, 510387, 511465, 509002, 509043, 
    508098, 508451, 508735, 507803, 507421, 506171, 505981, 506248, 505998, 
    506145, 505401, 504031, 503007, 505150, 503816, 502093, 502250, 501670, 
    502534, 500318, 500370, 499851, 500412, 500109, 498620, 499640, 499782, 
    499210, 498517, 497997, 498208, 498489, 497007, 497068, 496689, 497018, 
    497192, 495929, 495219, 495423, 495527, 495810, 495187, 495270, 495179, 
    493914, 492937, 493931, 492726, 494209, 493477, 494204, 493373, 493311, 
    491608, 492341, 492709, 492978, 492632, 493005, 492648, 492500, 492662, 
    491939, 492184, 491427, 491151, 492376, 491275, 491670, 490944, 491976, 
    492359, 490530, 490696, 491697, 491250, 491617, 491149, 490090, 489937, 
    488994, 491165, 490538, 491604, 491581, 491730, 493100, 491736, 492401, 
    490594, 491726, 491456, 491538, 491613, 491155, 491524, 491399, 492105, 
    491674, 491814, 492292, 490693, 492643, 492598, 492725, 492578, 491422, 
    492157, 491714, 491784, 492970, 493525, 494516, 493917, 493742, 494194, 
    494799, 493532, 494439, 495152, 495430, 495576, 495649, 496156, 495763, 
    495925, 496888, 497477, 496400, 496991, 496196, 498733, 499161, 498077, 
    499361, 499873, 498764, 498678, 500163, 499228, 500278, 501823, 500897, 
    500838, 501467, 502530, 502558, 502872, 502492, 503274, 505265, 503151, 
    505198, 505506, 504804, 505976, 505962, 506532, 507590, 508082, 507871, 
    508647, 509619, 508518, 508583, 511016, 510767, 510873, 512661, 512309, 
    512946, 513725, 514248, 514286, 514784, 516049, 516514, 516467, 516414, 
    518693, 518154,
  517624, 516906, 516766, 515854, 515144, 514662, 513486, 514277, 513859, 
    512762, 512883, 511104, 511877, 509010, 511356, 510922, 509166, 509956, 
    507895, 508250, 507192, 507889, 507642, 507336, 505510, 505044, 504315, 
    504609, 504063, 504007, 504012, 503104, 501923, 504700, 502141, 500929, 
    501861, 502544, 500862, 501882, 499658, 499750, 499933, 499797, 499432, 
    498894, 498215, 497276, 496907, 496681, 497231, 498719, 497065, 495852, 
    496199, 495852, 495897, 496701, 495042, 495650, 494566, 495486, 495043, 
    495994, 496120, 493364, 494005, 494638, 493507, 494263, 494589, 494360, 
    493162, 493483, 494053, 493459, 492796, 492264, 492396, 491185, 491494, 
    491899, 492180, 492598, 492001, 492219, 493143, 492394, 490960, 492211, 
    491142, 491951, 491458, 490406, 492415, 491583, 490819, 490691, 492113, 
    491416, 491532, 491629, 491492, 491910, 493139, 491553, 490594, 492139, 
    491180, 492035, 491539, 491493, 491598, 492440, 491470, 493479, 492181, 
    492580, 491624, 491645, 492967, 492048, 492502, 492626, 491953, 492937, 
    492803, 493640, 495075, 493161, 494025, 492779, 494447, 492844, 493695, 
    494811, 495326, 495834, 494535, 496289, 494910, 495839, 496685, 496215, 
    495506, 497752, 497202, 496588, 496794, 496880, 496933, 497297, 499695, 
    499411, 499133, 498624, 499190, 500954, 500676, 500166, 500058, 499670, 
    500848, 500739, 501837, 502745, 503438, 502704, 504807, 504955, 505048, 
    505336, 504680, 504402, 504800, 505217, 505803, 506409, 506561, 508671, 
    508403, 508233, 508769, 509851, 509755, 509273, 511626, 511099, 512179, 
    512276, 512561, 513111, 514308, 514411, 514257, 516408, 516051, 517034, 
    516767, 516999,
  516813, 516577, 516026, 515971, 514725, 513987, 513752, 514004, 513461, 
    513691, 511342, 511825, 510419, 510966, 509682, 510612, 509498, 508665, 
    508438, 507140, 506900, 507490, 506035, 504977, 507348, 504925, 505209, 
    505000, 503568, 503973, 504590, 501906, 503427, 503019, 503288, 503082, 
    501565, 501600, 501716, 499825, 500202, 499931, 499832, 499233, 498743, 
    498099, 499356, 498945, 497508, 497197, 498523, 498498, 498065, 496828, 
    495119, 497104, 495884, 496715, 495041, 494569, 494889, 495757, 494648, 
    493814, 494961, 494991, 493833, 493473, 494025, 493100, 494498, 494220, 
    494112, 492164, 493695, 494153, 493315, 492451, 493042, 491718, 492344, 
    491808, 492380, 493082, 492585, 492286, 491950, 491453, 492996, 491550, 
    492819, 491776, 492769, 491553, 492137, 492393, 491637, 491100, 490629, 
    491469, 491504, 491217, 491886, 492138, 491802, 492036, 491104, 492323, 
    491076, 490652, 491675, 491567, 491785, 491841, 492153, 492369, 491933, 
    492181, 491744, 491947, 492307, 493254, 492264, 494278, 493431, 494066, 
    491778, 493017, 494792, 493943, 494486, 492850, 494542, 494231, 495531, 
    494668, 495611, 495005, 495481, 495123, 495856, 496530, 495034, 496424, 
    497969, 497479, 497479, 495957, 497408, 498326, 498665, 498135, 497369, 
    499050, 499222, 499357, 500745, 498898, 500795, 500086, 501371, 500529, 
    502518, 501717, 501297, 500800, 503302, 503116, 502634, 502340, 504159, 
    503869, 504644, 504617, 506186, 505815, 505166, 506974, 508632, 506942, 
    508664, 507912, 508477, 509542, 508549, 509699, 510590, 511157, 512300, 
    511800, 513258, 512944, 513262, 514035, 514714, 514108, 515946, 516340, 
    516776, 516919,
  516542, 515117, 514752, 515314, 514289, 512731, 514159, 513363, 511670, 
    511427, 511261, 510058, 510494, 509511, 509623, 510094, 507664, 507430, 
    508591, 507850, 507673, 506530, 505847, 506236, 504617, 504329, 505575, 
    505092, 503287, 504734, 503208, 503897, 503432, 502361, 501814, 500667, 
    500753, 502012, 500983, 501029, 499016, 500138, 501026, 499135, 499117, 
    499700, 499327, 498990, 497808, 497648, 498409, 497573, 497112, 496910, 
    498070, 495994, 497145, 495739, 496721, 494543, 496001, 494315, 495232, 
    495057, 495307, 494870, 495831, 493569, 494913, 493465, 494823, 493684, 
    493982, 493216, 492437, 493313, 494400, 493800, 492766, 493578, 493164, 
    493660, 494091, 492726, 491812, 491955, 492439, 492781, 492358, 493037, 
    491772, 490878, 491546, 491777, 491349, 491653, 492117, 492575, 491958, 
    492233, 492016, 492600, 491823, 492968, 493188, 492687, 492267, 491955, 
    492162, 492615, 493209, 492730, 492423, 493476, 493083, 493710, 492506, 
    492728, 491955, 492503, 493742, 492353, 493155, 493665, 493343, 493890, 
    493491, 494230, 493297, 495646, 493931, 493799, 496315, 494510, 493722, 
    494853, 495356, 494965, 496042, 495912, 494852, 495896, 496398, 497095, 
    497573, 495616, 496200, 497171, 497043, 499479, 499136, 499635, 498301, 
    497136, 498943, 499135, 498553, 500272, 500451, 499202, 499867, 500807, 
    501655, 503109, 502565, 501632, 502531, 503701, 503072, 503037, 503654, 
    504296, 504708, 504381, 504977, 504923, 505643, 505492, 506289, 508516, 
    506649, 507826, 507304, 508052, 509419, 510613, 509565, 510916, 510617, 
    512136, 512438, 511717, 512619, 512810, 513180, 515491, 514236, 514386, 
    515736, 515949,
  515641, 515017, 514511, 513942, 513564, 511766, 512709, 512031, 512749, 
    511208, 510260, 510052, 509145, 508653, 509877, 509808, 507433, 509307, 
    506549, 507439, 506877, 506414, 505603, 505556, 505648, 504897, 505500, 
    504444, 503718, 504138, 504272, 502068, 502283, 503295, 501001, 500367, 
    501005, 501673, 501289, 501677, 500131, 501597, 500522, 499497, 498250, 
    498574, 499007, 498893, 496468, 497145, 497544, 496598, 496867, 497095, 
    497495, 496676, 497006, 496304, 496471, 497018, 496956, 494721, 496051, 
    495919, 496679, 494762, 495032, 493660, 493780, 493590, 495035, 494372, 
    492434, 493889, 493426, 493179, 493582, 493617, 493412, 493729, 493435, 
    493419, 492756, 494514, 491802, 492897, 493779, 493028, 492121, 493679, 
    491779, 493680, 493280, 490709, 493430, 492692, 493187, 493306, 490606, 
    493880, 492529, 491895, 492722, 492403, 491451, 492955, 492367, 493935, 
    492544, 493920, 493239, 492568, 492695, 493379, 493610, 493399, 492265, 
    493061, 492932, 492678, 492376, 494593, 492473, 493405, 494770, 493394, 
    494705, 493960, 494517, 493800, 494135, 495094, 493718, 495148, 495632, 
    495944, 495586, 494555, 496372, 496773, 496064, 496194, 496461, 496536, 
    496379, 497182, 497988, 496373, 498095, 497902, 498068, 497900, 498806, 
    498646, 499950, 497965, 499281, 499721, 499686, 501004, 500834, 501342, 
    500126, 501454, 502284, 501020, 502661, 502780, 502919, 502936, 504143, 
    503823, 503774, 504911, 504705, 505575, 504774, 507060, 507725, 507053, 
    507099, 506933, 507935, 509160, 508421, 509058, 508498, 510770, 510080, 
    512382, 511554, 511788, 512115, 511073, 513396, 513334, 513841, 514463, 
    515108, 515046,
  513004, 512490, 511310, 512007, 510829, 510502, 509965, 510528, 510047, 
    508612, 509367, 508007, 509167, 508162, 507600, 508021, 505656, 506694, 
    505864, 506328, 505704, 505664, 505689, 503898, 504588, 504601, 503082, 
    503491, 503428, 503346, 503092, 502202, 501474, 502154, 502185, 500148, 
    499714, 501192, 501796, 499458, 501310, 499820, 500597, 499162, 500302, 
    498729, 499532, 497879, 497822, 499494, 498585, 498338, 497968, 497528, 
    497171, 498585, 497797, 497308, 496113, 496643, 496303, 495485, 496049, 
    497082, 495649, 496634, 495015, 494138, 497614, 495667, 494609, 494887, 
    496578, 495410, 495380, 493593, 495762, 494625, 494438, 494652, 494505, 
    493757, 494456, 493749, 494853, 493590, 494644, 494578, 493286, 493308, 
    493305, 494141, 494542, 493771, 493450, 494174, 492716, 493825, 494688, 
    493928, 492847, 494166, 494165, 492934, 492580, 493459, 494013, 493382, 
    493658, 493510, 494424, 493416, 494614, 494120, 495337, 492821, 495004, 
    493714, 495176, 495550, 494776, 494055, 495414, 494648, 495034, 495173, 
    494839, 495406, 495487, 494881, 495096, 494737, 495030, 495204, 496944, 
    495847, 496341, 497385, 496745, 495925, 496257, 497584, 496774, 497684, 
    497465, 498059, 497307, 497696, 498113, 497035, 498161, 498700, 499067, 
    500087, 499532, 499577, 499711, 498739, 500487, 500108, 498998, 501346, 
    500813, 501698, 501253, 502655, 503440, 502877, 502729, 502719, 503086, 
    504341, 503720, 503167, 505104, 504346, 503506, 503999, 504083, 504423, 
    505437, 505797, 507057, 507270, 509044, 507214, 507491, 507829, 508520, 
    508673, 508686, 510230, 511410, 510439, 510115, 510702, 512145, 511984, 
    511864, 513204,
  510698, 510145, 512008, 507904, 509812, 509608, 509600, 507994, 508327, 
    507233, 508021, 506942, 506984, 506877, 506825, 506023, 505520, 506466, 
    504532, 505172, 505403, 503586, 504208, 503638, 503858, 504147, 504005, 
    503322, 502452, 502909, 502211, 502783, 502345, 501249, 502019, 501211, 
    501429, 500640, 499714, 500521, 500235, 501165, 499149, 499070, 499449, 
    498866, 497640, 499523, 499102, 498652, 498733, 498028, 498704, 498664, 
    499013, 498357, 498550, 496855, 496197, 496984, 497492, 496896, 496998, 
    497026, 495653, 497035, 496169, 495812, 495454, 495934, 495341, 497309, 
    496320, 494991, 495491, 494646, 496157, 495124, 494749, 496008, 495200, 
    494916, 496469, 495415, 495707, 496098, 496395, 494980, 494497, 493989, 
    493691, 494122, 494192, 494416, 495727, 494663, 493901, 495012, 494233, 
    494638, 494161, 494055, 494178, 494290, 495471, 492974, 495768, 495939, 
    494165, 493908, 495274, 495394, 494879, 495734, 493845, 497092, 495165, 
    493994, 495881, 495271, 496675, 494498, 496087, 495331, 495544, 495183, 
    495560, 495960, 494923, 495003, 495928, 495864, 497583, 496366, 495433, 
    496326, 496641, 497798, 497863, 497814, 497764, 497699, 496908, 497889, 
    498363, 497846, 497039, 498394, 497936, 499126, 499156, 498899, 499062, 
    497991, 499110, 499041, 500327, 499107, 499556, 499898, 500981, 500336, 
    500554, 501663, 500560, 502369, 500754, 502745, 502418, 502383, 501491, 
    504376, 502318, 502461, 503831, 503923, 503083, 504910, 505035, 505438, 
    504368, 505473, 505026, 507104, 506934, 506586, 506352, 505892, 507420, 
    507996, 508671, 507722, 508421, 508609, 508531, 509528, 511254, 510521, 
    510212, 510678,
  509418, 509111, 508920, 508329, 508585, 506640, 508690, 507954, 506996, 
    506983, 506435, 506632, 506032, 505867, 505550, 505313, 505734, 505342, 
    505000, 504726, 503568, 502676, 504295, 502940, 504155, 504056, 502947, 
    503024, 501409, 502035, 502542, 501250, 501571, 500495, 501431, 501748, 
    500443, 501579, 500725, 500517, 500135, 500565, 499344, 498833, 498608, 
    499455, 499957, 498828, 500329, 499265, 499208, 498806, 498788, 498289, 
    497253, 498352, 496864, 496448, 498061, 497441, 497256, 497177, 498267, 
    497570, 497577, 497798, 495624, 496978, 497879, 496728, 496533, 496695, 
    496089, 496123, 495694, 495850, 495650, 495806, 496634, 495818, 495415, 
    495356, 495954, 495849, 495811, 495110, 495288, 496357, 494916, 496271, 
    493907, 495774, 495312, 495590, 495814, 495815, 494822, 495770, 496171, 
    495100, 495738, 495838, 495022, 495291, 494763, 495181, 494852, 496527, 
    494860, 494686, 495602, 495299, 495187, 495986, 494864, 496441, 495858, 
    496340, 495540, 495580, 495324, 495137, 495317, 496403, 496952, 495403, 
    496971, 496484, 497088, 496196, 495496, 497346, 497459, 495980, 496357, 
    497830, 497280, 497553, 497720, 497733, 497742, 498254, 497331, 497608, 
    497040, 497023, 499187, 500071, 498022, 498198, 498278, 499690, 498765, 
    499928, 500377, 499653, 499684, 500612, 500091, 499515, 499702, 500617, 
    501365, 501612, 500365, 501294, 500801, 501890, 501753, 501832, 502094, 
    501928, 502898, 503284, 502386, 503566, 502793, 506814, 503521, 504138, 
    504774, 503671, 505154, 505329, 506173, 504470, 505388, 505981, 506616, 
    508071, 505720, 507270, 507587, 507597, 508379, 507747, 508474, 508654, 
    509605, 509493,
  508210, 508219, 507906, 506963, 508842, 506344, 506545, 506218, 507445, 
    506519, 505615, 506103, 506144, 504339, 505183, 505566, 504009, 503413, 
    503777, 504337, 503709, 503093, 503436, 503729, 502789, 503222, 503794, 
    500847, 502503, 501020, 502926, 501090, 501475, 501909, 502479, 499971, 
    501076, 500913, 500151, 500268, 499715, 499685, 499573, 500233, 500044, 
    499561, 500150, 499391, 498616, 498014, 498978, 498298, 497884, 499001, 
    498033, 498065, 498494, 498869, 498283, 497729, 497870, 498110, 496362, 
    497109, 496676, 497346, 497796, 496934, 496405, 496828, 498032, 497744, 
    496104, 496095, 496883, 496514, 495926, 497105, 495970, 496561, 496034, 
    497191, 497521, 497112, 496437, 494751, 495718, 496581, 496732, 497023, 
    495824, 495204, 494975, 496142, 496142, 495339, 494570, 496296, 495497, 
    496612, 496253, 495014, 496659, 494734, 495310, 495169, 496372, 495893, 
    496367, 495964, 496020, 496413, 495293, 494664, 495553, 496256, 497533, 
    496769, 496461, 496128, 496024, 496380, 495810, 496525, 497168, 496326, 
    496229, 496625, 496646, 497663, 498306, 495669, 497556, 496023, 496508, 
    498634, 497684, 497475, 497940, 499022, 496991, 497697, 498407, 498716, 
    497911, 498926, 498121, 497392, 499407, 498586, 499910, 498871, 499849, 
    499713, 500009, 499588, 499251, 499076, 500500, 500066, 498250, 501154, 
    501079, 500675, 501659, 501118, 502081, 502514, 501525, 502087, 501211, 
    501861, 502780, 502972, 501710, 502321, 503367, 503140, 504519, 504029, 
    504358, 504020, 504773, 503723, 504580, 505243, 505385, 505239, 505870, 
    505376, 505791, 507028, 506422, 507469, 506479, 506921, 507979, 508128, 
    507940, 508414,
  507710, 507071, 507546, 506878, 505448, 506662, 506714, 506207, 505335, 
    505578, 505911, 505237, 504780, 504426, 504519, 504508, 503537, 503291, 
    504364, 502950, 504216, 503273, 502720, 503178, 503012, 502648, 501259, 
    503259, 502099, 501400, 501547, 500052, 502613, 502349, 500495, 500470, 
    501343, 500034, 500898, 500538, 499656, 498876, 500264, 500507, 499372, 
    499502, 499051, 499420, 500203, 498943, 499698, 498792, 497952, 498635, 
    498474, 497847, 497864, 499473, 497923, 497648, 497567, 497658, 497882, 
    497642, 498098, 498499, 496823, 498163, 499844, 497498, 496133, 496547, 
    497917, 496330, 496775, 497057, 496813, 496677, 496671, 495811, 495459, 
    496864, 495855, 495642, 496968, 495078, 496251, 496769, 496671, 497112, 
    496346, 496947, 495938, 496062, 496510, 496649, 495631, 496141, 495909, 
    496674, 496480, 496115, 496215, 495689, 496156, 496178, 496551, 497041, 
    496329, 497495, 497004, 494935, 496623, 496550, 497167, 496151, 497746, 
    496132, 496127, 496496, 497465, 495999, 497187, 495726, 496482, 496070, 
    497497, 497728, 496429, 496699, 498764, 497253, 498286, 498141, 497520, 
    498300, 496197, 499719, 497690, 497733, 497962, 497867, 498034, 498654, 
    497985, 499046, 497951, 498387, 499305, 499407, 498304, 498751, 499402, 
    500552, 499618, 499176, 499227, 500530, 500168, 500356, 501399, 500110, 
    500558, 500211, 499952, 500263, 501452, 501503, 501938, 502350, 501848, 
    501964, 501523, 502641, 503130, 503685, 502658, 503722, 503210, 503008, 
    503127, 503996, 503862, 503334, 504720, 504604, 504229, 503903, 504902, 
    505978, 506473, 504589, 505228, 507223, 507285, 505703, 507015, 506896, 
    507541, 507463 ;

 true_corr_mean =
  -0.913533120455018, -0.843096077181069, -0.800226984195975, 
    -0.767710977561849, -0.739163880823788, -0.714912006930591, 
    -0.692859301735076, -0.673755746908881, -0.655146526898708, 
    -0.637460669698469, -0.621822923639206, -0.606870860621593, 
    -0.593337304219088, -0.578906658858212, -0.566258950123296, 
    -0.55294861335054, -0.541757290107362, -0.53032989212684, 
    -0.518622143662702, -0.508466064841381, -0.498114645096303, 
    -0.487969402052082, -0.47737684064841, -0.468950958289695, 
    -0.458882789655332, -0.451167190767064, -0.441038069278487, 
    -0.43255720275585, -0.423882508703808, -0.415052294016757, 
    -0.407702237498575, -0.399187289773097, -0.392130551586596, 
    -0.383759594895485, -0.375608595432397, -0.367505882086914, 
    -0.361192414235949, -0.353950377181781, -0.346405409675412, 
    -0.339723582127893, -0.331997708054946, -0.32522857335909, 
    -0.319696018908193, -0.311842525248471, -0.304967380774823, 
    -0.299066476702274, -0.292377978079589, -0.286521241429441, 
    -0.279101383143617, -0.272355868404347, -0.267077995212802, 
    -0.261447859080913, -0.255907983062271, -0.248683184442962, 
    -0.243551373667494, -0.2380481328704, -0.228862046424933, 
    -0.225127998822826, -0.218920221019191, -0.212512302038089, 
    -0.208122399360132, -0.202299017607585, -0.195343042085182, 
    -0.189930866796858, -0.18469459107826, -0.178651112003975, 
    -0.173626138705467, -0.167721738798722, -0.162834933255606, 
    -0.158240788782378, -0.152405303459335, -0.147612320849773, 
    -0.141747100987252, -0.135535934588959, -0.131531615377297, 
    -0.125710286482574, -0.119915802577165, -0.11564031597842, 
    -0.10876880798984, -0.103610792828107, -0.100898816548386, 
    -0.0941219268312776, -0.0874841969216722, -0.0846569819017256, 
    -0.079501645222881, -0.0750146319605614, -0.0694498445282589, 
    -0.0640419123405948, -0.0575088472461902, -0.0545005480195816, 
    -0.0494158333203924, -0.0434982683300794, -0.0384582481859887, 
    -0.0318290699834649, -0.0281297645485643, -0.0242687193436646, 
    -0.016298758934404, -0.013466593065544, -0.00874803854695804, 
    -0.00215816270308191, 0.0024777939480077, 0.00794326052976886, 
    0.0129365317540174, 0.0181999161333004, 0.0227064628639894, 
    0.0265433711439349, 0.0346905347153112, 0.0383773784125857, 
    0.0431944891290731, 0.048059033291719, 0.0542885670949517, 
    0.0581905084525709, 0.062622139008371, 0.0675806610163599, 
    0.0744675812720974, 0.078513143916142, 0.0837067634940263, 
    0.0888225228694915, 0.0931714577186573, 0.0979357392396977, 
    0.104399640131671, 0.109606906811346, 0.114918351812807, 
    0.119820200688956, 0.126023848005462, 0.131155356695721, 
    0.13710426328592, 0.141532151067017, 0.147780195820549, 
    0.152683586538147, 0.157788487825085, 0.163581083153665, 
    0.168492124734939, 0.17384232154136, 0.179538148614132, 
    0.184543090312679, 0.19090522358259, 0.196766192729411, 
    0.201557093898235, 0.207464920834022, 0.212870456569528, 
    0.219333952989217, 0.225918391089571, 0.23131080775466, 
    0.236609963413576, 0.242778250990662, 0.247337229677383, 
    0.255718820222734, 0.260538558251908, 0.267997703075238, 
    0.272992893785035, 0.279537609460446, 0.286999666495872, 
    0.29242455388284, 0.298689006350613, 0.306234501524128, 
    0.311895268517345, 0.318325187903983, 0.326667198208322, 
    0.332510324578859, 0.339944040613909, 0.347160312026797, 
    0.353205933993982, 0.361443872201707, 0.369383746359823, 
    0.37588858534597, 0.383621270532717, 0.391321481911873, 0.3991300857127, 
    0.407761970929946, 0.415623417601002, 0.42406022522342, 0.43248379880381, 
    0.440876997221026, 0.449273115101852, 0.459103656515662, 
    0.468378132035309, 0.478397515696717, 0.488265131737895, 
    0.497450590725965, 0.508538901271236, 0.519753784159855, 
    0.530067066433916, 0.541930309609859, 0.553423689950655, 
    0.566355269007855, 0.578987231053219, 0.59279343707387, 
    0.606911672007746, 0.622087708299949, 0.637979154964509, 
    0.654798766758482, 0.673487877413716, 0.693458661604457, 
    0.71482250718545, 0.739431177297288, 0.767064484303568, 
    0.800171619829262, 0.842987459050229, 0.913696895651076,
  -0.956038425985297, -0.901615056835609, -0.862963480780387, 
    -0.831711705433517, -0.804662886398226, -0.780325896532865, 
    -0.758375630798595, -0.738244138629596, -0.719304887091071, 
    -0.701323117246212, -0.684713247024421, -0.669053866954304, 
    -0.65389934028949, -0.639754122870923, -0.625473519948943, 
    -0.613185337836095, -0.599971503611794, -0.587578179928821, 
    -0.575696243250596, -0.563640434765195, -0.553134684146517, 
    -0.541236872065053, -0.531253697821117, -0.520724358469864, 
    -0.510977021937931, -0.500195304885074, -0.491081370047555, 
    -0.481112271813653, -0.472250827874463, -0.462398637079355, 
    -0.454109915975208, -0.443714396168826, -0.4366648093625, 
    -0.42765317135194, -0.419692966308148, -0.410526126675846, 
    -0.402974711192484, -0.395114961795676, -0.386603774338274, 
    -0.378045357327034, -0.371598941023155, -0.363830063893828, 
    -0.356310415424631, -0.348644314473082, -0.341325688592737, 
    -0.333877783061954, -0.325748438804933, -0.319055858151923, 
    -0.313243675822805, -0.305936864422135, -0.298968560444842, 
    -0.290877426533706, -0.285127006062649, -0.278306021246733, 
    -0.271565538883182, -0.26500301441576, -0.259943858897128, 
    -0.252096381299203, -0.24501699366837, -0.239401024040963, 
    -0.232329945388933, -0.226331279314149, -0.219784269910918, 
    -0.213005146999549, -0.20841951358632, -0.200527658747535, 
    -0.196165600355661, -0.188888695419647, -0.183070690595352, 
    -0.176652315588165, -0.170206501627788, -0.164216776394672, 
    -0.157767988385842, -0.152411168395638, -0.147060119784336, 
    -0.13992685911809, -0.134995845644391, -0.128287241285253, 
    -0.121624467037999, -0.117252389519305, -0.111836908212092, 
    -0.105115034839281, -0.0991766212840372, -0.09399911827609, 
    -0.0874461332355129, -0.0826179801601686, -0.0765341326768938, 
    -0.0704363906387308, -0.0654254789508003, -0.0593055473342918, 
    -0.0537250368397449, -0.0491729294548997, -0.0429988930681223, 
    -0.0373963280916576, -0.0316109352064619, -0.0257189258627343, 
    -0.0200610498908396, -0.0132188160680548, -0.00871812568540898, 
    -0.00144243643479377, 0.00288930719383454, 0.00864528799700643, 
    0.014533412975445, 0.0188837767367683, 0.0247388382800539, 
    0.0311789917552926, 0.0367489673205575, 0.042021086530463, 
    0.0471452473925742, 0.0543174757505479, 0.0585048545416291, 
    0.0659106813075236, 0.0704249674647338, 0.076338218551, 
    0.0821531944634836, 0.0884137957582706, 0.0946813230528476, 
    0.0999045798004723, 0.105064400719685, 0.111788667576962, 
    0.116199680957571, 0.123601330956418, 0.128227610219933, 
    0.134633884535772, 0.141054740354888, 0.146468478603791, 
    0.152065237948573, 0.158396573364946, 0.163896063456493, 0.169291142155, 
    0.176041487781908, 0.182481499971563, 0.189581806509559, 
    0.194685123810687, 0.200539071446769, 0.207390317242811, 
    0.21244615470321, 0.219568126617839, 0.225773762997592, 
    0.233499534791221, 0.238439770724859, 0.244668866695554, 
    0.252370182770676, 0.257280949846165, 0.265364791899061, 
    0.272065010489944, 0.27927808249744, 0.284426151456754, 
    0.290705842484824, 0.298926968160663, 0.305771518239923, 
    0.313055347240879, 0.31885345462933, 0.327204948942225, 
    0.333137909768229, 0.34250837495142, 0.349359213219381, 
    0.355569563767558, 0.363305887661416, 0.371244467007247, 
    0.378318769984081, 0.387017180412614, 0.395063570131904, 
    0.403626260314869, 0.411245887609638, 0.418733100011975, 
    0.427244815531757, 0.436837687272343, 0.444548165661842, 
    0.453827498410005, 0.461610935632946, 0.471593110768602, 
    0.481490779894616, 0.490412125988672, 0.500610592326314, 
    0.510536930911671, 0.520420574152443, 0.531138953618905, 
    0.54147801240838, 0.552908970937094, 0.563770698910377, 0.57553254396548, 
    0.587325233298829, 0.600524137116967, 0.613098350813151, 
    0.62600213030237, 0.639523027256492, 0.653892700707193, 
    0.668838386665514, 0.684378489743242, 0.701413547383001, 
    0.719148683156758, 0.737641318200023, 0.757971079163645, 
    0.780498345123092, 0.804476521374744, 0.831674454049134, 
    0.863084669970295, 0.90146514683704, 0.956025767805036,
  -0.972875369298955, -0.930984882824377, -0.898015875861099, 
    -0.869960320184338, -0.844514165002959, -0.821295579054382, 
    -0.800126654321435, -0.780609675575176, -0.761827986851584, 
    -0.744238484637487, -0.727479838163366, -0.712204072048578, 
    -0.696134157641036, -0.681936608538982, -0.667365564924766, 
    -0.653833045186656, -0.640954888995999, -0.62820552449428, 
    -0.615815626602188, -0.603692741869382, -0.592351398060364, 
    -0.581045153537965, -0.569501312069648, -0.559186611048769, 
    -0.547540548564049, -0.537699665172841, -0.527283557680221, 
    -0.516940552008266, -0.507479064558806, -0.497534695272446, 
    -0.48837750438672, -0.478876798875518, -0.469540595553353, 
    -0.460698878609607, -0.451352590075022, -0.44330329055583, 
    -0.433733177333566, -0.425615162566829, -0.416548937096451, 
    -0.409049829931424, -0.400794027371933, -0.392530475194818, 
    -0.384228868152336, -0.376499486096732, -0.368553751914797, 
    -0.360625695905508, -0.352791364648199, -0.345436754393399, 
    -0.337599336085228, -0.329468686273616, -0.322533774090197, 
    -0.316135742076311, -0.308356618606139, -0.301361337527223, 
    -0.293535003428822, -0.286649575919331, -0.279975014347917, 
    -0.272955735934299, -0.265532770995235, -0.258333041067697, 
    -0.252381312710053, -0.244446193003793, -0.237746110037562, 
    -0.23104233163576, -0.224532848958091, -0.217797016078774, 
    -0.211149551064787, -0.205035949068212, -0.198110180042228, 
    -0.191374154587567, -0.185221121404524, -0.178425532101044, 
    -0.171476081357623, -0.165131743936249, -0.15900607062449, 
    -0.152887059147792, -0.145407282043559, -0.139670370136895, 
    -0.13423592668563, -0.127202449020439, -0.121214777103625, 
    -0.114720069045819, -0.109190485575089, -0.101773469391062, 
    -0.0959034569881461, -0.0893244885800029, -0.0834707581894443, 
    -0.077435465451026, -0.0703412723325396, -0.0636565130152701, 
    -0.0588933102641885, -0.0523314836151334, -0.0460448738955201, 
    -0.0402312876978722, -0.0333171616490866, -0.0276235341473133, 
    -0.0208872302578275, -0.0150784762917254, -0.00992772416732606, 
    -0.00359665668854002, 0.00247918433031465, 0.00935185813515229, 
    0.0154380480762303, 0.0220336412741346, 0.0283836479409827, 
    0.0339691216246406, 0.0409345662325717, 0.0464993605264914, 
    0.0522829509177048, 0.0580534773575439, 0.0633256627096466, 
    0.0700291595786175, 0.0766431698357161, 0.0831193551343279, 
    0.0896799399243041, 0.0955988638757298, 0.101526681237365, 
    0.107308307630783, 0.114989621657791, 0.12095383550047, 
    0.127653691446987, 0.133966973120923, 0.140742985109436, 
    0.146074018346735, 0.152806418607374, 0.158729091378344, 
    0.165333641500746, 0.171885608443229, 0.178709736005664, 
    0.184727596059429, 0.191263396823815, 0.198174031031661, 
    0.205291855784572, 0.210882648880731, 0.216769220353002, 
    0.22415418503585, 0.230754003314043, 0.238196096633847, 
    0.244698763226338, 0.25225138246519, 0.258140140203732, 0.26603569728263, 
    0.271907453437402, 0.279963211816086, 0.286327340471215, 
    0.294390724385152, 0.301546683068406, 0.307841416854418, 
    0.315338556891707, 0.323629215372032, 0.330047043117534, 
    0.33799317331613, 0.346252470556072, 0.352669072974311, 
    0.361015571157255, 0.36866434601209, 0.377329199910292, 
    0.384080016117382, 0.392918408683119, 0.400543965324101, 
    0.408577646504704, 0.417018999362962, 0.425627512514781, 
    0.434455766595617, 0.44325250093764, 0.451461761432834, 
    0.460446578102352, 0.469489709330455, 0.479101270958581, 
    0.488631996927561, 0.497708776997426, 0.508372636747394, 
    0.516839297160366, 0.52616971977291, 0.537979452832255, 0.54866145610057, 
    0.558751022578098, 0.569672280228304, 0.580211293822789, 
    0.592281681345568, 0.604066744833477, 0.616349470209121, 
    0.628588112174866, 0.641270385707766, 0.65446228392665, 
    0.667527513293671, 0.681410907034482, 0.696762777399875, 
    0.712277904341595, 0.727446162874223, 0.744179850019586, 
    0.761423772496922, 0.780427604149307, 0.800389573849495, 
    0.821796093126291, 0.844316627628444, 0.86951313638381, 
    0.898075034217432, 0.931078977569854, 0.97297193579129,
  -0.980547568927585, -0.946949338860792, -0.918316563615793, 
    -0.892962472916511, -0.86971258489614, -0.84817680995109, 
    -0.828271737065628, -0.809304826886346, -0.791210671146473, 
    -0.774216736853529, -0.75806383641652, -0.742275202176755, 
    -0.727121358561797, -0.712541366127294, -0.698016520115308, 
    -0.684215056965067, -0.67184874522448, -0.658878654161492, 
    -0.645341907976448, -0.633516460711501, -0.62182758325613, 
    -0.610055023759638, -0.598643736624857, -0.587156865501295, 
    -0.576691279218972, -0.566177376091733, -0.555033384254019, 
    -0.544934151904346, -0.53448133176252, -0.525125644965088, 
    -0.515582663060571, -0.504790497302088, -0.495708818545893, 
    -0.486305222661558, -0.477226888634751, -0.467922600500366, 
    -0.458877304341969, -0.450074649796925, -0.44111529181221, 
    -0.432242717927323, -0.423719524199128, -0.414830799942035, 
    -0.406750522674261, -0.398178529742434, -0.389454427274589, 
    -0.381403463338732, -0.3732071774151, -0.365377728946215, 
    -0.358110407664129, -0.349783409894909, -0.341938474759671, 
    -0.33420633706563, -0.325877624202865, -0.31849360865377, 
    -0.310928691709204, -0.30354299573225, -0.29683928465154, 
    -0.289082887592968, -0.282142267072934, -0.274052909234266, 
    -0.267012540135185, -0.260321170936075, -0.251822602879275, 
    -0.244385454815305, -0.238172138861709, -0.230936955319349, 
    -0.223982447878692, -0.217230160473836, -0.210080688162591, 
    -0.203802881443246, -0.195783108732994, -0.189184708189739, 
    -0.182084323590431, -0.175750755879845, -0.168853192313404, 
    -0.161149008644414, -0.155282524326333, -0.148064717319094, 
    -0.141483147177789, -0.134733788288224, -0.128098440044203, 
    -0.122330466935284, -0.114228035727765, -0.108311155893241, 
    -0.101490197268763, -0.0946054859063776, -0.0877011387979962, 
    -0.0818453610980086, -0.0756643942319571, -0.0693385863665402, 
    -0.0616712410963574, -0.0555585483127386, -0.0489143691954302, 
    -0.0427859175034063, -0.0363144419307704, -0.0293045250126367, 
    -0.0234930868084438, -0.0162204075033162, -0.00982064846535498, 
    -0.00164745864786303, 0.00365614357090181, 0.00901236127962176, 
    0.0168890000046217, 0.0233498164213948, 0.0293269028126065, 
    0.0352833124497863, 0.0419136421754571, 0.0493271330564699, 
    0.0552208834827026, 0.0625814399042102, 0.0681307172624673, 
    0.0762021666459836, 0.0811729755110416, 0.0874193679723774, 
    0.0946135440147537, 0.101417822517973, 0.10820401237819, 
    0.114706036622099, 0.1219658095514, 0.128926382277669, 0.13509283779723, 
    0.142152833766473, 0.147874565105957, 0.15501521834628, 
    0.162186325251465, 0.168895405056041, 0.175527509896274, 
    0.182109446963392, 0.189429871227162, 0.195185744315935, 
    0.203116688889144, 0.210458000437899, 0.216816623055145, 
    0.224395969896082, 0.231748716074567, 0.238869882546687, 
    0.245769133080039, 0.252885039079663, 0.259977473440853, 
    0.266224107578193, 0.275263448198045, 0.281635770457428, 
    0.288678574083295, 0.296316763076775, 0.303915375849062, 
    0.311802815937496, 0.318126973089951, 0.326626151460566, 
    0.33456423850661, 0.341813058684399, 0.349115611720956, 
    0.357157031805008, 0.366603253041644, 0.374082173234436, 
    0.382685909806433, 0.389570671261948, 0.398219816046704, 
    0.406482178441086, 0.414910095752987, 0.423694251148701, 
    0.431934154317811, 0.440267301989466, 0.448367500405528, 
    0.458032803198124, 0.467273399497717, 0.476927394775193, 
    0.486407879703488, 0.496256047296122, 0.50518644656889, 0.51435392044264, 
    0.524933007602804, 0.534463617173758, 0.544602321521787, 
    0.555610687671846, 0.566107890016146, 0.576500180745224, 
    0.587410106015775, 0.599188086051818, 0.610361023017967, 
    0.621718781304712, 0.633640910813915, 0.64588373584219, 
    0.658961813137571, 0.671265392486252, 0.684647792882058, 
    0.697772885679536, 0.712603900773483, 0.72704749455847, 
    0.742188406963199, 0.757915212464939, 0.774289860036911, 
    0.79095995270815, 0.809148737094944, 0.828076436269897, 
    0.848367983463755, 0.869766721272766, 0.892997195788188, 
    0.918551434160441, 0.946989698799598, 0.980530690575195,
  -0.984494993128412, -0.956195077730587, -0.931077770394881, 
    -0.907899237372468, -0.886671487236368, -0.866630989932216, 
    -0.847389720499124, -0.829530778471359, -0.811883130921974, 
    -0.795233214442751, -0.779911333317084, -0.763998756680041, 
    -0.749583116896462, -0.735345246845249, -0.720537449394786, 
    -0.707305514139788, -0.694072161924291, -0.681343793014214, 
    -0.668744614092484, -0.65602236470126, -0.644457405223776, 
    -0.63234579457594, -0.620782184760923, -0.609720560887245, 
    -0.598753555282766, -0.587257621520618, -0.577051045370288, 
    -0.566138021111653, -0.555829250664086, -0.545374388825747, 
    -0.535550074599807, -0.52564056418521, -0.516040160190168, 
    -0.506138030845252, -0.497409938441386, -0.487596188060336, 
    -0.478429987095805, -0.469032431782506, -0.459945069196563, 
    -0.451053900058842, -0.441418497906201, -0.432994968437884, 
    -0.424536654191166, -0.416136193233317, -0.407139204102985, 
    -0.398914229618467, -0.389929024364424, -0.38172929095123, 
    -0.374023868364393, -0.365879943858037, -0.358241322209491, 
    -0.349494680096483, -0.341578159277242, -0.33343302198751, 
    -0.325666718578742, -0.317547367146417, -0.310787543035763, 
    -0.302695665303443, -0.294824385054521, -0.286927607420291, 
    -0.2790348015195, -0.27198503560092, -0.264344984066423, 
    -0.256077857948623, -0.249365718984139, -0.243029652378641, 
    -0.234556102214254, -0.227633376701395, -0.220155303445081, 
    -0.212720022273562, -0.205283779036916, -0.19801645799666, 
    -0.190883482063435, -0.183705516561917, -0.177151221977298, 
    -0.169363583359965, -0.162993703191229, -0.15537105291834, 
    -0.148209735751801, -0.141210373746915, -0.1342154026653, 
    -0.127968549646957, -0.120814835852641, -0.113677962747628, 
    -0.106484808115685, -0.0993557390973663, -0.0928693363892071, 
    -0.0854086486496493, -0.0791476901687242, -0.0716693868588062, 
    -0.0650237885702483, -0.0576199284244059, -0.0516577207046709, 
    -0.0451387794998479, -0.0374949894345329, -0.0307827981237776, 
    -0.0233799500968477, -0.0166734105763029, -0.0103290484400021, 
    -0.00314301189661183, 0.00361942565173752, 0.00938361238734802, 
    0.0173804143174495, 0.0234536123134993, 0.0309487641114619, 
    0.0375544024953129, 0.043948076507307, 0.0516509999013275, 
    0.0583423956905546, 0.0645184413832831, 0.0721699128777665, 
    0.0780506314513992, 0.0851572627579615, 0.0925474052835605, 
    0.099381702112034, 0.106415863065029, 0.113008642313846, 
    0.120416413161921, 0.127849305642001, 0.134723192606174, 
    0.142169074976001, 0.149389476664122, 0.156120247449481, 
    0.162333412943466, 0.170006766617108, 0.176732886128605, 
    0.183736853372242, 0.191309088550767, 0.197860339507547, 
    0.205229017831955, 0.212975826629851, 0.22016666895064, 
    0.226465691186359, 0.234179758687235, 0.241782281157918, 
    0.249300260038909, 0.256604912813577, 0.263509818838243, 
    0.27108305792902, 0.279422256244391, 0.287297224550856, 
    0.294507947333415, 0.302082520551716, 0.309224610828468, 
    0.31794879380652, 0.325474750639216, 0.333909384456815, 
    0.341167686459049, 0.348922020399585, 0.357425955418091, 
    0.36613076789581, 0.374208965623459, 0.381821848218267, 
    0.390565154365327, 0.39838187463748, 0.406974006340433, 
    0.415295105959503, 0.424481846942826, 0.432803156514095, 
    0.442405519595134, 0.450564084709045, 0.459136846333499, 
    0.468956912178639, 0.478310443514695, 0.487104806783928, 
    0.496805574619166, 0.506701837003951, 0.516021726232749, 
    0.525790579860279, 0.535612570432919, 0.545868494689695, 
    0.555971467925797, 0.566279107578859, 0.576560005569062, 
    0.58818579798577, 0.598546109050978, 0.610142138390241, 
    0.620885669611751, 0.632092117553836, 0.644019074328811, 
    0.656474875289122, 0.668588836177204, 0.681444953091481, 
    0.693924081843903, 0.707048643509093, 0.720884568211144, 
    0.734367324609556, 0.749209103789365, 0.764356522278871, 
    0.779664412614795, 0.795684984936318, 0.812184806961258, 
    0.829642659196338, 0.847591750628366, 0.86647326887211, 
    0.886649301609884, 0.908009161413891, 0.931139038874558, 
    0.956277643283081, 0.984563616046187,
  -0.986857326635862, -0.962141005669741, -0.939581226660411, 
    -0.918410891193877, -0.898575525359478, -0.879387052798839, 
    -0.861243600609534, -0.844198772208825, -0.827364986084213, 
    -0.811382284135802, -0.795929208971464, -0.780549859705593, 
    -0.766581134803068, -0.752152345888988, -0.738325511078811, 
    -0.725051267985978, -0.711910509212435, -0.699247129829712, 
    -0.686315582345957, -0.67395009885898, -0.662304673070733, 
    -0.650309223805045, -0.638551871000951, -0.627521305965226, 
    -0.616270132535126, -0.604984778355121, -0.594263405487677, 
    -0.583406209944731, -0.573888356962773, -0.562720449778519, 
    -0.552465713832672, -0.542195812251416, -0.532400536911511, 
    -0.522740988147527, -0.51255178782921, -0.503896429218117, 
    -0.494331645614017, -0.484400231735486, -0.474955677856409, 
    -0.465815478804461, -0.457228978976963, -0.447433614748483, 
    -0.439268778428888, -0.429682296009942, -0.421188978175196, 
    -0.412235884021309, -0.404186131428931, -0.395957735513786, 
    -0.386842712498312, -0.377687775256627, -0.369978923389967, 
    -0.361928290098778, -0.353303704730866, -0.345322453974168, 
    -0.337326184101501, -0.328865117222244, -0.320328075682995, 
    -0.313447993610989, -0.30470107220784, -0.297161111901012, 
    -0.289412753688399, -0.281391919579108, -0.273512867572261, 
    -0.265965863166602, -0.258856419839642, -0.251279558691762, 
    -0.242612511873915, -0.235748668412224, -0.228481633368406, 
    -0.221139415925897, -0.213696210923573, -0.205845404661586, 
    -0.198229345288882, -0.191503735957337, -0.183199038722053, 
    -0.175455390574534, -0.168197793676148, -0.16124953516414, 
    -0.154020843353511, -0.146658860927705, -0.140631395296553, 
    -0.132215558316584, -0.124472386539765, -0.118354897261092, 
    -0.10994112651029, -0.10239737202196, -0.0963855644250133, 
    -0.0890791493502671, -0.0822624646524971, -0.0738828073710105, 
    -0.0679928994098669, -0.0605735839945088, -0.0529394111139361, 
    -0.0460435654724498, -0.03960727329712, -0.031749664423445, 
    -0.0242436324801497, -0.0184308520505087, -0.010961144567005, 
    -0.00315221905019085, 0.00328177600356125, 0.0108630734105034, 
    0.0169870214874373, 0.025942295069716, 0.0315417980850972, 
    0.0393270724026448, 0.0455427441013728, 0.0534183233801293, 
    0.0607041843771286, 0.0674038022060333, 0.0747477329108538, 
    0.082218674238953, 0.0890491817601664, 0.0960903102143815, 
    0.103506948577574, 0.111628718577097, 0.118057308954755, 
    0.12544986735027, 0.13215288308591, 0.138953327793292, 0.146040286664206, 
    0.153986287409542, 0.160855890378869, 0.168315884636417, 
    0.176027304623495, 0.183630490372824, 0.190690058761713, 
    0.197432344036813, 0.206534074901825, 0.212690474782395, 
    0.220189442834265, 0.2280925921239, 0.235380334871861, 0.242923022854693, 
    0.251265211726655, 0.258568785791152, 0.265437219643981, 
    0.273231598237717, 0.28116563857234, 0.289773823488214, 
    0.298065290755044, 0.304792252358972, 0.312992229957303, 
    0.321569934269232, 0.329528952632318, 0.337486676359236, 
    0.345814087907996, 0.352937917309763, 0.361722786316493, 
    0.370631422596066, 0.378660345776107, 0.38699878269908, 0.39534422210522, 
    0.404346996676701, 0.412568477450909, 0.421394664435675, 
    0.430297878348913, 0.439127080934641, 0.447888087383286, 
    0.456436120173356, 0.465972628765872, 0.475293884577554, 
    0.483957227247036, 0.493784926475866, 0.503624562730617, 
    0.51244455723746, 0.522642938280696, 0.532350989591323, 
    0.542965322090088, 0.552225407852307, 0.562657710183261, 
    0.573236368161126, 0.584111331701501, 0.594737386672796, 
    0.605446485673233, 0.616010787613822, 0.627426117491339, 
    0.638968835968824, 0.650314695612906, 0.661942364378286, 
    0.674171797405325, 0.686613877052512, 0.699071358408498, 
    0.711677732258455, 0.72477465576958, 0.738093489615596, 
    0.752402596566972, 0.766361022294253, 0.780900175262973, 
    0.796130602706755, 0.811278006565135, 0.827696513933271, 
    0.844051284375713, 0.861160210321359, 0.879460706144681, 
    0.898387237875075, 0.918377256854842, 0.93939985929834, 0.96220524399198, 
    0.98687032985911,
  -0.989401127980446, -0.969044019577586, -0.949605691726086, 
    -0.931126689966527, -0.913311413251511, -0.896212267402858, 
    -0.879607543452206, -0.863916545453238, -0.84809818716436, 
    -0.83334245616693, -0.818107932791684, -0.804236232739155, 
    -0.790171574140868, -0.776490487125678, -0.763134102199047, 
    -0.749700753093848, -0.737042776901389, -0.724852006279291, 
    -0.712088748223117, -0.699765939293282, -0.688036310628007, 
    -0.676188168202237, -0.664551234122453, -0.653067180663329, 
    -0.642202894924528, -0.630926014041822, -0.620098556773465, 
    -0.609398460393422, -0.599056271220158, -0.588050233161207, 
    -0.577622446330843, -0.567424603819874, -0.557231683100689, 
    -0.546751113332801, -0.537269972966787, -0.527677589177586, 
    -0.51750563131236, -0.508428206752034, -0.498206480465584, 
    -0.489393622720704, -0.47949516586498, -0.47017211250578, 
    -0.461260969600304, -0.452237483988678, -0.44190461456564, 
    -0.434054434674783, -0.425226173026546, -0.415383871458067, 
    -0.406538027740756, -0.398846788432451, -0.389957608597726, 
    -0.381608589521657, -0.372182355797326, -0.363548885126456, 
    -0.35536649532955, -0.347297263043945, -0.339094761695222, 
    -0.329367671826832, -0.322026173384654, -0.313435523642995, 
    -0.305104496351912, -0.296996896056779, -0.28853400047705, 
    -0.281122479345159, -0.27330479324812, -0.26485925585192, 
    -0.256949814230808, -0.249197579366621, -0.240707396232055, 
    -0.231557033947573, -0.224997185553054, -0.216688467218222, 
    -0.209877716779516, -0.201803552234513, -0.193468529336203, 
    -0.185852087113032, -0.177945076858827, -0.170641479597599, 
    -0.162937914688617, -0.155279492938055, -0.147593360750977, 
    -0.139525295739053, -0.132102380472421, -0.124749982609462, 
    -0.116598720427398, -0.109319660879631, -0.10130961392967, 
    -0.0939840606523851, -0.0867506938554077, -0.0789371186770154, 
    -0.0726286230177281, -0.0643289748512315, -0.056927493955052, 
    -0.0492010276055979, -0.0413022647272922, -0.0337528843375244, 
    -0.0265002156939202, -0.0191294068772795, -0.0108267871425349, 
    -0.00332767773585459, 0.00390612728111918, 0.0110524408994918, 
    0.0189320930442489, 0.0264762021493374, 0.0343857584065964, 
    0.0412219254719641, 0.048088667878459, 0.0554507821210379, 
    0.0646324572147259, 0.0713787871921019, 0.0787075666453849, 
    0.0858891295769969, 0.093957109200888, 0.101811420798157, 
    0.109412274831325, 0.116639517044734, 0.123719383947861, 
    0.13132563178883, 0.139887427985919, 0.147424824052751, 
    0.155146903044258, 0.16268742072576, 0.170004314176357, 
    0.178533956820712, 0.186097906156757, 0.193954906996964, 
    0.20118002537305, 0.209950193178366, 0.216863810199797, 
    0.225066528118287, 0.233622390238902, 0.241145792998055, 
    0.248511697292411, 0.256613016854393, 0.264587885974751, 
    0.273206779365153, 0.281156714590521, 0.288742762437048, 
    0.297255174177897, 0.304792737969482, 0.31360114267543, 
    0.321515065397382, 0.330097911261818, 0.339001099242421, 
    0.346793195046552, 0.355054086584072, 0.364476530974795, 
    0.372279827109303, 0.380518012877339, 0.389569484032627, 
    0.39838572210612, 0.406859338367354, 0.41561232362833, 0.424684359719855, 
    0.433583241581145, 0.442900986038491, 0.451954494803275, 
    0.461052325531328, 0.470839483608596, 0.479189232499487, 
    0.489216579499544, 0.498653671311574, 0.508218099383886, 
    0.517582403745853, 0.52748316472015, 0.53731062255198, 0.547296767100716, 
    0.557538962074006, 0.567611662644354, 0.576840309907099, 
    0.588082668856896, 0.598134939123994, 0.609424881493853, 
    0.619951571604756, 0.630712704449258, 0.642317007162806, 
    0.653062243243112, 0.664605304191329, 0.676279298784009, 
    0.687933647194384, 0.700006139803007, 0.712049699482691, 
    0.724619361042972, 0.737139043706698, 0.749960771439277, 
    0.762937622035384, 0.776741672285235, 0.78996758686919, 
    0.804117508558262, 0.818288762024091, 0.83297028302431, 
    0.848322233710575, 0.863811347108292, 0.879808358374899, 
    0.896188935994858, 0.913400726692105, 0.931137163537089, 
    0.949607399679071, 0.968994793425654, 0.989394069554968,
  -0.990763316557802, -0.972731032605906, -0.955401928632989, 
    -0.938528590451031, -0.9222429876541, -0.90631833795049, 
    -0.891012588358373, -0.875800023656618, -0.861421703284748, 
    -0.847174632971394, -0.832670403667812, -0.819235380261287, 
    -0.805627602099647, -0.792251175447565, -0.77961899756148, 
    -0.766830604406776, -0.753977779978291, -0.741866764464742, 
    -0.729665809746013, -0.717620212867992, -0.705642081467423, 
    -0.693796162231833, -0.682376035700422, -0.67142932843777, 
    -0.659880385581727, -0.648710739499656, -0.63802299873146, 
    -0.627181283978405, -0.616461236922691, -0.60584172264411, 
    -0.595631442510995, -0.584565244722718, -0.574655123248925, 
    -0.56457276098926, -0.554764566260526, -0.544471030400091, 
    -0.534591113879333, -0.52497239399116, -0.515153798528913, 
    -0.505239607208552, -0.495737785147433, -0.486260165493727, 
    -0.476870008424915, -0.467554473271785, -0.458787226827319, 
    -0.449173811219696, -0.43987653137266, -0.430707050956025, 
    -0.422373263749701, -0.412581261697151, -0.403353652870853, 
    -0.395000008817188, -0.386026573556094, -0.377227460137739, 
    -0.369303880611023, -0.36020934382086, -0.351325408411371, 
    -0.342677833412542, -0.334167731346424, -0.325384440893668, 
    -0.31721508720639, -0.308618577856599, -0.300221261405323, 
    -0.291757604451049, -0.283269500874337, -0.275284175841429, 
    -0.267084200928611, -0.258394190672589, -0.250828357181376, 
    -0.242293163036132, -0.233874944935814, -0.225995536757197, 
    -0.217850868475619, -0.209886017579912, -0.20172458929414, 
    -0.194044188036502, -0.185199738462965, -0.177513565674135, 
    -0.169630892677158, -0.161508930882411, -0.154156146373256, 
    -0.145277654020026, -0.137889400958099, -0.129950423866533, 
    -0.121626779706364, -0.113628568594319, -0.10546829598411, 
    -0.0975857124985218, -0.0897172988895923, -0.0817984337361469, 
    -0.0744697543588626, -0.066682715344894, -0.0584713577472887, 
    -0.0512113594473242, -0.0430639512439842, -0.0352125116486071, 
    -0.0276581139491196, -0.0197533966267209, -0.0114227063035439, 
    -0.00394647395963456, 0.00352837697832586, 0.0113525599085309, 
    0.0200104767818413, 0.02723829891365, 0.0359199255413451, 
    0.0437271914877151, 0.0505521200449829, 0.0589602520916237, 
    0.0667723680377812, 0.0747974103512355, 0.0812641117460742, 
    0.0897922922848657, 0.0978920928781025, 0.105728137117629, 
    0.113442585454673, 0.121692817309661, 0.129737720385876, 
    0.137595828842102, 0.145064734155323, 0.152994213102405, 
    0.160881233145859, 0.169101679456018, 0.177339269304206, 
    0.185473330155416, 0.193859621633046, 0.201519629954082, 
    0.210118455742516, 0.218249507512367, 0.225704536172217, 
    0.23434772109342, 0.241797075763043, 0.250659873076742, 
    0.259226495087193, 0.267239195350319, 0.276045337972384, 
    0.283492031614052, 0.291470615787073, 0.300988042885703, 
    0.308970863165572, 0.317489435278786, 0.325214522747221, 
    0.333884629873174, 0.343011809486221, 0.350959958775418, 
    0.360275948317332, 0.36825500552018, 0.377503068695314, 
    0.385829582597587, 0.395119769844742, 0.402900316082435, 
    0.41331655914189, 0.422146917021105, 0.431127799631893, 0.44006000632349, 
    0.449009300692515, 0.458375725662631, 0.467177531874324, 
    0.476398019328868, 0.486190233264596, 0.49598785515137, 
    0.505292236225676, 0.515151366677841, 0.524870418207764, 
    0.535264257268931, 0.544583083726188, 0.554661745113796, 
    0.564963940932286, 0.574618992849742, 0.585099818144, 0.595324001346254, 
    0.606001883402227, 0.616469822993688, 0.627535187263527, 
    0.638362578676191, 0.648980837576141, 0.660080652669669, 
    0.671276063508625, 0.682672584803174, 0.694103535479909, 
    0.705893357425493, 0.717374418931897, 0.729337506374243, 
    0.741652464903256, 0.753934360653501, 0.766790546612941, 
    0.779303079373235, 0.7924806061541, 0.805381638744396, 0.81909636862155, 
    0.832939851466389, 0.846827197866773, 0.861150458015298, 
    0.875931275377371, 0.890906541069399, 0.906324073440383, 
    0.922308328383289, 0.938531534954145, 0.955328384713488, 
    0.972730609749026, 0.99076464370209,
  -0.991240839681095, -0.974034143560938, -0.95738466258806, 
    -0.941240309362998, -0.925522782657666, -0.910154716565344, 
    -0.895042416379228, -0.880385431782471, -0.866070024436343, 
    -0.851942966297101, -0.838247925767713, -0.824902069664784, 
    -0.811657178347422, -0.798386313753327, -0.785515894957144, 
    -0.773110167531619, -0.760454053753394, -0.748320493012125, 
    -0.736187345287587, -0.724438402808131, -0.712718519556359, 
    -0.701092889085074, -0.689674382893609, -0.678417968860631, 
    -0.667340557761518, -0.656309895623724, -0.645236003975398, 
    -0.633902116720682, -0.623496000243907, -0.61294608703687, 
    -0.602408556018206, -0.592325577083796, -0.581950086701443, 
    -0.571808770822966, -0.561526319169195, -0.551512742746393, 
    -0.541367520818759, -0.5313608255866, -0.522632627598182, 
    -0.512615173414245, -0.503138078043039, -0.492935673587151, 
    -0.48339686832097, -0.473977837914657, -0.464639535949316, 
    -0.455167620808684, -0.446639430371026, -0.437160199588337, 
    -0.42791535172049, -0.418717984933758, -0.409749215796699, 
    -0.401166814980344, -0.391529186044851, -0.383002892067618, 
    -0.374187415887354, -0.36523831652954, -0.357020072129482, 
    -0.348184701738612, -0.339236725915681, -0.331161868358896, 
    -0.322475159254833, -0.31351457422652, -0.30448652957018, 
    -0.296724077447309, -0.28779276427625, -0.279613297432465, 
    -0.271356667185113, -0.262490171222252, -0.254874203219539, 
    -0.246522942746326, -0.237284293654435, -0.229677056706991, 
    -0.221556304825533, -0.212985888468798, -0.205321164832975, 
    -0.19634802336407, -0.187654735377555, -0.179592360387252, 
    -0.171687103775143, -0.163693692825703, -0.155675000895078, 
    -0.147668123142117, -0.139571630677852, -0.131889648363779, 
    -0.122932465686333, -0.116134731943014, -0.107739626279296, 
    -0.0999006851334197, -0.0918496676128963, -0.0839742640227202, 
    -0.0755084671385028, -0.0674512160162239, -0.0592326380706089, 
    -0.0516907170721861, -0.0441321034076265, -0.03558795299707, 
    -0.0277577548857216, -0.0197716647890261, -0.0117591636450168, 
    -0.00413647978416014, 0.00412256627861376, 0.011935301443709, 
    0.0206252472551031, 0.0275861394224177, 0.0361973113410324, 
    0.0435867478847713, 0.0519410898569536, 0.0599754305879245, 
    0.0673581992228491, 0.0753845389792226, 0.0838483950891943, 
    0.0913344369364864, 0.099792742406966, 0.107825179924186, 
    0.115156044751727, 0.123935991342113, 0.131221170315224, 
    0.140018477971657, 0.147830364876536, 0.155686961358193, 
    0.163994394579271, 0.172341928568483, 0.180197773884884, 
    0.18794649657466, 0.197069872522581, 0.20481486868839, 0.213406208664412, 
    0.221077151598241, 0.229648344885797, 0.238137215364685, 
    0.245830396156955, 0.254183169712089, 0.262697626512874, 
    0.271120244893491, 0.279515655295381, 0.28863505614321, 
    0.296562867230025, 0.305080015516122, 0.31364058711889, 
    0.321668192002237, 0.330778207551232, 0.339134502190745, 
    0.347809748860325, 0.356236833371607, 0.365309731495725, 
    0.373761797303033, 0.382622195308678, 0.391811756172196, 
    0.401272326251477, 0.409979116401858, 0.418706199302485, 
    0.427640785548953, 0.436911923429368, 0.446375917919282, 
    0.455355615221104, 0.46469260680551, 0.473898034966547, 0.48342323724107, 
    0.492540400947848, 0.503135157490717, 0.512136851651649, 
    0.521942237792846, 0.53169070274401, 0.541776313485, 0.551319611854345, 
    0.56142701812417, 0.571193245474652, 0.58154957323712, 0.592123658194136, 
    0.602558039592065, 0.613058608032837, 0.624001109202438, 
    0.634454495103261, 0.644849786953089, 0.656119203482223, 
    0.667064654992253, 0.678325912309037, 0.68956684450242, 
    0.701129172415985, 0.712397554876073, 0.724803426694384, 
    0.736148351614562, 0.748618131553289, 0.760579328827879, 
    0.772969959514889, 0.785756126145524, 0.798273562820538, 
    0.811407249374166, 0.824690336580915, 0.838186493975752, 
    0.85211468081815, 0.866177765973629, 0.880485897211539, 
    0.895051956045583, 0.910152686519438, 0.925373227025153, 
    0.941137048114412, 0.957374646723518, 0.974040768260455, 0.991216501638886,
  -0.991592816388659, -0.975069536017506, -0.958973753994753, 
    -0.943418320905838, -0.92807960116829, -0.913162539702762, 
    -0.89859051750684, -0.884315675364595, -0.870248445532427, 
    -0.856475974193749, -0.842945898926823, -0.829652158958044, 
    -0.816546336087805, -0.803676723861877, -0.790978789808426, 
    -0.778378578298795, -0.76603018579114, -0.754199856734539, 
    -0.741850939306956, -0.730006942834007, -0.718813611316143, 
    -0.707163319238156, -0.695371665577528, -0.684212931074194, 
    -0.673290420455314, -0.662391433868153, -0.651210192540938, 
    -0.640285865249418, -0.630095467320148, -0.619344339563516, 
    -0.60867322508919, -0.598322130210736, -0.588231004777276, 
    -0.57786388804779, -0.568116213213754, -0.557778434482366, 
    -0.547913577934431, -0.538002987829504, -0.527919234170572, 
    -0.518015017428015, -0.508360208275744, -0.499273947316947, 
    -0.489394731810883, -0.480169503058023, -0.470063943679459, 
    -0.460875738693568, -0.451467873309232, -0.442357606717956, 
    -0.433596948431483, -0.424270724862459, -0.414312666213805, 
    -0.405528050659532, -0.396935547353373, -0.387598497628727, 
    -0.379276582716114, -0.370518617284273, -0.361124488445055, 
    -0.35234223995682, -0.34345138918693, -0.335136579331727, 
    -0.32624308630896, -0.31752584874994, -0.309062214803843, 
    -0.300539711812291, -0.291669189563597, -0.283440880389784, 
    -0.274742075709486, -0.265751554006836, -0.257916400066316, 
    -0.249494415281687, -0.24071967390206, -0.232276477775279, 
    -0.223435830049688, -0.215805990680925, -0.207574863152904, 
    -0.199474771521807, -0.191044428968663, -0.182838602411627, 
    -0.174703998508277, -0.166374429054869, -0.158144083013436, 
    -0.150014624179351, -0.141496109350658, -0.133256851538684, 
    -0.125231301422985, -0.117381761647701, -0.10892583476126, 
    -0.100807949763402, -0.0926492525502267, -0.0842047080308511, 
    -0.0767436769266842, -0.0685024652219492, -0.0606155187768198, 
    -0.0528485243417412, -0.0444611488741986, -0.0359542089035497, 
    -0.0284062866707116, -0.0198426137286606, -0.0126001998298151, 
    -0.00351926051403983, 0.00413667035810128, 0.0120233740835229, 
    0.0194072830908185, 0.0285291959139574, 0.035710236563988, 
    0.0437694065307552, 0.0522494802822727, 0.0612390503843099, 
    0.0687290948192431, 0.0769873488285141, 0.0851419225829878, 
    0.092784459453637, 0.101543859005291, 0.10901718309492, 
    0.117386122428708, 0.125249276766235, 0.132832351627566, 
    0.141411727034877, 0.149373368838507, 0.157669765644122, 
    0.16611020393313, 0.174106156754734, 0.182951327580296, 
    0.191135249979716, 0.199196247852639, 0.207456120722814, 
    0.216273379665083, 0.223980718242089, 0.232402938250497, 
    0.240864332431048, 0.248464608875589, 0.257563989044605, 
    0.266018209702062, 0.274510274299859, 0.283052370200077, 
    0.292084745624975, 0.300093910047912, 0.30859251277535, 
    0.317940629592458, 0.326211570608286, 0.335034983666075, 
    0.34320583363186, 0.352607570984055, 0.361116758933535, 
    0.370205862201953, 0.378552923533842, 0.388062835074052, 
    0.39707221042234, 0.405665018239593, 0.414797656253474, 
    0.424118913401548, 0.433339310135824, 0.442469256685249, 
    0.451922760353096, 0.46169501077454, 0.470462222533539, 
    0.479742995130013, 0.489431600163776, 0.498389515961605, 
    0.508317608140939, 0.518058831824593, 0.527880841501288, 
    0.53785632458434, 0.547492955338814, 0.55778025745155, 0.567291336181116, 
    0.577635066665329, 0.587681562376612, 0.597842785690479, 
    0.608364348344543, 0.619318262546884, 0.629643447325867, 
    0.640433329775022, 0.651319797917889, 0.662142432679735, 
    0.673483366693963, 0.684251459311689, 0.695971009529379, 
    0.70709693360342, 0.718651748458858, 0.730197952090835, 
    0.742086501800095, 0.754043425891564, 0.766310001116976, 
    0.778558703411884, 0.790939214090468, 0.80374501911541, 
    0.816594380869222, 0.829687658109691, 0.842923410717923, 
    0.856539701940647, 0.869997593107635, 0.884211870861407, 
    0.898351771640369, 0.91315484970097, 0.928075097591619, 
    0.943382765158495, 0.959016543789923, 0.97504938162602, 0.991591233679223,
  -0.992158268806891, -0.976705923872687, -0.961532153420316, 
    -0.946749089104026, -0.932192052612274, -0.91782520021099, 
    -0.904004730635426, -0.890203693709273, -0.876716715548907, 
    -0.86338884722344, -0.850220439244023, -0.837158598040746, 
    -0.824675620444673, -0.811898797607929, -0.799419060897225, 
    -0.787360574450307, -0.775103839488058, -0.763329670408469, 
    -0.751443810589262, -0.73975218370601, -0.728412257584474, 
    -0.716875015230179, -0.705731348725137, -0.694225524440839, 
    -0.683259937652296, -0.672362063447249, -0.661471109951454, 
    -0.650971586279615, -0.640142976096671, -0.629393721493506, 
    -0.618692806847623, -0.608544865631061, -0.598106575629967, 
    -0.588047989759127, -0.578173285304404, -0.568077156179963, 
    -0.557472859542907, -0.547535139678133, -0.537885452443423, 
    -0.527926278907851, -0.51798138505999, -0.50850679275067, 
    -0.498344962327383, -0.489263051917753, -0.479380154742802, 
    -0.470233211128941, -0.460524804339884, -0.451656970785108, 
    -0.44237678396782, -0.432986389885283, -0.423236583864335, 
    -0.414472748305169, -0.405784146412099, -0.395959956699428, 
    -0.386996975759483, -0.377885020360886, -0.369229542130689, 
    -0.360233670407148, -0.351655637827602, -0.341447550633219, 
    -0.333697770479607, -0.324602749234323, -0.316005934308332, 
    -0.307255656477443, -0.298580874729428, -0.289428757478409, 
    -0.281142302997629, -0.272642296632134, -0.263600993880742, 
    -0.255146510627607, -0.247142498751935, -0.237905913986342, 
    -0.229571664549174, -0.220702717291347, -0.212087558029286, 
    -0.20406645519754, -0.195464568932187, -0.187532685323392, 
    -0.178163163333491, -0.170418472887537, -0.162048077873159, 
    -0.153321858104327, -0.145018426246293, -0.137014091371492, 
    -0.128466100322431, -0.120163234253857, -0.111661638138009, 
    -0.104041201593493, -0.0951276052937488, -0.0866096208549397, 
    -0.0783079426410133, -0.0708273411327681, -0.0618478212119127, 
    -0.053287159408106, -0.0452553372872761, -0.0367065303300212, 
    -0.028393696968131, -0.0207106324762383, -0.012681066342607, 
    -0.0038615690341507, 0.00393797152327626, 0.0122285639541357, 
    0.020683800194019, 0.0286826204338627, 0.0370830677558465, 
    0.0454361295844916, 0.053321622468716, 0.0619655735492202, 
    0.0702179177782279, 0.0785840041183723, 0.0874519171107525, 
    0.095352494136218, 0.103314588957193, 0.111917161283891, 
    0.119925351230129, 0.127781850734597, 0.136218875355114, 
    0.14473709391406, 0.153073610649416, 0.161585526584615, 
    0.170319324686523, 0.177991293634441, 0.186848360120365, 
    0.196093476995734, 0.203889512422892, 0.21221971546494, 
    0.220494793756062, 0.229569747638788, 0.23840086737569, 
    0.246894004555776, 0.254969432832881, 0.263499728363842, 
    0.272374778366832, 0.280772900004717, 0.290144986371402, 
    0.297909150831987, 0.30678629383956, 0.315497186563416, 
    0.324747562520024, 0.334049260094591, 0.341916533749359, 
    0.350781907986222, 0.360331911785119, 0.369268930169068, 
    0.378001194168883, 0.387090601049781, 0.395936928243366, 
    0.405521375120388, 0.413946245625157, 0.423928214905508, 
    0.432649653117085, 0.442123686832083, 0.451251161242766, 
    0.460442509829832, 0.470389043663947, 0.479306627059206, 
    0.489549608034301, 0.498699731593864, 0.507954908930343, 
    0.518049844133901, 0.528375539318149, 0.537636825095062, 
    0.547982947887664, 0.557492257904566, 0.567573841435216, 
    0.577410494365978, 0.58789755944404, 0.598415519422181, 
    0.608639836387702, 0.618689114383389, 0.629406167253361, 
    0.640366184546243, 0.650717151580828, 0.661520627680096, 
    0.672435708413195, 0.683349069129953, 0.694322446751507, 
    0.705449875978802, 0.717025097333311, 0.7282865543114, 0.739875228880794, 
    0.75129722590754, 0.763352099730074, 0.775287320692339, 
    0.787227415473028, 0.799686140101917, 0.811991740894734, 
    0.824616001413798, 0.837483808900172, 0.850120711137762, 
    0.863249989518246, 0.876530453053219, 0.890110105225708, 
    0.903899252570287, 0.917950963394317, 0.932189911392703, 
    0.946759534476296, 0.961573324320965, 0.976695460072638, 0.992159881031145,
  -0.992559943284133, -0.977814942715452, -0.96342146117294, 
    -0.949173238753121, -0.935214644788119, -0.921403281229059, 
    -0.907922926910519, -0.894545049654939, -0.881419175048784, 
    -0.868443267353343, -0.855881733293465, -0.843098740160389, 
    -0.830688725808954, -0.818342975354141, -0.806227773693322, 
    -0.793846915504042, -0.782236807505551, -0.770332112885161, 
    -0.758738805189258, -0.747327516501909, -0.735844520616249, 
    -0.724441489011526, -0.713377874559213, -0.702344004069045, 
    -0.691021962701018, -0.680242571005795, -0.669540248314366, 
    -0.658817153635201, -0.648178704592521, -0.637585283277805, 
    -0.626826455158968, -0.61663180901601, -0.606041071719211, 
    -0.596111760221437, -0.585742004919716, -0.575775940750022, 
    -0.565715237435241, -0.555593569602165, -0.545358428618371, 
    -0.535994881069298, -0.525650649132138, -0.5161848061236, 
    -0.506552327204636, -0.496592622833241, -0.487201414184966, 
    -0.477503470968139, -0.468177599341182, -0.458190551916623, 
    -0.448899101827954, -0.440173540645851, -0.43013132657789, 
    -0.421205449667042, -0.412040556339008, -0.402588828727735, 
    -0.393893746833888, -0.384481715856863, -0.374890913336138, 
    -0.366519663908148, -0.356984081579446, -0.347998060451729, 
    -0.339053682769947, -0.329844334628497, -0.322010401063359, 
    -0.312525958979564, -0.30349554783708, -0.294642957753581, 
    -0.285705914690857, -0.27714954412006, -0.267937480494745, 
    -0.260112326935529, -0.250593237637854, -0.242430811912186, 
    -0.233487752418526, -0.225316913924801, -0.215538365618746, 
    -0.207507901586089, -0.19862403941789, -0.190676953461767, 
    -0.18233885594604, -0.173453340953991, -0.164931310610536, 
    -0.155921102649204, -0.148284358575553, -0.139273569247339, 
    -0.130775066520026, -0.122077246743089, -0.11358329573369, 
    -0.105536268483495, -0.0968214830367635, -0.0887419460485375, 
    -0.0799422041333904, -0.0711404659305965, -0.0632042475567691, 
    -0.0551170927240523, -0.046267489367627, -0.0383004767669875, 
    -0.0292992583198669, -0.0205982639971152, -0.0126977286571323, 
    -0.00458177196874682, 0.00438555819133699, 0.0129324867276516, 
    0.020795613926329, 0.0289644968528131, 0.0372872242333883, 
    0.0461161045627805, 0.0549987751835751, 0.0629264030372845, 
    0.0712947386890833, 0.0802074959111287, 0.0888873285805653, 
    0.0967898251393796, 0.105165279624867, 0.113656663797047, 
    0.122142413516308, 0.131135683431517, 0.139558049497067, 
    0.14748177646554, 0.156447591565037, 0.164663330990875, 
    0.173034849255745, 0.181865868864218, 0.190623273037989, 
    0.199322449032503, 0.207891759260983, 0.216590520779304, 
    0.224451423396369, 0.234157712638254, 0.242061980249078, 
    0.250795358004282, 0.259387526686755, 0.268396406077682, 
    0.276786637807962, 0.286067643190063, 0.295086764351898, 
    0.303662491771773, 0.312044322118699, 0.320830065097566, 
    0.330182712459342, 0.33921446926084, 0.348867613224647, 
    0.357130908220169, 0.366574293060328, 0.375368792938946, 
    0.384434782203294, 0.393995672974346, 0.402932159392301, 
    0.41197659517892, 0.421331325255165, 0.430508403923443, 
    0.439716924874665, 0.449193671383384, 0.458719733581237, 
    0.468313031972419, 0.478178288362638, 0.487220970519106, 
    0.49667325330839, 0.506059784232236, 0.516337987161305, 
    0.526089273456212, 0.53603883364033, 0.545845897703509, 
    0.555630242285416, 0.565521220075441, 0.575643575405821, 
    0.585496581190711, 0.596178768283604, 0.606015857361292, 
    0.616371202221034, 0.626761206085796, 0.637556506526724, 
    0.647912038045973, 0.658530973423253, 0.669444880084157, 
    0.680202966220845, 0.691278047763222, 0.702324664378082, 
    0.713030656642186, 0.724460446288115, 0.735958041281244, 
    0.747444952964149, 0.75861042648676, 0.770513621071816, 
    0.782065321794607, 0.794120085097186, 0.806142136179255, 
    0.818307734895039, 0.830596253660978, 0.843095193924635, 
    0.855708664030812, 0.868521508187656, 0.881485975898988, 
    0.894562097180771, 0.907968899507516, 0.921433611910683, 
    0.935213490613555, 0.949092065055862, 0.963421220348273, 
    0.977837952121192, 0.992564160437886,
  -0.99284682584359, -0.978710329781222, -0.964759339404004, 
    -0.951075611491931, -0.93758133694044, -0.924119657454404, 
    -0.911008541186391, -0.897969913467564, -0.885390181135349, 
    -0.872662896639184, -0.860056321152664, -0.847708868256484, 
    -0.835422252246606, -0.823302326457532, -0.811308980812497, 
    -0.799624497534251, -0.787735884696201, -0.775997529035969, 
    -0.764597569311425, -0.753124481212701, -0.741927326913679, 
    -0.730924818962061, -0.719434514063229, -0.708488364891499, 
    -0.697447816549213, -0.686728364316323, -0.675861528330173, 
    -0.665143432546945, -0.654513155742292, -0.64418367099386, 
    -0.633202376164517, -0.623422463128315, -0.612485515830363, 
    -0.602469270568279, -0.592301470237527, -0.581877844897295, 
    -0.57218401997853, -0.562165913717323, -0.551982562385559, 
    -0.542321876869511, -0.532406116768638, -0.522624176194797, 
    -0.51239653708342, -0.503097686889728, -0.493007991947693, 
    -0.48410027195727, -0.474440565289085, -0.464755658373057, 
    -0.455162937284224, -0.445979504635025, -0.436589030294081, 
    -0.427014896728824, -0.417892478733395, -0.408424333245707, 
    -0.398414651071865, -0.389598766198539, -0.380494947550303, 
    -0.37194404876019, -0.362480606826265, -0.353177852117333, 
    -0.343814034014522, -0.335566081245168, -0.326121456577743, 
    -0.317050375342694, -0.308162010093372, -0.299246396819178, 
    -0.289952314815391, -0.281359404559084, -0.272365722092527, 
    -0.263866481967071, -0.254585977339012, -0.24599546175517, 
    -0.236941739729247, -0.22794397584287, -0.219575595047931, 
    -0.211576241017417, -0.201797573973317, -0.193583407519205, 
    -0.184854215022013, -0.175674428033118, -0.167397513029801, 
    -0.159041168769567, -0.150183047412817, -0.141540917476561, 
    -0.132897121222634, -0.123921740871935, -0.11603563894622, 
    -0.107090867921927, -0.0981142944114582, -0.0893205384700079, 
    -0.0805793140966745, -0.0731611708166824, -0.0643013475211191, 
    -0.0555065584568982, -0.0469906443964098, -0.0384289506790955, 
    -0.0302218032885097, -0.0209397344641743, -0.0127768427382563, 
    -0.00464578906829091, 0.00463404374114444, 0.0127787609233342, 
    0.021445091175227, 0.0302807123328157, 0.0388883659074092, 
    0.0467773198161827, 0.0557683188893841, 0.0642077607916718, 
    0.072498843634985, 0.0808176283878675, 0.0893852781830561, 
    0.0981362396699367, 0.106623096441297, 0.115329118318148, 
    0.124230056434869, 0.132904357403826, 0.141403599293784, 
    0.150444568295305, 0.158512476822989, 0.167758895572628, 
    0.175536171203316, 0.184462574486252, 0.19318978900556, 
    0.201657094406384, 0.21083186044898, 0.219890329730819, 
    0.228279559367548, 0.237025080957649, 0.24621659775802, 
    0.254621690023218, 0.263683812480916, 0.272691104163775, 
    0.281546126064999, 0.290115372488356, 0.299728437615282, 
    0.308162285343379, 0.317361495944119, 0.32625512757896, 
    0.334384685184485, 0.343695145140492, 0.352824500013434, 
    0.362449097760673, 0.371133357995173, 0.380493666240532, 
    0.389827978478543, 0.399217862639248, 0.408006295169348, 
    0.417311371836878, 0.426778531794145, 0.436055829046189, 
    0.446145086817929, 0.455174274626196, 0.465008108023309, 
    0.474514537487431, 0.48362777901147, 0.493233753160225, 
    0.503398492152518, 0.512879512262515, 0.522520558794736, 
    0.53223390100143, 0.542614148909371, 0.552189466322157, 
    0.561941395771794, 0.572188105813632, 0.58225014190315, 
    0.592214539073465, 0.602835723839368, 0.612798541282464, 
    0.623135172570594, 0.633713047684711, 0.64377890493341, 
    0.654197286046694, 0.665221523597231, 0.675852353906517, 
    0.686651006413853, 0.697569362317741, 0.708445746921772, 
    0.719965725985925, 0.730744030226717, 0.74174862836375, 
    0.752851958920954, 0.764692503322575, 0.77608084752103, 
    0.787557387372344, 0.799644292614348, 0.811367971729588, 
    0.82338466202914, 0.835320218318615, 0.847921416590042, 
    0.860034768450684, 0.872593164525527, 0.885297727950199, 
    0.897998823093616, 0.911095260751388, 0.924259230962583, 
    0.937484007788645, 0.951031338197363, 0.964756462567466, 
    0.978713152820973, 0.992848919064886,
  -0.993089472861385, -0.979390599190324, -0.965877536453163, 
    -0.952541462901655, -0.939436063509416, -0.926321168757439, 
    -0.913521308214773, -0.900804198434831, -0.888309769274686, 
    -0.875886322604265, -0.863688155241226, -0.8513578498287, 
    -0.839255413920661, -0.827394675651936, -0.815690908348017, 
    -0.803921498961039, -0.792237785201515, -0.78079800846851, 
    -0.769417155148405, -0.757877490440131, -0.746742735771203, 
    -0.735866726103179, -0.724625254991542, -0.713583653357425, 
    -0.702707634958156, -0.691856660771539, -0.681196203224377, 
    -0.670379799093734, -0.660258371548018, -0.649267675623835, 
    -0.638895128372684, -0.628770713307262, -0.618077370979366, 
    -0.607982875638366, -0.597471243650769, -0.587420505649317, 
    -0.577193508137293, -0.567642146056035, -0.557389739610366, 
    -0.547392759497528, -0.537535067726232, -0.527668139918257, 
    -0.517875787364988, -0.508340721890347, -0.498407087781963, 
    -0.488870260012341, -0.47929954855786, -0.470114621803033, 
    -0.460176544361231, -0.450735215002181, -0.440978627353652, 
    -0.431879162704933, -0.422361121450237, -0.413024766060191, 
    -0.403531346660291, -0.394189098364999, -0.384741368124133, 
    -0.375493080480625, -0.366680180433652, -0.357360577507207, 
    -0.347921206154114, -0.338934779586073, -0.329992004837806, 
    -0.321163779483255, -0.311606682712679, -0.302593253484069, 
    -0.29382329725039, -0.284485060169468, -0.275456493227288, 
    -0.266469004816316, -0.258008861342683, -0.249316475645853, 
    -0.240139957580629, -0.231057344180964, -0.222086789250282, 
    -0.213234536333596, -0.204761542768459, -0.196228559294063, 
    -0.187251588274763, -0.178347785768398, -0.169348580986311, 
    -0.160857101558983, -0.15215687800004, -0.142923422528427, 
    -0.134607197313727, -0.12583917348178, -0.117298695656348, 
    -0.108331495987733, -0.0998770402303109, -0.0907854812484087, 
    -0.0820929179219281, -0.0734551794548024, -0.0647920609500563, 
    -0.0565951915212225, -0.0477592931282102, -0.0393149036073848, 
    -0.0306510637809865, -0.0210360900618276, -0.013483396297227, 
    -0.00447204822682961, 0.00457005585081153, 0.0132886728203735, 
    0.0209164580787642, 0.0305248455265212, 0.0389361421647189, 
    0.0477451546995962, 0.0566348867890812, 0.0647785528969747, 
    0.073022860780685, 0.082332053069804, 0.0907924742851189, 
    0.100097518452116, 0.108460146277156, 0.117054567123696, 
    0.125959306096028, 0.135005966634597, 0.14333415415474, 
    0.151763427693156, 0.160517643587673, 0.169544318740353, 
    0.178096412231876, 0.187298340025777, 0.195879416751568, 
    0.205065068338426, 0.213205162256757, 0.222812478757988, 
    0.230928974499711, 0.240156027465103, 0.248859337240073, 
    0.257898709040547, 0.267245117088982, 0.275919738074426, 
    0.284760423496737, 0.293533429700602, 0.30323412488217, 0.31208485128183, 
    0.320490350601654, 0.330158980493988, 0.339194236675837, 
    0.348531076588687, 0.356784682685575, 0.366493351807794, 
    0.375797444750425, 0.38483949412879, 0.394204925988847, 
    0.403733075790838, 0.412993884908782, 0.422379349764718, 
    0.431455018212156, 0.441201587770212, 0.450638938763379, 
    0.460116028875916, 0.469677522311394, 0.479153259191266, 
    0.488588198068913, 0.498240040174541, 0.508068923605444, 
    0.517968679598625, 0.527817863484007, 0.537408695358405, 
    0.547411260467803, 0.557401278639005, 0.56721632946382, 
    0.577358992096859, 0.587808526485126, 0.597861214029494, 
    0.608242233648603, 0.618068740534666, 0.628737202642922, 
    0.638571460671927, 0.649591066467869, 0.659835719940763, 
    0.670464360382678, 0.681368494514149, 0.69187984091045, 
    0.702779443454258, 0.713541750555843, 0.724871182883401, 
    0.735600939245038, 0.746921393802242, 0.757997117544586, 
    0.769381079108436, 0.780751945445026, 0.792269754174826, 
    0.803684504426267, 0.815518152348206, 0.827352383610143, 
    0.839180035039099, 0.851498325777827, 0.86354196804622, 0.87586664203437, 
    0.888297876410726, 0.900821815771409, 0.913562412952075, 
    0.926400705329411, 0.939359374662437, 0.952548706630848, 
    0.965878863995604, 0.979392435092826, 0.993094748891236,
  -0.993437144314528, -0.98040307780962, -0.967496908261908, 
    -0.954760655939374, -0.942118728638449, -0.929585886525324, 
    -0.917243106059281, -0.904951793121677, -0.892790637485763, 
    -0.880754325085541, -0.868686524186791, -0.857050771351156, 
    -0.845188252985932, -0.833534678860774, -0.822056035126118, 
    -0.810616197083192, -0.798985349572873, -0.787908749604284, 
    -0.776611360424323, -0.765327069336993, -0.754317262311211, 
    -0.743273512293729, -0.732515718443328, -0.72181121380543, 
    -0.710755681757205, -0.700305714218693, -0.689258512526199, 
    -0.678700882754054, -0.668156506556267, -0.658077003793341, 
    -0.647093954344003, -0.637177165316679, -0.626868036364562, 
    -0.616017860195875, -0.606129581804873, -0.595873807669101, 
    -0.585635252321776, -0.576076322083676, -0.56587411152891, 
    -0.555731261423244, -0.545934704053073, -0.535708155445, 
    -0.52632443368225, -0.516035493950476, -0.506407451479841, 
    -0.496717614911278, -0.487242852357526, -0.477584894721732, 
    -0.468229224580086, -0.457983992812251, -0.448627924580807, 
    -0.438917642777345, -0.429828111159238, -0.419901506638681, 
    -0.410483047070473, -0.401032713383497, -0.391854520425423, 
    -0.382449023449246, -0.372881620430689, -0.364355365410233, 
    -0.354690306785077, -0.345757969336753, -0.33595298650432, 
    -0.327275244722318, -0.317689061719446, -0.308718915446053, 
    -0.29944962517153, -0.29001430357135, -0.28128821316241, 
    -0.271720219085565, -0.262877343010448, -0.253606970487277, 
    -0.245015638903701, -0.235655736582083, -0.226893525852653, 
    -0.217476608523732, -0.209051253400438, -0.2001610069362, 
    -0.190772097607824, -0.181993454565428, -0.17305859550321, 
    -0.164507950669927, -0.154773248439308, -0.146001322013461, 
    -0.137331667720623, -0.128238444528031, -0.119460181806269, 
    -0.110327430269446, -0.101904940200967, -0.0928406822473589, 
    -0.0836754961721098, -0.0753835151468916, -0.0662599853835135, 
    -0.0578484055750119, -0.0487676652903338, -0.0397936517774861, 
    -0.0311541922220804, -0.0216092336791416, -0.0131759453287946, 
    -0.00442807341200986, 0.00427755286406891, 0.0130692673504969, 
    0.0222612320498353, 0.0317441068331264, 0.0398414895645453, 
    0.0492072771283941, 0.0572967932346559, 0.0661953745823624, 
    0.0754369599549081, 0.0842742562505947, 0.0922364930127311, 
    0.101309439597657, 0.111087873142816, 0.11934842598401, 
    0.128908738635649, 0.137472753200888, 0.146426713296281, 
    0.155410581239358, 0.163895164017598, 0.17290562962682, 
    0.182038164269308, 0.19125306092197, 0.199193468012907, 
    0.209116640601502, 0.217212764942237, 0.227092962777715, 
    0.235780513051602, 0.244328326936895, 0.253956621451282, 
    0.26266456839434, 0.272062478266034, 0.280985557340683, 
    0.290453873325546, 0.299203669879927, 0.308228527930365, 0.3174235969927, 
    0.326839228244645, 0.336352793391909, 0.34529765004017, 
    0.354571094989722, 0.36423869040062, 0.373198788422189, 0.38281636774978, 
    0.392242496241883, 0.40116193518207, 0.410726955793213, 
    0.420130802799095, 0.429960472353695, 0.439483636322869, 
    0.448442075713018, 0.458175071676684, 0.467853927265335, 
    0.477458495571169, 0.486622552685884, 0.496594572004865, 
    0.506531392598591, 0.516312352846219, 0.52616707182896, 
    0.535910442307284, 0.545835379698001, 0.555821933966839, 
    0.56596803584544, 0.576138031871232, 0.58589190370742, 0.595990976174715, 
    0.606220906869988, 0.616485246986928, 0.626735506797646, 
    0.636853889467487, 0.647420705014266, 0.657813650469662, 
    0.668307101774366, 0.678654986660272, 0.689396908638292, 
    0.699986276408455, 0.71068386749708, 0.721527187769762, 
    0.732360756100534, 0.74342576629933, 0.754355886526489, 
    0.765201103256323, 0.776529801996659, 0.787899556563469, 
    0.79917617315266, 0.810174318767645, 0.821999994720768, 
    0.833622298638239, 0.845155133391957, 0.856988323725206, 
    0.868845158085121, 0.880801441449887, 0.892727867336035, 
    0.904899211350107, 0.917245840247996, 0.929695501032729, 
    0.942080020909184, 0.954756201339399, 0.967504782210566, 
    0.980396926703797, 0.993439560060179,
  -0.99357195233891, -0.98079026166487, -0.968121581637716, 
    -0.955546216466658, -0.943191418471886, -0.930797000707581, 
    -0.918623342225227, -0.906447159670613, -0.894543527209219, 
    -0.882613918395288, -0.870832691155138, -0.859020747620768, 
    -0.847463611796997, -0.835893094103806, -0.824584350398912, 
    -0.813040683280445, -0.801737057341161, -0.79044006081581, 
    -0.779369520850911, -0.768392647022409, -0.757294806167503, 
    -0.746393687647799, -0.735487660187717, -0.72460014387876, 
    -0.713925705175572, -0.703301730226648, -0.692590178567822, 
    -0.68206215784483, -0.671742186810109, -0.661040528623423, 
    -0.650792247576769, -0.640288788358697, -0.629805136624723, 
    -0.619838414863661, -0.609743656729502, -0.599565465008088, 
    -0.589438533346543, -0.579117897323213, -0.56908486954168, 
    -0.559102394166684, -0.549093387218802, -0.539294381908772, 
    -0.529385813725524, -0.519871759848538, -0.509679117134859, 
    -0.499938579157994, -0.489929205529519, -0.480645743218613, 
    -0.470843434535631, -0.461195416800722, -0.451809327678235, 
    -0.442443521162587, -0.432492631497935, -0.423069250007337, 
    -0.413603863153315, -0.404051467037685, -0.394596169626796, 
    -0.384923383869929, -0.376296393227937, -0.366504736469843, 
    -0.357310869906643, -0.347793444480941, -0.338371866012374, 
    -0.32903654286172, -0.320118149953709, -0.3107965022755, 
    -0.301307310908743, -0.29281469785742, -0.283379905918418, 
    -0.274086806497705, -0.265328380510827, -0.256361897001633, 
    -0.246526001426852, -0.237439663537819, -0.22872522556446, 
    -0.219290041128338, -0.210274960469538, -0.201207740179657, 
    -0.191939371597861, -0.183342415600423, -0.173813659294833, 
    -0.165368197134595, -0.15658374994748, -0.147352476896367, 
    -0.138415214034259, -0.129657182413007, -0.120661853797379, 
    -0.111408608528811, -0.102700716207706, -0.0938404919558644, 
    -0.0844663708007978, -0.0757088505787894, -0.0669548687062303, 
    -0.0575876483327843, -0.0487988627052648, -0.0402704608260537, 
    -0.0311038452628929, -0.0221306227904838, -0.0140136180416773, 
    -0.00456359322277087, 0.00447488033511175, 0.0138658708681255, 
    0.0222635104397929, 0.0309175051911923, 0.0397970485218434, 
    0.0488990331112006, 0.0576972776649837, 0.0664404112903877, 
    0.0758141046908005, 0.084501891710764, 0.0931980086316229, 
    0.102810270441386, 0.111893934077809, 0.121034642374563, 
    0.129749229382991, 0.138208634455566, 0.147215916731933, 
    0.155845607195255, 0.165145706207792, 0.174506479770711, 
    0.18369649475005, 0.192342278627221, 0.201163074882523, 
    0.210303223807012, 0.219573858599243, 0.228360734876295, 
    0.237545816838108, 0.246729428859512, 0.256147379784164, 
    0.264716637718142, 0.274009210485576, 0.283197314610982, 
    0.292552080391114, 0.301382567745261, 0.311019621109519, 
    0.319886067223734, 0.329426557888462, 0.338698284941505, 
    0.347755352865594, 0.357538225083085, 0.366399179491241, 
    0.375970271774163, 0.385212243911483, 0.394759767197388, 
    0.404042964172026, 0.413583429037005, 0.423107497097211, 
    0.432721710130083, 0.44213703282684, 0.452060041407799, 
    0.461186264809201, 0.471076697742791, 0.480531508081371, 
    0.490417418571096, 0.500179382908764, 0.509994319692893, 
    0.519859502044269, 0.529340433670014, 0.539213242088661, 
    0.548976229942087, 0.559263224359779, 0.569517237266269, 
    0.578988447638802, 0.589137604011533, 0.599595793009384, 
    0.609299941823048, 0.619473904956974, 0.630160466213848, 
    0.640289398146193, 0.650792058994905, 0.661059446638382, 
    0.671531538116799, 0.682080879395069, 0.692684015367969, 
    0.703374849415592, 0.714131798700945, 0.724700555026801, 
    0.735588684179229, 0.746329050414167, 0.757401281843465, 
    0.768351816115448, 0.779608496676825, 0.790426986792614, 
    0.801811804222466, 0.812988038303232, 0.824458780500032, 
    0.835982490000773, 0.847490639256569, 0.858958324142502, 
    0.870880087677781, 0.882611784365786, 0.894478900821587, 
    0.906493091465884, 0.918682247769331, 0.930809707162745, 
    0.943130489198284, 0.955573916450487, 0.968144924598768, 
    0.980798364218818, 0.993570567567715,
  -0.993670811725793, -0.981107122007405, -0.968635132936609, 
    -0.956256564042192, -0.943992018889023, -0.931868741384798, 
    -0.919853294901609, -0.907832672099897, -0.895922580671829, 
    -0.884148099174846, -0.872618729637424, -0.860965301323443, 
    -0.849476049373765, -0.837988663858334, -0.826679766815968, 
    -0.815198465527969, -0.803965194685049, -0.792849488837784, 
    -0.781811722636107, -0.770846389501056, -0.760032054568606, 
    -0.748907666018835, -0.738146718561044, -0.727298630732475, 
    -0.716712168618386, -0.706248818696633, -0.695156715302857, 
    -0.684702535691644, -0.6744404085132, -0.664176393882422, 
    -0.653507017170565, -0.643200279700954, -0.632924098019182, 
    -0.622514991782093, -0.612600086193565, -0.602424108491834, 
    -0.592235324493045, -0.58208701533427, -0.572034783868958, 
    -0.562198750339083, -0.551856675541021, -0.542349738319261, 
    -0.532481540017823, -0.522536216126315, -0.512834631867154, 
    -0.50316797611197, -0.492939687086535, -0.48315153774182, 
    -0.473517484839574, -0.463826539459284, -0.454466605706625, 
    -0.445088459601359, -0.43527455304038, -0.425870107880441, 
    -0.416291438569229, -0.406738830251205, -0.39739480881695, 
    -0.387715325557316, -0.37841870042783, -0.369296317024603, 
    -0.359368753662443, -0.349726286057132, -0.341028692089011, 
    -0.331602209205701, -0.322258691550744, -0.313136104842328, 
    -0.304022592623885, -0.29432972491378, -0.284966114544855, 
    -0.27601166638528, -0.266549266601634, -0.257557031750055, 
    -0.248662168079912, -0.239103527157298, -0.230007552369053, 
    -0.22087081384867, -0.212367038608537, -0.202805419402979, 
    -0.193819015844346, -0.184619133974507, -0.175476605076861, 
    -0.16655243998803, -0.157444722587247, -0.148264114811287, 
    -0.138917240627132, -0.130457562144887, -0.12119794567625, 
    -0.112203524305217, -0.10339360862365, -0.0941550225359836, 
    -0.0854519742628028, -0.0760198735578923, -0.0676424173378723, 
    -0.0584615599597382, -0.0493432499938493, -0.0403996867528263, 
    -0.0312763213200051, -0.0226449790520623, -0.0135711903909933, 
    -0.00444132023055572, 0.00477330750912166, 0.0134296020779171, 
    0.022062610920177, 0.0319379009288712, 0.040921068869122, 
    0.049361205659372, 0.0582083454240827, 0.0672297296832042, 
    0.0762496642869155, 0.0853113157188298, 0.0943253020277521, 
    0.103465651411185, 0.112550578816327, 0.121305788432309, 
    0.130888694809678, 0.139669665895072, 0.148453278999968, 
    0.157748801700629, 0.166762500262689, 0.175516745752674, 
    0.184876118451137, 0.194120105134258, 0.202663787381928, 
    0.211619245353351, 0.221322268227277, 0.229773491201591, 
    0.239337813815221, 0.24844301703291, 0.257844037162275, 
    0.266989194208904, 0.27603804717424, 0.285154878156114, 
    0.294480223254341, 0.304003462532914, 0.312779857254312, 
    0.322389104083715, 0.331423567345213, 0.340843077356865, 
    0.350018227424749, 0.359840455716675, 0.369023286400975, 
    0.378331198949022, 0.387416405585078, 0.397242492667097, 
    0.406816641322928, 0.416117156653224, 0.425487610205777, 
    0.435176519184111, 0.44489771272219, 0.454565777727078, 
    0.464269990334275, 0.47358144610419, 0.483603162908575, 
    0.492935474205748, 0.503021256493036, 0.512834989867464, 
    0.522422011666885, 0.532284529882801, 0.542050432297141, 
    0.55202232734664, 0.561886563490342, 0.572109999891131, 0.5821819117986, 
    0.592120573960298, 0.60244672850026, 0.612582348369751, 
    0.622685218162058, 0.633022877008565, 0.643176792401692, 
    0.653582480962566, 0.664243715839893, 0.674607931877555, 
    0.684799466536442, 0.695535234191528, 0.705993069493362, 
    0.716835168740258, 0.727359312726633, 0.738172096650772, 
    0.74903524197002, 0.759862790928403, 0.770779590094274, 0.78173243956202, 
    0.793105711993139, 0.803982104858324, 0.815309927149123, 
    0.826541928897584, 0.837911020927421, 0.849492506033205, 0.860968285161, 
    0.872508740962136, 0.884236254501981, 0.896003853930202, 
    0.907867304970846, 0.919820664888985, 0.931820970454318, 
    0.944035689245635, 0.956238842113792, 0.96864161083502, 
    0.981109013005454, 0.993678322205219,
  -0.993852857989574, -0.981620519339406, -0.969443501387105, 
    -0.957391751820713, -0.945466363599336, -0.933568128247873, 
    -0.921726273716227, -0.910149235092955, -0.898488108747968, 
    -0.886780416605524, -0.875360013887673, -0.864060725718747, 
    -0.85262007288261, -0.84126056964499, -0.830129571640335, 
    -0.818824545866127, -0.807911846293757, -0.796866448127758, 
    -0.785860359232445, -0.77496964201067, -0.764133239377303, 
    -0.75334150997459, -0.742589025626488, -0.731687937943123, 
    -0.7210663600657, -0.710530524927516, -0.699952764018968, 
    -0.689703152266832, -0.679201686585471, -0.668804002147194, 
    -0.658562547659324, -0.647942422049377, -0.637747034381689, 
    -0.627409490108964, -0.617317348699358, -0.607242941543508, 
    -0.59706022895003, -0.587009607878566, -0.57715035082852, 
    -0.566879111587897, -0.556661119409999, -0.547276261200233, 
    -0.537114281332654, -0.527060776260125, -0.517489399778982, 
    -0.507571890638964, -0.497476363082569, -0.487924508396762, 
    -0.478128825674651, -0.468486309473039, -0.458766226921355, 
    -0.449469818437267, -0.439790398155251, -0.429989786869963, 
    -0.420288537611205, -0.410829474662787, -0.401505930848562, 
    -0.39169275302102, -0.382245185913884, -0.372992533424047, 
    -0.363269613932157, -0.353993499587144, -0.344380930564907, 
    -0.335099633350338, -0.325790632839966, -0.31644195712416, 
    -0.307234635859128, -0.297804435379563, -0.288175162870419, 
    -0.279092422231157, -0.269960361805289, -0.260615744740455, 
    -0.251443396308174, -0.242030172359077, -0.232626828443045, 
    -0.22350858382369, -0.21475135420141, -0.20512267721535, 
    -0.195993700231955, -0.186954885706376, -0.177801664163453, 
    -0.168224011054189, -0.159102456062424, -0.149773494499242, 
    -0.141119765967355, -0.131795111892101, -0.122870459204468, 
    -0.11374038457884, -0.104798316882281, -0.095328287797785, 
    -0.0864773438149466, -0.0773786536721297, -0.0679245509578405, 
    -0.0588824111530857, -0.0499029903476317, -0.0409643694990185, 
    -0.0319715417945569, -0.022505632457377, -0.0133993973516746, 
    -0.00474581687054433, 0.00447744037650955, 0.0135596657287461, 
    0.0226881523014374, 0.0317537047721388, 0.0410177556602205, 
    0.0498555141071513, 0.059367331898751, 0.0678430201694437, 
    0.0771332161331945, 0.0863317110361446, 0.0951310801775719, 
    0.104618732010171, 0.113847469748204, 0.123004734312049, 
    0.131969468864865, 0.141091269766544, 0.150239169672527, 
    0.158949520672679, 0.168205931877891, 0.177552325083774, 
    0.187039970057886, 0.195978141417996, 0.204829797445145, 
    0.214424737170195, 0.223935298314924, 0.232442322572898, 
    0.242140941633652, 0.251377050901988, 0.260362313413228, 
    0.269912393939022, 0.278923029172262, 0.288385466518485, 
    0.296994076051947, 0.306718663624281, 0.316401309239124, 
    0.325632857401768, 0.33479312877339, 0.344685046088172, 0.35363129344609, 
    0.363354544818768, 0.372919979696735, 0.382265228452202, 
    0.391704560424075, 0.401413393071713, 0.411016679393084, 
    0.420636128563653, 0.429969747115961, 0.439432509974263, 
    0.449150708121146, 0.45898957767295, 0.468416473037022, 
    0.478207420716979, 0.488054541288682, 0.497341057775207, 
    0.507367850179087, 0.517548542180051, 0.52716315314188, 
    0.537026307341295, 0.546672595793068, 0.556863026826954, 
    0.566790742988008, 0.576989429724143, 0.586993402019585, 
    0.597445034748053, 0.607272931803127, 0.617345568726304, 
    0.627803449275518, 0.63782130668633, 0.648057025525614, 
    0.658276326592008, 0.668602530406075, 0.678942805576936, 
    0.689525430175061, 0.700023941823082, 0.710704469220697, 
    0.721089198042184, 0.731677576640946, 0.742609123605689, 
    0.753328644051119, 0.764150684268002, 0.774920189483912, 
    0.78602275833649, 0.796824010424352, 0.807795357794876, 
    0.818918740804981, 0.830126518217746, 0.841445711687319, 
    0.852561509028703, 0.863916465860213, 0.875371395972019, 
    0.886890220484922, 0.898478642553966, 0.910120448524871, 
    0.921736036588369, 0.933569436667159, 0.945471556642625, 
    0.957419458103052, 0.96946833829445, 0.981607076396915, 0.993845036343051,
  -0.99399235586758, -0.982009093952408, -0.970111511304203, 
    -0.958282287737963, -0.946537960758367, -0.934864956370653, 
    -0.92331537956771, -0.911746911177809, -0.900274175069531, 
    -0.888961013908183, -0.877438635177484, -0.866290785177248, 
    -0.855147033249116, -0.843898293221713, -0.832861073115296, 
    -0.821693146315049, -0.810882014685805, -0.799842055252876, 
    -0.788781474884853, -0.778151628041193, -0.767471717082435, 
    -0.756690628080431, -0.746063866082679, -0.73531082814878, 
    -0.724730897020067, -0.714143645820058, -0.703782034796291, 
    -0.693368151835425, -0.682889814548257, -0.672490852996383, 
    -0.662056970239644, -0.651765016097378, -0.641548062393773, 
    -0.631124059120198, -0.620950019199411, -0.61109630167239, 
    -0.601032126553342, -0.590585139380302, -0.580940220173522, 
    -0.570813239257826, -0.561105285478828, -0.550614697055401, 
    -0.541144260575422, -0.531067317550055, -0.521301922242751, 
    -0.511445882610499, -0.501497751324635, -0.49156942908241, 
    -0.481826242712148, -0.472159428958111, -0.462142800009537, 
    -0.452699104014021, -0.442973233139249, -0.433496163693806, 
    -0.423540610640799, -0.414405934090092, -0.404447762912622, 
    -0.394856697857161, -0.385717051030058, -0.376067614206125, 
    -0.36648776540551, -0.356931047936415, -0.34731981401247, 
    -0.338072615916586, -0.328434568207003, -0.319255023862721, 
    -0.31005520505747, -0.300359329614449, -0.290849343112344, 
    -0.281887823836565, -0.272355519667085, -0.262609439352727, 
    -0.253511083017009, -0.244116996886719, -0.234580290647235, 
    -0.225942364029265, -0.216624987225704, -0.207221858697227, 
    -0.197625242349703, -0.188417104677424, -0.179286171680999, 
    -0.170065601864609, -0.160991795991372, -0.151693560457002, 
    -0.142158069238132, -0.133079323448332, -0.123843506316451, 
    -0.114645115973885, -0.105610994296687, -0.096109207145507, 
    -0.0872776458146735, -0.0780221243964431, -0.0690131283226568, 
    -0.0590819333523119, -0.0509397491993543, -0.0409465782536978, 
    -0.031858454108904, -0.0227960397428999, -0.013826143770519, 
    -0.00476303074849872, 0.00469050586384981, 0.014066423834374, 
    0.0229767948167355, 0.0323113830261886, 0.0412959109825173, 
    0.0503309306219801, 0.0596272076629069, 0.0687580579416872, 
    0.0779492372088297, 0.0869081337496139, 0.0964762188921094, 
    0.105323492623897, 0.11450956124289, 0.123990664638806, 
    0.133200356930838, 0.142187147900271, 0.151811012938937, 
    0.160529713909059, 0.170062946067894, 0.179295986451253, 
    0.188237681109778, 0.197879300390116, 0.207135355205087, 
    0.216464628421383, 0.225630062655279, 0.23487198163629, 
    0.244422558157467, 0.253811380728611, 0.263050784980011, 
    0.272139185755195, 0.281427906375785, 0.290988442019537, 
    0.300437101862713, 0.309731344872939, 0.318790382474367, 
    0.328664734559257, 0.338003809413467, 0.347067298350039, 
    0.356816169075007, 0.36634261226927, 0.376189822698112, 
    0.385710306492726, 0.395035911437338, 0.404830200606832, 
    0.414131362821442, 0.424018897384756, 0.433622361166683, 
    0.442873285647318, 0.45284404813696, 0.462312760182079, 
    0.472108632580791, 0.481880533975669, 0.491888359915912, 
    0.501356855383211, 0.511309296358555, 0.521017180039036, 
    0.531027574433875, 0.540930316499287, 0.550768210783453, 
    0.560858163049437, 0.570928811754404, 0.580731025853349, 
    0.591060382178877, 0.600893544505069, 0.611105528789681, 
    0.621254233176041, 0.631379414201468, 0.641696041877454, 
    0.65195626583201, 0.662135444217923, 0.672530233220422, 
    0.682868703873262, 0.693272768070603, 0.703628035577276, 
    0.71442164904163, 0.724816600581015, 0.735514806465542, 
    0.746093753097109, 0.756766575504045, 0.767254342182294, 
    0.778035204518034, 0.789046812754134, 0.799758411866511, 
    0.810936891562997, 0.821731804442874, 0.832805119163806, 
    0.843845728097376, 0.855184184018753, 0.866315200047299, 
    0.877597505581322, 0.888889848456739, 0.900269443629478, 
    0.911679574633866, 0.923225546194738, 0.9348267154246, 0.946576685468896, 
    0.958292198836739, 0.970114386496548, 0.982012781218649, 0.993990616291913,
  -0.9940898855687, -0.98232405265742, -0.970622843063481, 
    -0.958945875830684, -0.947419981703779, -0.935935997271335, 
    -0.924446676912607, -0.913133078186143, -0.901742254469617, 
    -0.890435139000586, -0.87929139351304, -0.86817063461093, 
    -0.857029614553182, -0.846037507275588, -0.83503323154788, 
    -0.824087025906733, -0.813134546405457, -0.802344560737853, 
    -0.791572290370135, -0.780716763744614, -0.770193893761511, 
    -0.759425925152101, -0.748855515440058, -0.738249219722366, 
    -0.727803007099966, -0.717310204791889, -0.706743550551873, 
    -0.696112829440055, -0.685975022156664, -0.675509709903944, 
    -0.665321727026555, -0.655192494558228, -0.644846985592488, 
    -0.634478952312105, -0.624391297746727, -0.614106778004095, 
    -0.604303177029702, -0.594084144122313, -0.583939881474858, 
    -0.573986337914203, -0.563953545559472, -0.553753897475849, 
    -0.544266411061014, -0.534240416831516, -0.524274951266498, 
    -0.514538348841025, -0.504469441724419, -0.494483242109683, 
    -0.485124041623586, -0.475176978083076, -0.465469191282809, 
    -0.455863256543611, -0.445866299364569, -0.436229425854331, 
    -0.426380129248682, -0.416796855460011, -0.407219645611237, 
    -0.397665917037624, -0.388059007070732, -0.378652867823975, 
    -0.369335468855368, -0.35960627396829, -0.349914993971318, 
    -0.340462741310535, -0.330561693685084, -0.321782687090787, 
    -0.311879087874603, -0.302137226550708, -0.292720725143666, 
    -0.283548984094091, -0.274414495063257, -0.265214706877156, 
    -0.255492339149546, -0.24587295672067, -0.236799885051085, 
    -0.227237577348646, -0.218336621197, -0.208572063929451, 
    -0.199166109496116, -0.189989043183618, -0.180615814389846, 
    -0.17147300254926, -0.162175231686044, -0.152558181215651, 
    -0.143128206233251, -0.134487053202583, -0.124740786973747, 
    -0.115803321189014, -0.106329009142155, -0.0967292034942328, 
    -0.0879173290129833, -0.078200838379786, -0.0694209622392746, 
    -0.0605789402753451, -0.0506139555397783, -0.0414547839810814, 
    -0.0321215585578779, -0.0231539393242452, -0.0137530941563338, 
    -0.00443773737683175, 0.00438240340012489, 0.0137742180878844, 
    0.0228427359028806, 0.0323192026958473, 0.041944319070984, 
    0.0507235337217357, 0.0599348549519362, 0.0691076260853019, 
    0.0784054354504138, 0.0878099593565607, 0.0969770256251587, 
    0.106620538426189, 0.115582854774154, 0.124751818515898, 
    0.134237080434411, 0.143504046838729, 0.15291470330169, 
    0.161857791302094, 0.170850786857698, 0.180403976108759, 
    0.189867548113477, 0.199888724494592, 0.208293675292732, 
    0.217853868503605, 0.227459749900463, 0.23650164169056, 
    0.245761007830408, 0.255515978498165, 0.264932556114403, 
    0.274630467631409, 0.283785078297937, 0.293067664438147, 
    0.302336132341768, 0.311826888830434, 0.32124882847816, 
    0.330812498299912, 0.340028594428648, 0.349991365534671, 
    0.35955215201795, 0.368776593474745, 0.378687383466799, 0.38824751635533, 
    0.39762695618611, 0.407155708920637, 0.417406732485129, 
    0.426717922054122, 0.436131492652553, 0.445997565639311, 
    0.455493963710728, 0.465434361293542, 0.474900564292472, 
    0.484653453214709, 0.494793588086752, 0.504845300306157, 
    0.514374399490023, 0.524172838367414, 0.534263127634698, 
    0.544143452155127, 0.553937421651125, 0.564098408283114, 
    0.573831342150765, 0.58381395506079, 0.594037977494027, 
    0.604259650219811, 0.614145147493818, 0.624359114596097, 
    0.634398618391905, 0.644782833347004, 0.654962115101154, 
    0.665279407112887, 0.675427784745398, 0.686068492406556, 
    0.696328412923823, 0.706496229791895, 0.717203498102404, 
    0.727624330820427, 0.738193290851427, 0.748838107834687, 
    0.759533414372086, 0.770069654021024, 0.780865676631971, 
    0.791621256109808, 0.802335380299534, 0.81310346296179, 
    0.824030114977176, 0.835112698562594, 0.845925503499704, 
    0.857191809271118, 0.868139608999217, 0.879336055719169, 
    0.890476986651188, 0.901705645442151, 0.913121747913099, 
    0.924488666786992, 0.935903503719839, 0.947386257493916, 
    0.958999672373446, 0.970628160230369, 0.982312909555019, 0.994095530489521,
  -0.994180320116048, -0.982578373345538, -0.971051430374406, 
    -0.95953604490674, -0.948094198010165, -0.936774919519556, 
    -0.925473360658044, -0.914219499268652, -0.903015295522967, 
    -0.891813010198907, -0.880791419878959, -0.86956075067575, 
    -0.858618175069742, -0.84768636459257, -0.836804848578638, 
    -0.826079989265911, -0.815112864356245, -0.80435258858126, 
    -0.793582423536753, -0.782945136487983, -0.772227640337976, 
    -0.761552428218736, -0.751120537643256, -0.740452368042143, 
    -0.73020735498293, -0.71962316548031, -0.709175616194236, 
    -0.698766729162634, -0.688500683849696, -0.678168464935944, 
    -0.667835193906051, -0.657364565661113, -0.647473219429412, 
    -0.637341700569629, -0.627274733217717, -0.616737524685603, 
    -0.606787320176663, -0.596741024262475, -0.586265581283538, 
    -0.576439951953674, -0.566443502575309, -0.556630145546609, 
    -0.546712543413477, -0.53694339976451, -0.526627252671243, 
    -0.517154086725352, -0.506808746313492, -0.497319450288127, 
    -0.487287876281457, -0.477525892769509, -0.467787304018641, 
    -0.458160373634678, -0.448366828891194, -0.438605051751478, 
    -0.429107165713119, -0.419454617406483, -0.409454638822187, 
    -0.39999573199533, -0.389970707213413, -0.380641828135114, 
    -0.371105062563182, -0.361374995569867, -0.352113575389522, 
    -0.342503248773102, -0.332633367955105, -0.323545098636832, 
    -0.314020172287506, -0.304261825926332, -0.294676739316088, 
    -0.285438484256986, -0.275546277279396, -0.26641277547105, 
    -0.256938324320682, -0.247466761003162, -0.238718904579619, 
    -0.228488803414101, -0.219469113395999, -0.210178703091471, 
    -0.200773528222765, -0.191172268372426, -0.181533078219445, 
    -0.17272137305191, -0.16302340136269, -0.153744876188885, 
    -0.144030324085835, -0.135201679295775, -0.125623830217475, 
    -0.116507275735999, -0.107009100663897, -0.0976118248885627, 
    -0.0887538248691111, -0.0787636855056859, -0.0693872570943232, 
    -0.0602168860356512, -0.0511775951571192, -0.041966657686492, 
    -0.0324850121577763, -0.023267380983556, -0.0140766602099245, 
    -0.00471058778601602, 0.00475322025053029, 0.0141883514867603, 
    0.0233406291647012, 0.0325577918093713, 0.0417987153081216, 
    0.0511948179130562, 0.0607083280343173, 0.0697248857059957, 
    0.0791397380462086, 0.088278199771381, 0.0979625762291091, 
    0.106948018492396, 0.116137575703697, 0.125819965337221, 
    0.134752503192672, 0.144727242927343, 0.153188463716417, 
    0.163311817353436, 0.172398061932959, 0.181802450894881, 
    0.191318447789662, 0.200678577224805, 0.209837445621071, 
    0.219344696622245, 0.228556025829019, 0.238486287506076, 
    0.247470358098497, 0.256929662182698, 0.266431117074523, 
    0.275811973699619, 0.285349500724362, 0.294999109519159, 
    0.304333945457753, 0.313865950024548, 0.32323037474304, 
    0.332961028198794, 0.342542507389664, 0.352127033816236, 
    0.361426608283477, 0.370977159456176, 0.380734101198373, 
    0.390393608204466, 0.399755298355038, 0.409686747529327, 
    0.419226456310846, 0.428877240492472, 0.438448929327004, 
    0.448419003080174, 0.458127345802956, 0.467770723855046, 
    0.477564178244451, 0.487254094591812, 0.497377772216655, 
    0.507294768222743, 0.517110219542317, 0.526667729022375, 
    0.536682382599613, 0.546552731242419, 0.556758920389262, 
    0.566454625490876, 0.57637237730526, 0.586665069686775, 
    0.596694343406572, 0.606825193559027, 0.616744110929265, 
    0.626970286252167, 0.637231638181578, 0.647435528668661, 
    0.65748678739814, 0.667947916248285, 0.678107083177262, 
    0.688384615815951, 0.698747372128915, 0.709224348894518, 
    0.719987581127962, 0.730072348146959, 0.740515987577642, 
    0.751117431083585, 0.761778340941019, 0.772373910135216, 
    0.78295388128022, 0.793468232247318, 0.804456634122361, 
    0.815206699946773, 0.825998729020638, 0.83684546677294, 
    0.847831958002796, 0.858740993026943, 0.869656213024215, 
    0.880738728209338, 0.891899876827953, 0.903048931787986, 
    0.914219886830299, 0.925437032772961, 0.936743028292809, 
    0.948131440199671, 0.959542371265991, 0.971044165523127, 
    0.982573183154855, 0.994179684393818,
  -0.994205251197892, -0.982630677512829, -0.971128030124449, 
    -0.959657269102974, -0.948295283762373, -0.936940285911383, 
    -0.925676114642262, -0.914495463919707, -0.903262619606647, 
    -0.892188384753987, -0.881067675994507, -0.870040956536965, 
    -0.859005928057763, -0.848084614028688, -0.837184864519869, 
    -0.826482744310908, -0.815536410692628, -0.804889764131382, 
    -0.794071176683209, -0.78348740644839, -0.772750250151836, 
    -0.76231217489835, -0.75152329008605, -0.741076495542544, 
    -0.730593364697267, -0.720146442319556, -0.709564545191388, 
    -0.699248432812516, -0.689010598271537, -0.678953375288736, 
    -0.668551508136, -0.658254420392505, -0.64791810127212, 
    -0.637737164293283, -0.62757327001002, -0.617493491679924, 
    -0.607239123236257, -0.597066006030868, -0.587318187015155, 
    -0.577270039191044, -0.566917346407535, -0.55719535924372, 
    -0.547101572000369, -0.537553468120404, -0.527295201803381, 
    -0.517580076345698, -0.507451312298588, -0.497628049768983, 
    -0.48806038312695, -0.478276841246444, -0.468448141083259, 
    -0.458488312910277, -0.448872880013699, -0.439140731751204, 
    -0.429277395570733, -0.419907714016697, -0.410269349751845, 
    -0.400393118459354, -0.390615284874399, -0.381494709523079, 
    -0.37137953290017, -0.361947106128128, -0.352424491994542, 
    -0.342716634927135, -0.333225358580109, -0.323820653479012, 
    -0.314319635753061, -0.304670063832776, -0.295291004023768, 
    -0.285724665317765, -0.276312102071261, -0.266946780846963, 
    -0.257478863880987, -0.248079826025228, -0.238460545826383, 
    -0.229005087881063, -0.220017789811426, -0.210208986734575, 
    -0.200789943181123, -0.191770109735835, -0.181826483062971, 
    -0.172269856457951, -0.163124648237523, -0.153674047075521, 
    -0.144905487248568, -0.135202186384465, -0.125631329723294, 
    -0.116575119747083, -0.106946259766435, -0.0977460177559602, 
    -0.0885853869728377, -0.0794917432070585, -0.0699410500365746, 
    -0.0608343104401409, -0.0511458103418556, -0.0420526316972344, 
    -0.0328655949421407, -0.0230343319818862, -0.013895991077369, 
    -0.00463507814140766, 0.00492075819718679, 0.0138256081389213, 
    0.0233927867204663, 0.0326095016207166, 0.0421306503671489, 
    0.051206833205636, 0.0605540328714566, 0.0699432508783909, 
    0.0791664204484631, 0.0882930674338234, 0.0982460942022292, 
    0.107132685110504, 0.116496894690028, 0.125919317967764, 
    0.135354753641078, 0.144699238460606, 0.15402603962917, 
    0.163169325151132, 0.172622601638774, 0.181944807598143, 
    0.191379637232123, 0.200448553558979, 0.210232063557631, 
    0.219744187050915, 0.229354053161611, 0.238406955831336, 
    0.248555437468114, 0.25750873833031, 0.267147579746965, 
    0.276041271677846, 0.285695471267484, 0.294982993017815, 
    0.304670705622612, 0.314159715859064, 0.323576443526542, 
    0.33303333750086, 0.342738652639668, 0.352106443346377, 0.36197139753281, 
    0.37154686795255, 0.381136006531501, 0.390628936745173, 
    0.400509795304305, 0.410082023712298, 0.419854302734479, 
    0.429517475095425, 0.439206666727916, 0.448875055333726, 
    0.45877321622914, 0.468687539605844, 0.478067544890893, 
    0.487924422302178, 0.497926572922735, 0.507946922310652, 
    0.517345712681434, 0.527390940820316, 0.537232485581665, 
    0.547157746292512, 0.556906399897445, 0.56712707243563, 
    0.577308702035581, 0.587015696239409, 0.597221439639825, 
    0.607424073374717, 0.617250882990905, 0.62762251359641, 
    0.637649687596386, 0.648018728526026, 0.657970229860586, 
    0.668106511712429, 0.678609117404228, 0.688937882431056, 
    0.699381413278516, 0.709735143659181, 0.720186121482939, 
    0.730556292335146, 0.741073983363587, 0.751754498495295, 
    0.762147652551858, 0.772748865767221, 0.783451274250173, 
    0.794100092086412, 0.804741557740932, 0.81553243721442, 
    0.826477298438087, 0.8372542029519, 0.848042410962537, 0.859087025696858, 
    0.870056100752622, 0.881032120375082, 0.89211283806936, 
    0.903221614404977, 0.914444487637105, 0.925717324249837, 
    0.936932042387161, 0.948292758793886, 0.959660358874437, 
    0.971122171831697, 0.982633133477723, 0.9941956946729,
  -0.994215810249361, -0.982688933042893, -0.971175041984606, 
    -0.959775096621377, -0.948480357617225, -0.937122099831545, 
    -0.925846980528595, -0.914704448919362, -0.903464823649012, 
    -0.892373986355242, -0.88137600607143, -0.870324994445397, 
    -0.859386525559334, -0.848523589366369, -0.83761201926173, 
    -0.826831639617237, -0.816034951979508, -0.805289822113661, 
    -0.794477429734437, -0.783926276592683, -0.77328943711815, 
    -0.762655430162049, -0.752160527070841, -0.7415670288688, 
    -0.731225151370713, -0.720720275120769, -0.710231813286875, 
    -0.699828130875022, -0.689534704390932, -0.678987607369597, 
    -0.668873398670539, -0.658625972746599, -0.648616464874681, 
    -0.638127028650339, -0.628164831178385, -0.617997427411913, 
    -0.608049691748643, -0.598048436292705, -0.587501911579996, 
    -0.577744477206771, -0.567868959943476, -0.557787525510299, 
    -0.547848514226456, -0.53792491570515, -0.527799415882695, 
    -0.517857230610947, -0.508331096963804, -0.498119348145647, 
    -0.488323201425878, -0.478812012459952, -0.46880993113085, 
    -0.459164280452315, -0.449209218047378, -0.439835365671032, 
    -0.429967138965381, -0.420069962758632, -0.410536581335349, 
    -0.400806895820297, -0.391349102820511, -0.381510352168201, 
    -0.371864012688361, -0.362464176582759, -0.352653623815045, 
    -0.343430083358811, -0.334053561218669, -0.323973794673924, 
    -0.314359330331291, -0.305515604004818, -0.295754077045609, 
    -0.28628047244064, -0.276795627013524, -0.267039301721266, 
    -0.257736151451469, -0.248373516647259, -0.238430940890602, 
    -0.229366094998011, -0.219848741781235, -0.210360304443203, 
    -0.201297187125291, -0.191658807962178, -0.182211864809878, 
    -0.173140757069909, -0.163512364053875, -0.154318528821079, 
    -0.144806584466411, -0.135308339146443, -0.125770922352138, 
    -0.11674845402398, -0.107414621473604, -0.0981255595787839, 
    -0.088653252516577, -0.0795203441097797, -0.0697658586862902, 
    -0.0605680405039837, -0.0511230309424852, -0.0420204713727906, 
    -0.0325038270017554, -0.0232828390253435, -0.0140916545271526, 
    -0.00448245603926831, 0.00456124969540251, 0.0140752659778364, 
    0.0233344571546968, 0.0328803607016116, 0.0419580468272549, 
    0.0514285328231682, 0.0604998298851272, 0.0700871978716614, 
    0.0794576349679901, 0.0885360489965268, 0.0976701068084981, 
    0.107233763786332, 0.116840418587431, 0.125883411552956, 
    0.135581263795838, 0.144989631796557, 0.154292801291917, 
    0.163517564910292, 0.17283569429194, 0.182255916290571, 
    0.191712334988847, 0.201117942260872, 0.210837599967794, 
    0.220061157731801, 0.229517942141437, 0.238790102304918, 
    0.248171469066108, 0.257819224936982, 0.267082765922937, 
    0.276552543243109, 0.286323952143953, 0.295608940409258, 
    0.305219653826442, 0.314519956155112, 0.323974968366787, 
    0.33364854593855, 0.3431132378295, 0.352427249135702, 0.362643114411149, 
    0.371815916783682, 0.381631006954823, 0.391468649838047, 
    0.400901666300573, 0.410574805120226, 0.420225499258323, 
    0.430034584551253, 0.439895576984801, 0.449595106494009, 
    0.458891281871567, 0.468942401441356, 0.47848992495238, 
    0.488260102076409, 0.498439272329726, 0.507974964116276, 
    0.518146547730272, 0.527998815033236, 0.537901476917677, 
    0.547849419981732, 0.557627583686919, 0.56751473129201, 
    0.577821529940944, 0.587945290269864, 0.597531588615629, 
    0.607992679854752, 0.617975045726882, 0.628221785459578, 
    0.638494054789943, 0.64842832345788, 0.658737916985252, 
    0.668714251529959, 0.679192511510977, 0.689460458618056, 
    0.699954485534454, 0.710201777109464, 0.720597033588786, 
    0.731035512464489, 0.741546663200275, 0.752089299451543, 
    0.76280264045933, 0.773271643223385, 0.783890416889918, 
    0.794585547955372, 0.805279439572211, 0.81597727753715, 
    0.826671583812377, 0.837374794881697, 0.848547157317635, 
    0.859383858681737, 0.870369933004034, 0.881343014075309, 
    0.892462281173214, 0.903509527495866, 0.914649535033316, 
    0.925848031025777, 0.937133917582796, 0.948407707505814, 
    0.959817167940818, 0.971210982439852, 0.982677550295914, 0.994215221584715,
  -0.994251058626677, -0.982777640041624, -0.9713754361327, 
    -0.960020371865999, -0.948741139075352, -0.937454114444355, 
    -0.92625608584296, -0.915145397946785, -0.903958526076652, 
    -0.893022601707041, -0.881898188074008, -0.871030966294071, 
    -0.859908279641674, -0.849139073161801, -0.838303472305174, 
    -0.827528706505704, -0.816714939499625, -0.806150290138213, 
    -0.795419119925642, -0.78467809600162, -0.774185974789098, 
    -0.763554297882127, -0.753010870820941, -0.742579176523943, 
    -0.731916428390258, -0.721776703055971, -0.711132909805687, 
    -0.700781865055668, -0.690648609061863, -0.680220641558305, 
    -0.66999085424538, -0.659943908948568, -0.649570020560331, 
    -0.639198522688516, -0.629102051556337, -0.619086414409087, 
    -0.608988369824454, -0.598762673774623, -0.589113034670128, 
    -0.578800731053994, -0.568875316322454, -0.558794721890305, 
    -0.548742595439479, -0.53872571133792, -0.529070802501346, 
    -0.518936057315577, -0.509016729340018, -0.499430626923155, 
    -0.489583204349042, -0.479725197211033, -0.469969102767223, 
    -0.460282237710495, -0.450422037426781, -0.440641753605136, 
    -0.430901968431268, -0.421222848231307, -0.411924545716873, 
    -0.402058573877122, -0.392231020023687, -0.382428847025854, 
    -0.373048196848851, -0.363426498965524, -0.353731256067548, 
    -0.344403386754764, -0.33453435873011, -0.324843011820605, 
    -0.315451819334052, -0.305575507229621, -0.295962939309843, 
    -0.28664487910305, -0.277426870632625, -0.267896528292416, 
    -0.258606891826944, -0.248792631847293, -0.239475364765111, 
    -0.229797424956071, -0.220468952030069, -0.211251072400609, 
    -0.201846709642275, -0.192105029945751, -0.18310899685908, 
    -0.173478496782745, -0.164183412438588, -0.154567670943362, 
    -0.145325203318513, -0.135671396023033, -0.125989125727909, 
    -0.117076073742988, -0.107662102221431, -0.0986357627845401, 
    -0.0891287940707045, -0.0794394164037493, -0.0701929480095626, 
    -0.0609666177901873, -0.0513380862016951, -0.0418253749485021, 
    -0.0329611753471765, -0.0233935228721137, -0.0140224355053873, 
    -0.0046843298912887, 0.00446037741644204, 0.0141751815978044, 
    0.0238728407254441, 0.0328302635958499, 0.0419467834698059, 
    0.05140440681788, 0.0609517073595973, 0.070315160422087, 
    0.0794168926444618, 0.0888581141198221, 0.0983887897207404, 
    0.107766674880514, 0.11697377412025, 0.126084727402415, 
    0.135456225206845, 0.144817696000204, 0.154690314264015, 
    0.163929339640691, 0.173320849343968, 0.182897067780304, 
    0.192446457928478, 0.201450877772469, 0.211165453390326, 
    0.220272349681062, 0.229868712784769, 0.239548389049971, 
    0.248827529155052, 0.258194208131516, 0.267845177286668, 
    0.277503581141909, 0.286725539805162, 0.296137545705906, 
    0.305637298929859, 0.315571105185053, 0.324931704371669, 
    0.33493369164333, 0.344048667157934, 0.353696865199199, 
    0.363190516677303, 0.373009699248996, 0.38232714221291, 
    0.392236897809132, 0.401904950651255, 0.411525147802969, 
    0.42108892685294, 0.43121577086313, 0.440389608588148, 0.450406531358912, 
    0.460487946072634, 0.470253497655302, 0.479728518885724, 
    0.489416712360443, 0.499351918912441, 0.509032269559411, 
    0.519064082539528, 0.529108488864014, 0.539084343279124, 
    0.548722715060096, 0.558845528891268, 0.568749082182345, 
    0.57855218017893, 0.588732758007412, 0.598721275401343, 
    0.608888127039066, 0.61910156277725, 0.629252916507176, 
    0.639381887537984, 0.649501164379409, 0.659892979330005, 
    0.669878817958717, 0.68033118650808, 0.690650771933587, 
    0.700901862330302, 0.71129595427997, 0.721539252149015, 
    0.732054832110591, 0.742580896819032, 0.753031205834931, 
    0.763581737943524, 0.7741349988916, 0.784735311805191, 0.795282611758814, 
    0.806137757950131, 0.816763148935367, 0.827539881959857, 
    0.838298535720483, 0.849208755808617, 0.860044399530641, 
    0.871035990237025, 0.881928976282313, 0.892916124722219, 
    0.903971704069835, 0.915116712731001, 0.926258683552434, 
    0.937441533237879, 0.948715426066321, 0.960018024940174, 
    0.971363461993029, 0.982780966088085, 0.99425069111322,
  -0.994305839112685, -0.982958705608895, -0.971656902636937, 
    -0.96042589044033, -0.949231334686774, -0.938068023196386, 
    -0.926952125675894, -0.915892636723738, -0.904946522236156, 
    -0.893935886599432, -0.883044217724624, -0.872072785890053, 
    -0.861210519936221, -0.850288856908243, -0.839633288590469, 
    -0.828806087143347, -0.81820206702974, -0.807375983899824, 
    -0.796913415410068, -0.786286114063749, -0.775610292779286, 
    -0.765328440314357, -0.754580134754314, -0.744346186670064, 
    -0.733658648006106, -0.723566629260255, -0.712942156703729, 
    -0.702621889479134, -0.692393743034667, -0.682086296615229, 
    -0.671951391007322, -0.661690062054542, -0.651355557443243, 
    -0.641172322990558, -0.631044808729292, -0.620984263025427, 
    -0.610993441675696, -0.600817926440017, -0.590651497994881, 
    -0.580949596331651, -0.570592092112412, -0.560508825601438, 
    -0.550576888726454, -0.540727035493131, -0.530906830425615, 
    -0.520893573585075, -0.511136581011717, -0.501391435108098, 
    -0.491455454681452, -0.481563300137402, -0.471586536878602, 
    -0.461783870893858, -0.452270206288093, -0.44251263977846, 
    -0.432632250706964, -0.423119235298241, -0.413355181207292, 
    -0.403754569528287, -0.393838199541527, -0.384239853349299, 
    -0.374262067449606, -0.364671009841117, -0.355210502196682, 
    -0.345371378649639, -0.336093089224011, -0.326340563814095, 
    -0.316865840733957, -0.307012967892635, -0.29760440490306, 
    -0.288135827774373, -0.2784992809284, -0.269303992382475, 
    -0.259575897923231, -0.250027063741566, -0.240781473894923, 
    -0.230682239218248, -0.2216817505178, -0.211814993025906, 
    -0.202374241868726, -0.1932209813483, -0.183844700573061, 
    -0.174296856339221, -0.164413560925473, -0.155445071151073, 
    -0.145809906802639, -0.136344366656229, -0.126866652132768, 
    -0.117818896032601, -0.10826375280381, -0.0988197849567091, 
    -0.0892934766415057, -0.0795675804983429, -0.0702986500298178, 
    -0.0608975855507811, -0.0518995637674918, -0.0420966551333911, 
    -0.0326156196903788, -0.0232066778594625, -0.0142377173663334, 
    -0.00471388809754097, 0.00455172882012177, 0.0141003744609063, 
    0.0235090915334673, 0.0328518898911647, 0.0422593588834762, 
    0.0518589071380365, 0.0609859325628226, 0.0706466942725165, 
    0.0799868785484145, 0.0893130591693822, 0.0988196790943402, 
    0.10822015548678, 0.117783381238041, 0.127027973489005, 
    0.136677503329787, 0.145887601441915, 0.15512027435939, 
    0.164531602181096, 0.174104520352917, 0.183794723784359, 
    0.193132741528673, 0.202878987855564, 0.212077151386555, 
    0.221636029909765, 0.230825954300336, 0.240307692794601, 
    0.249910072196502, 0.25959504802375, 0.268921122707413, 0.27854296521733, 
    0.288276466029753, 0.297523854248874, 0.307471590714305, 
    0.316723319318324, 0.326588587244321, 0.335667943589196, 
    0.345287257320676, 0.355110293066117, 0.364752678417146, 
    0.374477459084563, 0.384176467673819, 0.393839184343409, 
    0.403541493349799, 0.413228520100386, 0.422984952765973, 
    0.432706632871183, 0.442155700168733, 0.452038851501253, 
    0.46207722237082, 0.471740472892251, 0.481603938957407, 
    0.491446702524673, 0.501062494181697, 0.511190956381211, 
    0.521139915842187, 0.530849164785934, 0.540818203251949, 
    0.550517225649788, 0.560838655723549, 0.570640048668458, 
    0.580717103147992, 0.5906303335619, 0.600924968597856, 0.610728396495612, 
    0.621029298386893, 0.631058752406834, 0.641133949059946, 
    0.651223308683242, 0.66162071486786, 0.671771943113047, 
    0.681968209759916, 0.692365273673761, 0.702537163276415, 
    0.71308343543755, 0.72327162709901, 0.733741931845686, 0.744095869744908, 
    0.754488774545039, 0.765214707789887, 0.775693016648587, 
    0.786244863630292, 0.796857130891972, 0.807457969122693, 
    0.818225244993133, 0.828791923439271, 0.839619915155039, 
    0.850396278066674, 0.861144955646796, 0.872054892187708, 
    0.882893857688948, 0.893875753257554, 0.904868225407823, 
    0.915820196435544, 0.926956029606823, 0.938045959850794, 
    0.949233266785094, 0.960404307568535, 0.971679594681523, 
    0.982967507518685, 0.994307334347735,
  -0.994364680402046, -0.983117326689602, -0.97191867238597, 
    -0.960732268134912, -0.949666977293364, -0.938545932727415, 
    -0.927507883247026, -0.91655289285252, -0.905632459014091, 
    -0.894685295795353, -0.883755927316026, -0.872975903602821, 
    -0.8622089152559, -0.851481009822746, -0.840671969653473, 
    -0.829959531688647, -0.819347619930551, -0.808865615842081, 
    -0.798106833141089, -0.787448472686084, -0.776956576466535, 
    -0.766604811189194, -0.756176156969963, -0.745788458177586, 
    -0.735207893916594, -0.724950150982796, -0.71462672822686, 
    -0.704211664510269, -0.693996540581925, -0.683682900436693, 
    -0.673298718538706, -0.663287384640967, -0.653054867409584, 
    -0.642837194336622, -0.632575963326351, -0.622630782928022, 
    -0.612545213522075, -0.60224969332122, -0.592082908593462, 
    -0.582410330585684, -0.572186953457134, -0.562155260797813, 
    -0.552511566424996, -0.542490731404854, -0.532606252005559, 
    -0.52271572477929, -0.512639691338484, -0.502842386729219, 
    -0.492955390338291, -0.482786100814254, -0.473299358028401, 
    -0.463220498371294, -0.453910812125391, -0.443822603649643, 
    -0.434099485388127, -0.423923606808238, -0.414743080638134, 
    -0.404779059912434, -0.394952528635474, -0.38534926072808, 
    -0.375834175302737, -0.366094260947474, -0.356480693831099, 
    -0.347021878661644, -0.337153365940918, -0.327493109061825, 
    -0.318171821206708, -0.308465446655336, -0.298899509766359, 
    -0.289334328518697, -0.27962304264206, -0.269988715954918, 
    -0.260536022066455, -0.250996791607716, -0.241480134416044, 
    -0.231693967899042, -0.222444482459366, -0.212795011742399, 
    -0.202891565836689, -0.193833744795385, -0.184404747272486, 
    -0.17484145939371, -0.165388106119027, -0.155909383661595, 
    -0.146351043388795, -0.136859056146967, -0.127572003918893, 
    -0.118599162375718, -0.108635957995186, -0.0990143750237975, 
    -0.0895094128646067, -0.0803495520831832, -0.0705878868985519, 
    -0.0611866471987474, -0.0521461805060993, -0.0422370465846016, 
    -0.0330638075913751, -0.0233705342116362, -0.0142139713661093, 
    -0.00457073854735093, 0.00470274666977389, 0.0140813353576556, 
    0.0235375224075688, 0.0329033571869713, 0.0423364170927573, 
    0.0517114255347712, 0.0613784429026271, 0.0708711243808705, 
    0.0803106288263332, 0.0899401725414386, 0.0993054259429038, 
    0.108540468208576, 0.117988429116301, 0.127648584984137, 
    0.137040875657756, 0.146507687025067, 0.155855404771257, 0.1655542167077, 
    0.175047119479326, 0.184286694264679, 0.193655969060319, 
    0.203392704402046, 0.212984871612676, 0.222622540845447, 
    0.23176458331499, 0.241399616123401, 0.251080277031265, 
    0.260519159976535, 0.270151736798884, 0.279836843422209, 
    0.288968922093377, 0.29876175496712, 0.308384460955119, 
    0.318133168721632, 0.327343275231316, 0.337446517102511, 
    0.346804497754563, 0.356846756169803, 0.366075227352124, 
    0.375658958587282, 0.385474007431856, 0.394939511759418, 
    0.404805236623876, 0.414597784287392, 0.424445391078911, 
    0.433999539011235, 0.443974718705957, 0.453570440456652, 
    0.463673310590578, 0.473289763494219, 0.483143328900656, 
    0.493000343742639, 0.503004209696365, 0.512734940784773, 
    0.522702378626121, 0.532353719266345, 0.542414453908921, 
    0.552319785336448, 0.562157707163994, 0.572458211175427, 
    0.582333080901978, 0.592321186513531, 0.602371654759042, 
    0.612506941955389, 0.622457366749096, 0.632808424293181, 
    0.642790391532564, 0.652980667524449, 0.663193336479671, 
    0.673483973394137, 0.683641369876409, 0.694106174899777, 
    0.704321862249267, 0.714556231997194, 0.724898133683455, 
    0.735209144688288, 0.745525054723244, 0.756194917635683, 
    0.766683096637199, 0.777052651448146, 0.787694163525445, 
    0.798212567466285, 0.808680599307665, 0.819344433548998, 
    0.830028529330858, 0.840679250153734, 0.851403550143987, 
    0.862252159138758, 0.87286474895185, 0.883837174424747, 
    0.894647509363259, 0.905655237717545, 0.916568802095146, 
    0.927527095030371, 0.938526950814911, 0.949641157941892, 
    0.960755039848537, 0.971910096909946, 0.983095890420401, 0.994350316890369,
  -0.994407436744374, -0.98325011529954, -0.972122386401945, 
    -0.961012526735077, -0.949984383572526, -0.938982703534898, 
    -0.928025154509051, -0.917094119395912, -0.906194438094638, 
    -0.8953459347446, -0.884565340525044, -0.873797170183317, 
    -0.862964298682967, -0.852366198844955, -0.841678158077467, 
    -0.831038916872836, -0.820280330316203, -0.809685655352745, 
    -0.799296024205461, -0.788686546387136, -0.778186432389394, 
    -0.767754688273576, -0.75743180509914, -0.746901626660341, 
    -0.73661015265405, -0.726180474638391, -0.715841082294994, 
    -0.705503132738742, -0.695345936432363, -0.684980929405154, 
    -0.674806729390881, -0.664558732706618, -0.654317299058969, 
    -0.644213007843178, -0.634314841486347, -0.623889883285963, 
    -0.613845202721628, -0.604010816776451, -0.593959712215315, 
    -0.583628551060343, -0.573916980551525, -0.56371358736442, 
    -0.553701203109028, -0.543746771684273, -0.534134075344361, 
    -0.52387321561445, -0.51398246483714, -0.504428567930078, 
    -0.494169171018172, -0.484522421712896, -0.474630162528963, 
    -0.464796535574928, -0.454873635780338, -0.445007386148279, 
    -0.435436367176886, -0.425411813799754, -0.415740900273507, 
    -0.406371269232893, -0.396487327216933, -0.386754723343812, 
    -0.377039054378916, -0.366966436785992, -0.357785826477728, 
    -0.347982362265903, -0.338146804598352, -0.328740503321029, 
    -0.31914951231607, -0.309313791138711, -0.299781890544373, 
    -0.289938552404328, -0.280462473083055, -0.271002206439545, 
    -0.26140009279698, -0.252048818933818, -0.242011285126436, 
    -0.232473021086326, -0.223523860616652, -0.213503458493319, 
    -0.204277413631955, -0.19427747541144, -0.184881154253561, 
    -0.175210150535879, -0.165800491051372, -0.156366473352798, 
    -0.146907041844017, -0.137438461210167, -0.127982412935993, 
    -0.118769748109103, -0.10942198908752, -0.0992899724265214, 
    -0.0898748854183811, -0.08034469599527, -0.0714041829332714, 
    -0.0615562575927597, -0.0519318415327981, -0.0428419903369155, 
    -0.0335195474364665, -0.02367335816633, -0.0146716148190043, 
    -0.00498981953555876, 0.00495961451502233, 0.0138379922596585, 
    0.0236324468195313, 0.0332027097311703, 0.0426708289776069, 
    0.0520575791066205, 0.0616860171177248, 0.0709927930745333, 
    0.0805777247916934, 0.0903969383436003, 0.0994470881085312, 
    0.108853906877234, 0.118474137674815, 0.127637216373333, 
    0.137543759871937, 0.146952980537594, 0.15642685520158, 
    0.166176594887405, 0.175340885664754, 0.185260683135592, 
    0.194585030916316, 0.203825584105423, 0.213722118868547, 
    0.222915682356929, 0.232847803098188, 0.242534806879757, 
    0.251625663948967, 0.261197149958485, 0.271065704752813, 
    0.28102693793268, 0.290237733494129, 0.299649140274335, 
    0.309450537536491, 0.318951378490334, 0.328998337991812, 
    0.338140736734249, 0.348079985257667, 0.357558993569729, 
    0.367239844551856, 0.376875155515488, 0.386770355980144, 
    0.396429923585986, 0.406344786728712, 0.415925536461778, 
    0.42556664615917, 0.435169424181357, 0.444936698026874, 
    0.454830372193596, 0.464629898165025, 0.474525819735045, 
    0.484533956140991, 0.494392528503823, 0.503894628544232, 
    0.514221945001108, 0.523801539744762, 0.533815926162915, 
    0.543688877252336, 0.553874920550398, 0.563807446855903, 
    0.573663879112679, 0.583654058697966, 0.593902745879068, 
    0.603770208129802, 0.613770129426579, 0.624128716543559, 
    0.634163573413295, 0.644208202649233, 0.654485217304036, 
    0.664484979393299, 0.67476735018719, 0.684881391449163, 
    0.695369486388878, 0.705537408861594, 0.716037940196481, 
    0.726172489906692, 0.736440904318839, 0.746944627703474, 
    0.757336603264167, 0.767787809636908, 0.778181586427027, 
    0.788708000422453, 0.79926008608972, 0.809876873518608, 
    0.820398855453275, 0.830910401620645, 0.841593695035248, 
    0.852356430578238, 0.863025348140625, 0.873724089595912, 
    0.884520575857648, 0.895391284646497, 0.906222066195783, 
    0.917144720245836, 0.9280183321056, 0.938988644342562, 0.950019840689921, 
    0.961044783568663, 0.97212537338249, 0.983234246571395, 0.994403379370963,
  -0.994466019313238, -0.983410076209977, -0.972393480695827, 
    -0.961411583460133, -0.950471498580968, -0.939572507800569, 
    -0.928694026027913, -0.917845742967385, -0.907041663864347, 
    -0.89624163264008, -0.885492953174411, -0.874773324491491, 
    -0.864091627212043, -0.853419823793197, -0.842874760936296, 
    -0.832307061415635, -0.821789775895697, -0.811154933433488, 
    -0.800598838650461, -0.790262110619642, -0.779820214210931, 
    -0.769247206092192, -0.758919566761204, -0.748691010433877, 
    -0.738068651602638, -0.727740665444704, -0.717380158230547, 
    -0.707366492319089, -0.697053140482077, -0.686809227488364, 
    -0.676552189934189, -0.666429754209883, -0.656332194199748, 
    -0.646196390444506, -0.635923521061735, -0.626050875009239, 
    -0.615720415373492, -0.605577880267454, -0.595468744380335, 
    -0.585668751524772, -0.575540986477178, -0.565565134961704, 
    -0.555624237281674, -0.545490680023489, -0.535698678760635, 
    -0.525988560984956, -0.515949373144571, -0.506094953359351, 
    -0.49581459427797, -0.486236640084451, -0.476319825064218, 
    -0.466492032152619, -0.456550556118906, -0.446809547655118, 
    -0.437141521512728, -0.427286294134308, -0.417380455211007, 
    -0.407868100059729, -0.39811498523359, -0.388011004391761, 
    -0.378424766108114, -0.368918192645157, -0.359217041697443, 
    -0.349433858897886, -0.339804163167161, -0.329913363477733, 
    -0.320430356903939, -0.310707722584755, -0.301277300696418, 
    -0.291483569733568, -0.281734742159083, -0.272358979148625, 
    -0.262343841811132, -0.25320670516297, -0.243319844918383, 
    -0.23358066080453, -0.224035537797862, -0.214384514736058, 
    -0.204785354913466, -0.195220434875784, -0.185723491160325, 
    -0.176266858540527, -0.166428051764292, -0.157367456050355, 
    -0.147904614802964, -0.137947449945512, -0.128536885929193, 
    -0.118842788488222, -0.109365457635242, -0.100131246927666, 
    -0.0905047099308258, -0.0808335612700739, -0.0713452915145985, 
    -0.0619069663245469, -0.0522697960859925, -0.0428262792043543, 
    -0.0330380093515606, -0.0236707660883511, -0.0142752193589314, 
    -0.00458574693333493, 0.00486620618866865, 0.0143995104526075, 
    0.023774314685693, 0.0333287142806459, 0.042776135882427, 
    0.052431535502207, 0.0618977600296324, 0.0712656306173698, 
    0.0809880576311441, 0.0905395276615356, 0.0997700950421575, 
    0.109450014866457, 0.119095083847601, 0.128660996813725, 
    0.138067224760419, 0.147651366201825, 0.157247360824856, 
    0.166805638068636, 0.176533378396547, 0.185690556113222, 
    0.195479845853869, 0.20486275033407, 0.214219190051392, 
    0.224086564823227, 0.233370692606838, 0.243344398643161, 
    0.253131150365512, 0.262572875228387, 0.272191516134487, 
    0.281596807842158, 0.291334976440029, 0.301146368381795, 
    0.310820091733844, 0.32020669998293, 0.330299188448136, 
    0.339844788751589, 0.349304439049699, 0.358905770050587, 
    0.368931390461964, 0.378537970074857, 0.388333179775699, 
    0.398050300175008, 0.407772491135242, 0.417697364043331, 
    0.427413645092013, 0.437059407279782, 0.446853361035797, 
    0.456773525757564, 0.466480072480004, 0.476521973270563, 
    0.486186369662033, 0.495949733050623, 0.506043423452427, 
    0.515842895373304, 0.525701517091193, 0.535790420308158, 
    0.545811034885819, 0.5555493809124, 0.565440864097718, 0.575681415127978, 
    0.585455444602198, 0.595595786914679, 0.605678938246409, 
    0.615677844835639, 0.6259021152924, 0.635931731824654, 0.645726281196817, 
    0.656375687035627, 0.666418470614718, 0.676737916413713, 
    0.686831222569219, 0.697188948636243, 0.707371429333097, 
    0.717518329176499, 0.727796298736497, 0.738127127652419, 
    0.748517990069279, 0.758759673810933, 0.769347550451823, 
    0.779692487076505, 0.790179467540708, 0.800756363384154, 
    0.811130034913706, 0.821652489498252, 0.832213659342447, 
    0.842857053048436, 0.853505033465127, 0.864109835252252, 
    0.874790915086665, 0.885513344816247, 0.896178526478118, 
    0.90702817996463, 0.917837175573193, 0.928708233143012, 
    0.939521272296887, 0.950458972644727, 0.9613962535629, 0.972375979882271, 
    0.98340669680311, 0.99445802765831,
  -0.994480034978883, -0.983452783797433, -0.972472543238291, 
    -0.961516948543938, -0.950599249355848, -0.939731162761756, 
    -0.928851583203956, -0.918023436552532, -0.907294916432091, 
    -0.896559113812576, -0.88581252936377, -0.875035322527193, 
    -0.864416123310209, -0.853879670224784, -0.843186168833968, 
    -0.832644820690152, -0.82212117371491, -0.811626254187264, 
    -0.801081446657361, -0.790600166951834, -0.78019034585487, 
    -0.769789695673819, -0.759373002890819, -0.748964015057731, 
    -0.738540908622551, -0.728392463139468, -0.717983032396764, 
    -0.707780234210086, -0.697569771885205, -0.687251059770956, 
    -0.67711267901497, -0.666828823403474, -0.656677867058341, 
    -0.646595404083327, -0.636615237809018, -0.626334143630178, 
    -0.61628225685352, -0.606210860098601, -0.596151654125968, 
    -0.586065317136322, -0.576180556717852, -0.566057901596181, 
    -0.556306387172121, -0.546010856527102, -0.536451757854637, 
    -0.526532556479619, -0.516315757327428, -0.506269705843812, 
    -0.496467368917015, -0.486648701435053, -0.476939766574801, 
    -0.466915162878629, -0.457024081565697, -0.447277503084294, 
    -0.437567404131141, -0.427841238699922, -0.418165929144913, 
    -0.408080363238764, -0.398642069780699, -0.388745172611843, 
    -0.378985061942102, -0.369498393266131, -0.359603726054083, 
    -0.349806764439897, -0.340175227536085, -0.330412713513818, 
    -0.320241510876172, -0.310866293491593, -0.301438008515207, 
    -0.291738797921608, -0.282120181777834, -0.272705270294788, 
    -0.26295386983794, -0.253169153119044, -0.243641519389026, 
    -0.234036144223721, -0.224496552005399, -0.214994979640935, 
    -0.205277459363372, -0.195622022352147, -0.185877794361994, 
    -0.176409751765809, -0.166735444602603, -0.157327151715824, 
    -0.147718577418741, -0.138466315570481, -0.128800965127588, 
    -0.11904986910198, -0.109935575869281, -0.0999094194409271, 
    -0.0907756676182827, -0.0810171731782913, -0.0710937561715044, 
    -0.0618923861984281, -0.0524771802273781, -0.0429619163362962, 
    -0.0335599996093589, -0.0237145083185169, -0.013901611721891, 
    -0.00442728241027656, 0.00456936913708036, 0.0145464680376151, 
    0.0239331313774852, 0.0334748776251078, 0.0431167494411597, 
    0.052491030726164, 0.0618169989949861, 0.0714137490024067, 
    0.0810073869574476, 0.0906499980527674, 0.0998734891205858, 
    0.109632158320766, 0.118930964287106, 0.128831335871975, 
    0.137972953045173, 0.147952607845961, 0.157342510616793, 
    0.166749950369861, 0.176403416146307, 0.186020498713535, 
    0.195678230199876, 0.205180653313998, 0.214659461183409, 
    0.224662390551199, 0.23406424568851, 0.244032027221444, 
    0.253309797208892, 0.262888836768003, 0.272691416024045, 
    0.282187384590827, 0.291693767894376, 0.301460832715214, 
    0.311402503343036, 0.320790658312171, 0.330366197610741, 
    0.340242014134369, 0.349519875313863, 0.35967482351958, 
    0.369520447941889, 0.378887918613608, 0.388608271553843, 
    0.398264843548436, 0.40784958151066, 0.417969774837726, 
    0.427766763543976, 0.437585252893276, 0.447434201013532, 
    0.457108365352325, 0.466974969551316, 0.476864092364184, 
    0.486811777495822, 0.496695175109519, 0.506454420262842, 
    0.516308609230485, 0.526103883002517, 0.536113343818331, 
    0.546314375668149, 0.556103870116636, 0.566113648068019, 
    0.576129645925575, 0.586282935321775, 0.596140659783287, 
    0.606122284745005, 0.616231600859537, 0.626225689893182, 
    0.636581962785948, 0.646710000027993, 0.656758645202076, 
    0.66694218775038, 0.677121808183279, 0.687287268788672, 
    0.697476227248902, 0.707821045118254, 0.718017296115215, 
    0.728503248043337, 0.738603469930445, 0.749046654061583, 
    0.759263545012773, 0.769704518346619, 0.780192302832024, 
    0.790528310421542, 0.801100842834881, 0.811578007574024, 
    0.822121884736137, 0.832522749455426, 0.843222029182135, 
    0.853824489184209, 0.864453997341378, 0.87509774864635, 0.88583684517574, 
    0.896491428076463, 0.907197887075165, 0.918037168295424, 
    0.928884187145115, 0.939699494239607, 0.950604021340674, 
    0.961514803613852, 0.972462787879153, 0.983450159173136, 0.994474519463263,
  -0.994531851440943, -0.983613921746897, -0.972731129281934, 
    -0.961869961551452, -0.951086075744997, -0.940262383605067, 
    -0.929499602644797, -0.918751984575371, -0.90809649731512, 
    -0.897393693157155, -0.88678661728335, -0.876161969569044, 
    -0.865530820661012, -0.854968439303116, -0.844446442024205, 
    -0.833963790024296, -0.823450841918895, -0.812925959809827, 
    -0.802443001960733, -0.792175791274813, -0.781687074729336, 
    -0.771347932487976, -0.760973715480531, -0.750709669602932, 
    -0.740419875752255, -0.729942045671794, -0.719609501440866, 
    -0.709403853220231, -0.699364515144566, -0.689211796086513, 
    -0.678952259554508, -0.668809022743158, -0.658694944871837, 
    -0.648538018482495, -0.638359243863189, -0.628360212953284, 
    -0.618246564409799, -0.608242675058243, -0.598197337018961, 
    -0.588041514134539, -0.578091698160526, -0.567946599521535, 
    -0.558253518452927, -0.548093625687523, -0.538092816617885, 
    -0.528134434999739, -0.518219506109161, -0.508398897118043, 
    -0.498483607740128, -0.488571647691999, -0.478646591051922, 
    -0.468811691258851, -0.458889809253395, -0.449298027600624, 
    -0.439164904321893, -0.429523718101111, -0.419612461164051, 
    -0.409856999963703, -0.400000960082614, -0.390392264757826, 
    -0.380547293416975, -0.370775714357587, -0.360966400436606, 
    -0.3512825824857, -0.341761838060289, -0.331718349988391, 
    -0.322040983133709, -0.312598794578818, -0.302893475883547, 
    -0.293048948103879, -0.283238127264622, -0.273881998582161, 
    -0.264118859731348, -0.25437501085034, -0.244771988718103, 
    -0.234610091241904, -0.225534629812283, -0.215686876220673, 
    -0.206051605425623, -0.196695312009842, -0.187183670680614, 
    -0.177469845613394, -0.167846169867814, -0.158089578596042, 
    -0.148336093485777, -0.138761690732433, -0.129423026117575, 
    -0.119852542562713, -0.110232911464034, -0.100348993948638, 
    -0.0910300725607176, -0.0813887590009382, -0.0718285451667314, 
    -0.0622830809758558, -0.0526704606424595, -0.0430006121311525, 
    -0.033498240100882, -0.0240182374908857, -0.0144697929504149, 
    -0.00508162976917849, 0.00475252530816062, 0.0145387067629353, 
    0.0240483811584262, 0.0334536522306038, 0.0431518552466235, 
    0.0525885910798413, 0.0623269944632693, 0.0719962141199413, 
    0.0813208982884772, 0.0911568407042454, 0.100508146120773, 
    0.110072507829324, 0.119432531672875, 0.129103780533194, 
    0.138967316249163, 0.148418872991588, 0.158147512316111, 
    0.167589923492311, 0.177377530439784, 0.187272854444484, 
    0.196695692303841, 0.206254811655886, 0.216024825921593, 
    0.225317015562252, 0.234807126167613, 0.244668539180018, 
    0.25420198818494, 0.264050834989918, 0.274055511511734, 
    0.283325413498274, 0.293241736846745, 0.302813576267216, 
    0.312300085861157, 0.322189254487504, 0.331836477035877, 
    0.341629753725386, 0.351454306086864, 0.361004507554137, 
    0.370926310449262, 0.380553322150184, 0.390355157906727, 
    0.399913871044144, 0.409965346839522, 0.419918011766261, 
    0.429219058391919, 0.439224794192811, 0.449299440960122, 
    0.459206539138731, 0.468795358285428, 0.478849261860805, 
    0.488791364003937, 0.498385412550705, 0.508208028137217, 
    0.518227526389844, 0.528105997981328, 0.538135596655139, 
    0.548189495690209, 0.557994086264177, 0.567958087816533, 
    0.578177902882295, 0.587795364015275, 0.598185451679348, 
    0.608017594241406, 0.61821895326881, 0.628154771116842, 
    0.638335267116123, 0.648543947017187, 0.658668760299666, 
    0.668753641824237, 0.67893294595843, 0.689058173469273, 
    0.699398391404354, 0.709478416701371, 0.719764218082125, 
    0.730112322791859, 0.740362514710419, 0.750733131967076, 
    0.761013559448989, 0.771380512938029, 0.781629634424384, 
    0.792168066163237, 0.802486370640223, 0.812967828777382, 
    0.823416087846534, 0.834001060208744, 0.844364206181341, 
    0.854931064312527, 0.865617148188412, 0.876211852671859, 
    0.886760715713296, 0.897434020957511, 0.908091629767438, 
    0.918807402336778, 0.929510987094881, 0.940265986831271, 
    0.951072847632997, 0.961882111496181, 0.972731095435741, 
    0.983622953546275, 0.994532546651181,
  -0.994558391228747, -0.983688622239569, -0.972850764472399, 
    -0.962048035085906, -0.95128227292376, -0.940518215651286, 
    -0.929759609010524, -0.919127316407889, -0.908466567366888, 
    -0.897775997748252, -0.887142501040449, -0.876572122336935, 
    -0.866015396466161, -0.855538474299032, -0.844964846433042, 
    -0.834530486300615, -0.824001955945632, -0.813478459890231, 
    -0.803231665572084, -0.792794864926225, -0.782240975560438, 
    -0.772029997674731, -0.761667832536963, -0.751298942775411, 
    -0.741141911714583, -0.730669381710767, -0.7205604796158, 
    -0.710175886967347, -0.700115812168683, -0.689883388999323, 
    -0.67991759899747, -0.669584100877038, -0.659359189126819, 
    -0.649314770088608, -0.639073377439905, -0.629002631423765, 
    -0.619010474454915, -0.608969705699232, -0.598742509548363, 
    -0.588789765307732, -0.57892956814859, -0.568936469585832, 
    -0.558797500218881, -0.548709084129831, -0.53892912454548, 
    -0.529014599478837, -0.519060075307134, -0.509077197807577, 
    -0.499215751951437, -0.489247987195908, -0.479411186280667, 
    -0.469678444130185, -0.459726187364635, -0.449578757713991, 
    -0.44015258699711, -0.430384522395253, -0.420610913786875, 
    -0.410578430593476, -0.4006640122286, -0.391064590314468, 
    -0.381232312227378, -0.371342386666818, -0.361933636765222, 
    -0.352072611523622, -0.342478909678899, -0.332376441570625, 
    -0.322760124135825, -0.313278084842315, -0.303386108708069, 
    -0.293401931612347, -0.283947524677819, -0.274607053180351, 
    -0.264675802372765, -0.254923798164295, -0.245370251515057, 
    -0.235549776081422, -0.225691416934281, -0.216286473418995, 
    -0.206734049671917, -0.196784137980226, -0.187617219824828, 
    -0.177318352632728, -0.168037506886237, -0.158514969575002, 
    -0.148856002023445, -0.139300562469302, -0.129500375128866, 
    -0.119822458322472, -0.110339006663293, -0.100664225232907, 
    -0.0911256732338305, -0.0814269542205042, -0.0718951744930996, 
    -0.0623676421026188, -0.0527839902153731, -0.0431757580610727, 
    -0.0333993340032678, -0.0240928605712367, -0.0143415025077004, 
    -0.00508258992366757, 0.00471992817137372, 0.0143373089903147, 
    0.0241678015272247, 0.0336786721416975, 0.0430737717196158, 
    0.0526678214443833, 0.0623719601407372, 0.0720764430646051, 
    0.0815722052067265, 0.0910983584009677, 0.100965608095743, 
    0.110436017141045, 0.120143505914268, 0.129781746859177, 
    0.139266643091424, 0.148771065916963, 0.158385303617465, 
    0.167900498892362, 0.177709852742384, 0.187355761192658, 
    0.19719907835586, 0.206006331858904, 0.216388846570762, 
    0.225890777336468, 0.235185505521869, 0.245109909071846, 
    0.255403568988427, 0.264702916214629, 0.274490355661018, 
    0.284114062366585, 0.293567654066405, 0.303494022401672, 
    0.312915820905486, 0.322558727934078, 0.33249748905164, 
    0.342348833140752, 0.351939210511517, 0.361498818217263, 
    0.371400263380001, 0.381090702207239, 0.390934826373871, 
    0.400765833589215, 0.410700899197232, 0.420308942493772, 
    0.43022975596423, 0.440150484472352, 0.449907240184359, 
    0.459691072207308, 0.469657314266021, 0.479419083104638, 
    0.489133453662698, 0.499178873116005, 0.508787642644581, 
    0.518982939427584, 0.529078402393345, 0.53903957752295, 
    0.548936439472971, 0.558906526071693, 0.568730619849451, 
    0.578806027563778, 0.588867247704894, 0.598853362221121, 
    0.609187847031824, 0.619041255938352, 0.629060306258793, 
    0.639108090849503, 0.649314241436906, 0.659374603206223, 
    0.669516599340165, 0.679781108666135, 0.689793383073288, 
    0.700098587862125, 0.71034767206533, 0.720360900030066, 
    0.730824010499799, 0.74110572242554, 0.751347126514798, 
    0.761594080446338, 0.772059601218818, 0.782283547660682, 0.7928086020021, 
    0.803154692860209, 0.813628672729369, 0.823953309746155, 
    0.834510237600865, 0.844999428621846, 0.855527720494038, 
    0.865943913956869, 0.876595002105721, 0.887173162254921, 
    0.897770430442691, 0.908443008799926, 0.919084561428488, 
    0.929785415599211, 0.940510960187125, 0.951268365683368, 
    0.962053086125389, 0.972855051340467, 0.983689170290896, 0.994560267809094,
  -0.994579013778687, -0.983755288873741, -0.972957789198039, 
    -0.962184303624715, -0.951432643026565, -0.940736765189836, 
    -0.930086022175229, -0.919391900192408, -0.908721372904366, 
    -0.898129215180948, -0.887550764269506, -0.877019998557414, 
    -0.86651019491997, -0.855884005075258, -0.845477000015255, 
    -0.834912715079584, -0.824494071035524, -0.814028674132261, 
    -0.803809972219732, -0.793300087824428, -0.782947767060978, 
    -0.77259079405976, -0.762250305407208, -0.751948898571638, 
    -0.741770430645883, -0.731425748560384, -0.721168279498546, 
    -0.711009654380987, -0.700644827227157, -0.690562067091893, 
    -0.680371630669465, -0.670203004989096, -0.660069763168263, 
    -0.649955490899368, -0.639884527188594, -0.629839883976876, 
    -0.619694123657662, -0.609560170312059, -0.599605625339615, 
    -0.589502554906482, -0.579588988799567, -0.56957417884928, 
    -0.559625182008307, -0.54972073880947, -0.53965359995479, 
    -0.52985197982226, -0.519783493236377, -0.509878055991532, 
    -0.500136391970819, -0.490039615909855, -0.480320543478217, 
    -0.47032260392313, -0.460405934561483, -0.450679208451863, 
    -0.440735449580055, -0.431124482121724, -0.421253848132425, 
    -0.411189210009097, -0.401507816263075, -0.391727137347153, 
    -0.381928901395115, -0.372047643840677, -0.362128139207754, 
    -0.352619274220761, -0.342574326691529, -0.332900609849984, 
    -0.323120027563055, -0.313505294632844, -0.303942277993853, 
    -0.293884886126277, -0.284670559899482, -0.274971513626484, 
    -0.265114980293747, -0.255098625768988, -0.245936698258298, 
    -0.235830300127986, -0.226337484361444, -0.216732069534103, 
    -0.207179591352739, -0.19716268736253, -0.187826078875998, 
    -0.178015431221987, -0.168245497130425, -0.158738185250737, 
    -0.1491803355716, -0.139550072862651, -0.130065747442632, 
    -0.120214683804295, -0.110576546413938, -0.101070121238912, 
    -0.0912233589333799, -0.081909961299411, -0.0720907252188298, 
    -0.0625563264456831, -0.0527047042235438, -0.0433361515228231, 
    -0.0336300433185205, -0.0238763834976608, -0.0142522064758843, 
    -0.00466825521305901, 0.0050024440456141, 0.0145056050170416, 
    0.0241638984970743, 0.0335200485238123, 0.0431565645349308, 
    0.052951805190073, 0.0625803313547142, 0.0719271907742564, 
    0.0815340884415484, 0.0912925660630688, 0.10134321161062, 
    0.110493090196394, 0.120020008263369, 0.129920974170994, 
    0.139550129956595, 0.149113432951177, 0.158780432385558, 
    0.168369203484087, 0.178017251141553, 0.187807174083646, 
    0.197506876547423, 0.207031043081108, 0.216796999949823, 
    0.226467331991486, 0.236142750983126, 0.245795410032246, 
    0.25535422904111, 0.264922476298161, 0.274696047558529, 
    0.284338194988238, 0.294175548985312, 0.303967718442632, 
    0.313498396236428, 0.323490739206006, 0.333217437936555, 
    0.342646081965798, 0.352469901146952, 0.362367891027181, 
    0.372087433020222, 0.381906735402571, 0.391636904721614, 
    0.401284472790834, 0.41130393277158, 0.421001537087913, 
    0.430877114683263, 0.440621814590152, 0.450680261156974, 
    0.460385094145965, 0.470294884781978, 0.480191932327918, 
    0.490000840617523, 0.499863970594604, 0.509807915111486, 
    0.519701238792646, 0.529805728005007, 0.539742036615498, 
    0.549620424749594, 0.559642704808723, 0.569640880391429, 
    0.579562584298681, 0.589429101839449, 0.599710328203515, 
    0.60988677554319, 0.619665162110599, 0.629733503052943, 
    0.639839849937806, 0.649996180770997, 0.66023263659287, 0.67017948469015, 
    0.680468029520617, 0.690569959856107, 0.700652255576128, 
    0.710935652552839, 0.721280181039229, 0.73142868051612, 
    0.741694954594678, 0.751962042370301, 0.762347718983361, 
    0.772637107055159, 0.782898555910541, 0.793362860936482, 
    0.803732930468295, 0.814092911061553, 0.824528281688547, 
    0.834971406322015, 0.845439426662945, 0.855925017412249, 
    0.866368679336969, 0.87698284839772, 0.887549067966017, 
    0.898114059794444, 0.908712364033837, 0.919424970154818, 
    0.930045773691323, 0.94070643618097, 0.951441016556097, 
    0.962193855577997, 0.972964060150581, 0.983766878005189, 0.994584136879682,
  -0.994593410725575, -0.983791925855685, -0.972999763752363, 
    -0.962283460787516, -0.95152002581735, -0.940848824170802, 
    -0.930167390730054, -0.919526487998647, -0.908877173822184, 
    -0.89831385249568, -0.887732003897668, -0.877146873484995, 
    -0.8667476783545, -0.856083545251036, -0.8455468714122, 
    -0.835191694964816, -0.824763619097987, -0.81426726129587, 
    -0.804024581587764, -0.793510402625898, -0.783259857135759, 
    -0.772961944594139, -0.762666772051677, -0.752297526029959, 
    -0.74208265104521, -0.7317930673175, -0.72156230152762, 
    -0.711287618058132, -0.701145000618623, -0.691011744212515, 
    -0.68061066277808, -0.670602678248564, -0.660488912535918, 
    -0.650298400622273, -0.640312123713359, -0.630302457730933, 
    -0.620019439851422, -0.610227523372811, -0.600003677075864, 
    -0.589901691475478, -0.579981140083945, -0.569858256042113, 
    -0.559726368770357, -0.549661175529781, -0.539911910539427, 
    -0.529909336760353, -0.519997816351499, -0.510304803610555, 
    -0.500264936444775, -0.490229044278493, -0.480524615925011, 
    -0.470702633375305, -0.460798209198135, -0.450867674852088, 
    -0.441082818403269, -0.430967801117192, -0.421390744344343, 
    -0.411522243402831, -0.401760319494164, -0.392020439988993, 
    -0.382083788766151, -0.372546176329965, -0.362473449670845, 
    -0.35294487204846, -0.342846977723807, -0.333282705109883, 
    -0.323701503414297, -0.313905852161618, -0.304088290421227, 
    -0.294288203901563, -0.284487519468528, -0.274806972038387, 
    -0.265330729409586, -0.25563156045023, -0.245902737306279, 
    -0.236410041242564, -0.2264392569736, -0.217028401700817, 
    -0.207199990952376, -0.197716388463607, -0.187920869340414, 
    -0.178227607090697, -0.168626189860518, -0.159004365748095, 
    -0.149435341958052, -0.139886611334799, -0.130080210563042, 
    -0.120163358344779, -0.110652084640023, -0.101175546634951, 
    -0.091397731195707, -0.0818344766861801, -0.072108916903213, 
    -0.0625831259630572, -0.0529636208864684, -0.0432894255203167, 
    -0.0336908787502299, -0.0241576140391728, -0.0143935690641361, 
    -0.00496278251710957, 0.00463568637867463, 0.014576954902202, 
    0.0241336979427148, 0.0336292117679221, 0.0434018653363169, 
    0.0529811915267713, 0.0624553215779554, 0.0722931341497467, 
    0.0815604620147247, 0.0913084835572827, 0.100810281065356, 
    0.110915848428428, 0.120295457101141, 0.130074162849313, 
    0.139772862826409, 0.149348183739421, 0.158651322672294, 
    0.168407360599126, 0.178125652386328, 0.187760504456071, 
    0.197369401062981, 0.207031732800284, 0.216743595822552, 
    0.226373775211998, 0.236135368676421, 0.245906828334194, 
    0.255634698700429, 0.265354466343213, 0.275109578537446, 
    0.284601133691254, 0.294495193987244, 0.304043349413569, 
    0.313900647424301, 0.323241947463576, 0.333113851327501, 
    0.343091270301952, 0.352689606462916, 0.362623322642785, 
    0.372298014938054, 0.382151980626208, 0.391909824896955, 
    0.401643290728378, 0.411538997491114, 0.421283362173451, 
    0.431322715411889, 0.441092146039668, 0.451182929261676, 
    0.460798621028222, 0.470597137344542, 0.48041687482054, 
    0.490317956999933, 0.500356376760483, 0.510074191529382, 
    0.520016457350536, 0.530093766524316, 0.540080858011887, 
    0.549924465851974, 0.55996125497757, 0.56996813321959, 0.580047277613255, 
    0.590031203934125, 0.600231561020259, 0.609927322782481, 0.6201314191003, 
    0.630169459616487, 0.640186511081181, 0.650317654399966, 
    0.660441654793893, 0.670679513944458, 0.680771602145024, 
    0.690982894766102, 0.701112282082251, 0.711348735383323, 
    0.721502847288472, 0.73179594536172, 0.741955348243902, 
    0.752307996115825, 0.762631371060666, 0.772921826063078, 
    0.783257776725765, 0.793529744877309, 0.80396639595794, 
    0.814389713269203, 0.824793350285289, 0.835242514743884, 
    0.84564347710873, 0.856108962436743, 0.866619477463372, 
    0.877159299407191, 0.887729441601086, 0.898311557236544, 
    0.908860610652394, 0.919517628321829, 0.930176004480367, 
    0.940828452859985, 0.95154744225901, 0.96224338922006, 0.973001902200766, 
    0.983787659797746, 0.994592034736824,
  -0.994611194199906, -0.983861938532704, -0.97313277803233, 
    -0.96244213702908, -0.951744120994893, -0.941109959114978, 
    -0.930462147749416, -0.91985460013942, -0.909287071048147, 
    -0.898718017270393, -0.888162631140203, -0.877615069088468, 
    -0.867205703222449, -0.856695942896003, -0.846330996209286, 
    -0.835819278124341, -0.825418826502104, -0.815089818019841, 
    -0.804685560485883, -0.794278586083882, -0.783889713201306, 
    -0.773747493579174, -0.763384291833111, -0.753024646177393, 
    -0.742863116136273, -0.732606562191878, -0.722376359869209, 
    -0.712181286704747, -0.702075830106827, -0.691657561104404, 
    -0.681550612397475, -0.671557175553214, -0.661280651599086, 
    -0.65139702626043, -0.64109872084836, -0.631234974068325, 
    -0.620986274787526, -0.610920964223647, -0.600903282546888, 
    -0.590876841849647, -0.58093802679167, -0.570869891261899, 
    -0.560838039356799, -0.550943504345255, -0.540974031966135, 
    -0.530954668856732, -0.52090216178747, -0.51111881233164, 
    -0.501127666756368, -0.491283032066558, -0.481429016525638, 
    -0.471450920865687, -0.461420371707365, -0.451976050740438, 
    -0.441745914206877, -0.431965547904293, -0.422216966114857, 
    -0.412362972397372, -0.402429036228457, -0.392783019121478, 
    -0.383118448976554, -0.372936949118777, -0.363218538856444, 
    -0.353475877990739, -0.343751432859864, -0.334098349834937, 
    -0.324294166975361, -0.314482271648991, -0.304834153634075, 
    -0.295030231352142, -0.285331768101836, -0.275627946188552, 
    -0.265795208378644, -0.256207611252105, -0.246480156892289, 
    -0.23672095705312, -0.227183828635757, -0.217449440498111, 
    -0.207472634740823, -0.197888267876184, -0.188030482061383, 
    -0.178658298438443, -0.169029881695178, -0.159110766860445, 
    -0.149691097397294, -0.139951040522784, -0.13022726644425, 
    -0.120551234410099, -0.110826895866068, -0.101256199260584, 
    -0.0916080595649317, -0.0822296354079936, -0.0724511220844237, 
    -0.0629502056800617, -0.0529563792544004, -0.0431061496832589, 
    -0.0337288256096337, -0.0241127411387142, -0.0145678845740229, 
    -0.00497554539224609, 0.00472345005715194, 0.014574569759672, 
    0.0238203823455291, 0.0338575391146014, 0.043382268541482, 
    0.0529344037095982, 0.0627366952803713, 0.0719467982046649, 
    0.0820798145628585, 0.0911839125247817, 0.101296210974764, 
    0.111011828186408, 0.120645705667196, 0.130449800638771, 
    0.140037891893438, 0.149620481675946, 0.159024767672162, 
    0.168729576897435, 0.178560206425032, 0.188191561020943, 
    0.198010914500896, 0.20792298790499, 0.217408617053162, 
    0.226856788576233, 0.236575100274649, 0.246168287660288, 
    0.256316886811816, 0.265904286945388, 0.275299496066948, 
    0.285326979959389, 0.2953098065812, 0.304809687588456, 0.31451118547019, 
    0.324369082131604, 0.333870633250153, 0.344066202616154, 
    0.353684809457679, 0.363387329513461, 0.373173538777676, 
    0.382914688054815, 0.392839093472067, 0.402447466691816, 
    0.412363127909256, 0.422202431589211, 0.432296754714946, 
    0.441790358694112, 0.451894892502634, 0.461718361256747, 
    0.47124069380612, 0.481405468943892, 0.491222670572569, 0.50116519988153, 
    0.511233171655961, 0.521026408742662, 0.531037316237017, 
    0.54075463172786, 0.550990113058526, 0.560877560395834, 0.57088515798064, 
    0.580958812768567, 0.590864127964338, 0.600968360033114, 
    0.610744192530868, 0.621106987808908, 0.631021103723165, 
    0.641138764037088, 0.651262601272468, 0.66141198095542, 
    0.671542263329952, 0.681631113785438, 0.691793281293661, 
    0.701988333303315, 0.712234235942102, 0.722430486987598, 
    0.732603999349727, 0.742816469014515, 0.753167447643859, 
    0.763362234230811, 0.773596231634574, 0.784011896204445, 
    0.794326682376295, 0.804645396110392, 0.815051301684792, 
    0.825495095586229, 0.835756530272936, 0.846181202967219, 
    0.856633086864829, 0.867148536933042, 0.877704605887489, 
    0.888168745028819, 0.898760926135409, 0.909318267982125, 
    0.919856748068425, 0.930468582515188, 0.94111355401332, 
    0.951764573193508, 0.962444072823493, 0.973141860065256, 
    0.983864956285232, 0.994616833054946,
  -0.994630447771906, -0.983908831598932, -0.973192893577807, 
    -0.962544984415862, -0.951899252858313, -0.941263764623101, 
    -0.930685087505012, -0.920098851915375, -0.909545609492572, 
    -0.899015717695306, -0.888495010712619, -0.877976481661964, 
    -0.867506879921691, -0.857071962578833, -0.846585280020835, 
    -0.836280018882649, -0.825852511992366, -0.815456877275198, 
    -0.805120247845036, -0.79480445888243, -0.784441183826221, 
    -0.774122963880943, -0.763840651842496, -0.753591616351881, 
    -0.743351492467123, -0.7331369428473, -0.722867538258399, 
    -0.712650750214143, -0.702476124135712, -0.692307006429233, 
    -0.682178393600063, -0.671995299842321, -0.661941850820899, 
    -0.65188519558472, -0.641800729615405, -0.631527493113216, 
    -0.621615302284355, -0.611560904361057, -0.601618428093889, 
    -0.59140068354237, -0.58145133807292, -0.571431824983418, 
    -0.561501369582247, -0.551377297778809, -0.541461360844406, 
    -0.531446405220201, -0.521516172079862, -0.511682509915034, 
    -0.501740760129987, -0.491885289786571, -0.481953973561926, 
    -0.472314738715556, -0.462178690560017, -0.452197351344514, 
    -0.442356369462184, -0.432897678336708, -0.422879215813403, 
    -0.413073424508736, -0.403027652794831, -0.393193714097362, 
    -0.383545682441575, -0.373703122341274, -0.363936187315382, 
    -0.353903458873899, -0.344137202526677, -0.334394349091801, 
    -0.324507252057428, -0.314856555851602, -0.305338434685608, 
    -0.295526968948871, -0.285842120753657, -0.275897870460225, 
    -0.266343371625811, -0.256453022884992, -0.246785317046487, 
    -0.237317557535563, -0.227512940226758, -0.217557058471183, 
    -0.207825399552088, -0.198347402071597, -0.188522961519688, 
    -0.178915663703617, -0.169319192988678, -0.159711063199013, 
    -0.149869350927937, -0.140254959206891, -0.130404871323972, 
    -0.120826916847988, -0.110996538047167, -0.101390142124612, 
    -0.091726390397148, -0.0821656362201286, -0.0724794163394961, 
    -0.0628455675559594, -0.0534695221116148, -0.0433809668416659, 
    -0.0341474729429223, -0.0242705380535561, -0.014638141021502, 
    -0.0047682452127018, 0.00478510177816319, 0.0143295451312918, 
    0.0243537538591658, 0.0339992039808094, 0.0435284408288746, 
    0.0527681823668157, 0.0627185142319357, 0.0722467291184104, 
    0.0822007849430604, 0.0915071359249108, 0.10164784088119, 
    0.111190367274627, 0.120663131842887, 0.130355367073986, 
    0.140045178453063, 0.149815555718921, 0.159307427227459, 
    0.169027166620309, 0.178984717324809, 0.18854166540463, 
    0.198173773696768, 0.207817168799194, 0.21759150323443, 
    0.227304196663352, 0.237001701258839, 0.246779712601487, 
    0.256524764627223, 0.266315724573145, 0.276081796601457, 
    0.285478975990393, 0.295469286554171, 0.304927678472806, 
    0.315076287785152, 0.324996795091321, 0.33451196819327, 
    0.344399569286142, 0.35407880583325, 0.363739413237167, 
    0.373792149514071, 0.383391017935098, 0.393107662956724, 
    0.403051855514709, 0.412783916736622, 0.422816040315614, 
    0.432662747601775, 0.442230298429167, 0.452441772990355, 
    0.462099686826837, 0.471967722916787, 0.481968405299332, 
    0.491698054935417, 0.501581129902273, 0.511629194837667, 
    0.52164055940057, 0.531437988158109, 0.541482084906051, 
    0.551498350689441, 0.561421794718424, 0.571553790577492, 
    0.581426698296793, 0.591310585508828, 0.60148907811235, 
    0.611633735973412, 0.621506167206922, 0.63163762344916, 
    0.641717961649346, 0.651839338099346, 0.661955331793134, 
    0.672083673808706, 0.682197099250142, 0.692253578564968, 
    0.702380436113222, 0.712685209937035, 0.722813793761346, 
    0.733066066795659, 0.743339282368636, 0.753611475433157, 
    0.763835841574423, 0.774123771496251, 0.784392660612702, 
    0.794743265510035, 0.805088393123016, 0.815447576171137, 
    0.825862971622556, 0.836210588457692, 0.846672381207727, 
    0.857041437940187, 0.867468708048689, 0.878005312162417, 
    0.888488501309798, 0.899013842571442, 0.909508477415027, 
    0.920114651301483, 0.930671820618466, 0.941292782050813, 
    0.951903164287363, 0.962549609357703, 0.973218501222434, 
    0.983920104523937, 0.994634810433412,
  -0.994694182246884, -0.984099166095322, -0.973522403226017, 
    -0.962971272008372, -0.952444340540434, -0.941914910901269, 
    -0.931412931972264, -0.920956073973018, -0.910482126791642, 
    -0.900045133344298, -0.889606242525607, -0.879258204104509, 
    -0.868837095674043, -0.858423656942331, -0.848089110427242, 
    -0.837681572504259, -0.827398570112221, -0.817112011574875, 
    -0.806740977758401, -0.796491615936874, -0.786270608799684, 
    -0.776136598447064, -0.765740717256731, -0.755465836473279, 
    -0.745259595136026, -0.735109927749505, -0.72488521812334, 
    -0.714663552329718, -0.704688039797642, -0.694545958981063, 
    -0.684401988594397, -0.674235000585506, -0.664129983710097, 
    -0.65409366169305, -0.643957237416892, -0.634078009910534, 
    -0.623993755114089, -0.613890359576081, -0.603715694726025, 
    -0.593659310543985, -0.583887563685441, -0.57371271539465, 
    -0.563686367676053, -0.553779408534652, -0.543692342484749, 
    -0.533787033947696, -0.523729825394491, -0.513811424279366, 
    -0.503927348570816, -0.494063503183811, -0.484083987424097, 
    -0.474307287316419, -0.464338328938002, -0.454486487506414, 
    -0.444601176362202, -0.434450205047074, -0.424848333901144, 
    -0.414986733415156, -0.40506455572087, -0.395151655229203, 
    -0.385319455606564, -0.375526742161562, -0.365659095350139, 
    -0.355686313200388, -0.346025365407425, -0.336155335757166, 
    -0.32646986846727, -0.316640950103587, -0.306517540521335, 
    -0.297123234801246, -0.287324528487555, -0.277471432053945, 
    -0.267857737455988, -0.258003049311146, -0.248172792638581, 
    -0.238665103639762, -0.228566108296976, -0.218721427258061, 
    -0.208785816367094, -0.199379161595251, -0.189586528264357, 
    -0.179755602125755, -0.170221876933545, -0.160220622482511, 
    -0.150727143224567, -0.140879949838713, -0.130981672610954, 
    -0.121414763299848, -0.111846277535995, -0.102149459679616, 
    -0.0923824090330273, -0.0826102655836689, -0.0728371800140145, 
    -0.0630830285455302, -0.0533898986767289, -0.0437316359226316, 
    -0.0340845375746679, -0.0244057431954076, -0.0146876679959861, 
    -0.00478761741870605, 0.00474845559809092, 0.0145693423247992, 
    0.0243530837385377, 0.0338507222383155, 0.0439373578296853, 
    0.0534581734405978, 0.0630176401315458, 0.072827582179564, 
    0.0828585057758141, 0.0921580064002939, 0.101965277652176, 
    0.111831620430093, 0.121239915149529, 0.131326606893815, 
    0.140852531941982, 0.150798928722556, 0.160522077366389, 
    0.170099136556676, 0.179803845412472, 0.189760496966271, 
    0.199205797298498, 0.209028347755097, 0.218867711031739, 
    0.228669843930535, 0.238098056924593, 0.248100736159725, 
    0.258042092705996, 0.267553779399921, 0.277454182730479, 
    0.287290508733242, 0.296999887263543, 0.306806562832562, 
    0.316465508937647, 0.326421514724141, 0.336150302646254, 
    0.345998257790824, 0.355793759702537, 0.365730873997327, 
    0.375650488940115, 0.385278104790174, 0.395152276767115, 
    0.405164258578882, 0.415011688705053, 0.42447992594258, 
    0.434600090368624, 0.444742769164155, 0.454121605272988, 
    0.464299318465419, 0.474174089375368, 0.484109030278379, 
    0.493919294630207, 0.504010477434431, 0.513882526818777, 
    0.523944558990561, 0.533857465686257, 0.543797620092008, 
    0.553711412803314, 0.563676641816526, 0.57370502172235, 
    0.583727021483643, 0.593678792391568, 0.603768200592222, 
    0.613694809867662, 0.623816385463647, 0.633756148874669, 
    0.643978190027587, 0.654069564884117, 0.664286326877252, 
    0.674185538566536, 0.684559370643148, 0.694644601232969, 
    0.704712512532488, 0.714764033235629, 0.724997533376346, 
    0.735171538980164, 0.74541333884402, 0.755558474836011, 
    0.765790037287862, 0.776053275291095, 0.786307132926009, 
    0.796455077139159, 0.80675914627069, 0.817120074049172, 
    0.827363604780514, 0.837677187926937, 0.848067055613501, 
    0.858510191944428, 0.868760989173496, 0.879175823938103, 
    0.889585981624171, 0.900009977225504, 0.910473727035331, 
    0.920947929464182, 0.931427236920758, 0.941925488597552, 
    0.952434613852882, 0.962970706013415, 0.973526631104752, 
    0.984095783923086, 0.994692444206207,
  -0.994744136971824, -0.984243836455627, -0.973744669299788, 
    -0.963265046968628, -0.952820399885881, -0.94240049516178, 
    -0.931941641426355, -0.921514139899763, -0.911166004011096, 
    -0.900771450329224, -0.890398549564881, -0.880075840472971, 
    -0.869700494792618, -0.859436839903748, -0.849101033591748, 
    -0.838815282319887, -0.828568522648094, -0.818259319976366, 
    -0.807956996920879, -0.797748336587122, -0.787496621972783, 
    -0.777310322248543, -0.767082882059885, -0.756936353886887, 
    -0.746868628155218, -0.73663754482703, -0.726317754759035, 
    -0.716274268028651, -0.706143751472239, -0.696076120623272, 
    -0.685841063565708, -0.6758072668996, -0.665689002547998, 
    -0.655543504456488, -0.645546392957567, -0.635538821864322, 
    -0.625514536621247, -0.615378575309581, -0.605336631106675, 
    -0.595336067418169, -0.585347178579864, -0.575434156116686, 
    -0.565241976291344, -0.555260703954595, -0.545335387817901, 
    -0.535451024111291, -0.525321461954854, -0.515508493962544, 
    -0.5055418352517, -0.495695038394408, -0.485826006548925, 
    -0.475838918130142, -0.465704892913484, -0.455940030527077, 
    -0.445939904681816, -0.435966926368652, -0.426165575585778, 
    -0.416271411459794, -0.40634631253874, -0.396749648800077, 
    -0.38676439813823, -0.376878629102946, -0.366913832206517, 
    -0.357049701334038, -0.347463924249558, -0.337325392805368, 
    -0.327545116073302, -0.317710154337063, -0.307857327235722, 
    -0.298109001589703, -0.2885200806903, -0.278785464206034, 
    -0.268898677007291, -0.258611482752931, -0.249126752473714, 
    -0.23950893064398, -0.229485140344274, -0.219719214490354, 
    -0.209997537615297, -0.200046979553335, -0.190341261038226, 
    -0.180363213764573, -0.170826089442747, -0.161051730036036, 
    -0.151125423725656, -0.141555732540656, -0.131886210110755, 
    -0.12200718249265, -0.112119472872917, -0.102627439111026, 
    -0.0928272137454633, -0.0828207981077821, -0.0733519110953639, 
    -0.0633677598031223, -0.0536031341271215, -0.0439382728129183, 
    -0.034133644252019, -0.0241321909492238, -0.0146058876875026, 
    -0.00509833652052196, 0.00472632320588959, 0.0144378653076708, 
    0.0243969815722766, 0.0343063690103649, 0.0439487992706406, 
    0.053725166222745, 0.0633497230863377, 0.0732982806444437, 
    0.082877792069296, 0.0927642279595195, 0.102283005342417, 
    0.1121031310197, 0.121867164362528, 0.131789229169441, 0.141698627822818, 
    0.151360219547126, 0.160874788553651, 0.170895616148524, 
    0.180709924812117, 0.190337025531381, 0.200187359479196, 
    0.209844185819226, 0.219707709372489, 0.22937595555958, 
    0.239316819720142, 0.248915417023519, 0.258985074771385, 
    0.268916991165979, 0.278655375300963, 0.288353983520322, 
    0.298009794085901, 0.307959618018171, 0.317724579774626, 
    0.327676031550891, 0.337531983649163, 0.347341450484173, 
    0.357222325471791, 0.367071911012042, 0.376866293960447, 
    0.386892077614257, 0.3965428676215, 0.406333091761022, 0.416305459258888, 
    0.426308645594361, 0.436070158801753, 0.445954213242971, 
    0.455996837889759, 0.465747101462405, 0.475803270013006, 
    0.485582179558521, 0.495668733121707, 0.505597828215163, 
    0.515465977826767, 0.525380708235332, 0.535453736201439, 
    0.545281577521213, 0.555383031136358, 0.565269036610601, 
    0.575405451134272, 0.585414748822044, 0.595416184410865, 
    0.605366693544521, 0.615493751010194, 0.625326719640693, 
    0.635541086629236, 0.645592856265308, 0.655601650791708, 
    0.665690062070725, 0.675753268489123, 0.685892039538735, 
    0.695991210547321, 0.706168389094367, 0.716306709842004, 
    0.726436854543487, 0.736603939256173, 0.746681226652746, 
    0.756887412673229, 0.767108667071859, 0.77724262888499, 
    0.787479486782588, 0.79774141229471, 0.807987212685337, 
    0.818215038742303, 0.828550233928544, 0.838787100162222, 
    0.849069674529344, 0.859407866003497, 0.869735295216097, 
    0.880029378421767, 0.890407552667767, 0.900787170353523, 
    0.911165940632745, 0.92152650396169, 0.931942999945397, 
    0.942355594631857, 0.952795038516049, 0.963259652496289, 
    0.973751199013294, 0.984245467229543, 0.994744566894841,
  -0.99477710167711, -0.984336801907834, -0.973912001278027, 
    -0.963511228799046, -0.953100970275106, -0.942726478454335, 
    -0.932348685589247, -0.922028004415207, -0.911636388297688, 
    -0.901310432281893, -0.891026219483714, -0.880675626530322, 
    -0.870408013017321, -0.860119161370202, -0.849868879500939, 
    -0.83959876192162, -0.829301612784589, -0.819088311286853, 
    -0.808935371245824, -0.798666062651557, -0.788526261339633, 
    -0.778274113889536, -0.768199281383849, -0.758009006057039, 
    -0.747710085650838, -0.737613733729311, -0.727394853360051, 
    -0.717273811001213, -0.707231789385677, -0.697153196465849, 
    -0.687073987476675, -0.677014760586032, -0.666934447076094, 
    -0.656804750128867, -0.646883283671215, -0.636788313793721, 
    -0.626610313312538, -0.616642612061117, -0.606685738560067, 
    -0.59663521665665, -0.586539073282192, -0.576471467009767, 
    -0.566545551054389, -0.556554387502173, -0.546605703550319, 
    -0.536597121141035, -0.526511897407058, -0.516673183865524, 
    -0.506764067967201, -0.496934724464931, -0.486721826881325, 
    -0.476894067363842, -0.467200564927621, -0.457005102676843, 
    -0.447029122628878, -0.437298072834699, -0.427349758595802, 
    -0.417436557106153, -0.407511618709, -0.397628972220545, 
    -0.387834377359077, -0.377905754081533, -0.36800891575769, 
    -0.358065113163251, -0.348109535737467, -0.338349817849735, 
    -0.328532745035032, -0.318916661859696, -0.308820882545402, 
    -0.298978910216241, -0.289077263559905, -0.279278928690671, 
    -0.269487183488867, -0.259839496794536, -0.249896254134928, 
    -0.240048495747017, -0.230124485518156, -0.220545119783778, 
    -0.210606659799498, -0.200654363401012, -0.190890113197237, 
    -0.180930769373965, -0.171363540282574, -0.161598545646344, 
    -0.151774559185138, -0.141753361256156, -0.132144965934802, 
    -0.122265477046447, -0.112633657105536, -0.102615697344761, 
    -0.0930239247636891, -0.0833567866094235, -0.0734047872660528, 
    -0.0636174322931081, -0.0537961638371431, -0.0438646475390571, 
    -0.0342460572842292, -0.0245047821306409, -0.0148796083406308, 
    -0.00476054156883379, 0.00492688868721914, 0.0148116204514408, 
    0.024395410310457, 0.0343186362337029, 0.0440092695164986, 
    0.0539066100927644, 0.0636442488975796, 0.0733372617607293, 
    0.0830201525272478, 0.0929214381719107, 0.102715630930104, 
    0.112656382915281, 0.122255879671889, 0.132083646908693, 
    0.141980682727684, 0.151838524983549, 0.161562912521254, 
    0.171409096770863, 0.180991605943874, 0.190964484678276, 
    0.200684843303332, 0.210359639893846, 0.22040048453801, 
    0.230344754314515, 0.239956916728478, 0.249724326226797, 
    0.259577322662555, 0.269473327952586, 0.279417439877504, 
    0.28908810512088, 0.299088476071204, 0.308730315763953, 
    0.318665083220442, 0.328547050126186, 0.338404746511534, 
    0.348500922480487, 0.357887844993284, 0.368059351414541, 
    0.377827700169821, 0.387864671622016, 0.397603003368493, 
    0.407481238694661, 0.417471620070317, 0.427355021580345, 
    0.437207628987481, 0.447037572282714, 0.457068149896447, 
    0.467093109020725, 0.476939855460736, 0.486786230262419, 
    0.496663086586097, 0.506797615276478, 0.516723187288886, 
    0.526641199112078, 0.536663046544673, 0.546553705212093, 
    0.556477869977839, 0.566514050060397, 0.576603972026723, 
    0.586558774622509, 0.596505492671259, 0.60663917211721, 
    0.616621567401843, 0.626617364042515, 0.636726036375193, 
    0.646750978702413, 0.656806572801861, 0.666968069207969, 
    0.67699615316937, 0.687026319416905, 0.697244837860672, 
    0.707282487807145, 0.71729732491746, 0.727513994327745, 
    0.737620999539897, 0.74773961826797, 0.757983862343323, 
    0.768142017610099, 0.778174147425243, 0.788503616543952, 
    0.798633988049461, 0.808959190376076, 0.8191175075665, 0.82936804301023, 
    0.839662603371586, 0.849867240860214, 0.860107977684209, 
    0.870415642220907, 0.880692633335634, 0.891002425076391, 
    0.901339978727254, 0.911608487263155, 0.922009483075548, 
    0.932358071005065, 0.942729713304913, 0.953081819406105, 
    0.963503472584482, 0.973900603290484, 0.984333277634754, 0.994775108007685,
  -0.994803824644056, -0.984416756505597, -0.974035579095254, 
    -0.963676836757954, -0.95331372492289, -0.942978780842939, 
    -0.932654776615598, -0.922322771495273, -0.912022871254781, 
    -0.901757560778523, -0.891424779900476, -0.881181539237402, 
    -0.870908545013648, -0.860630165744525, -0.850432202598101, 
    -0.840193930203666, -0.829960664624803, -0.819753032688907, 
    -0.809597377173866, -0.799390349538532, -0.789239049747755, 
    -0.779044179846492, -0.768917248567993, -0.758711547068538, 
    -0.748632652415962, -0.738436855368331, -0.728327785127145, 
    -0.718213704059506, -0.708130498578061, -0.697960745251774, 
    -0.687925663754715, -0.677889521190995, -0.66776632986241, 
    -0.657763853645391, -0.647613973595461, -0.637547318812313, 
    -0.62757191599849, -0.617519305943945, -0.607573189300652, 
    -0.597527229270706, -0.587554175626346, -0.577516507228584, 
    -0.567548143328573, -0.557459881576765, -0.547514194062478, 
    -0.537516720315198, -0.527622850439276, -0.51750528503226, 
    -0.507564257601666, -0.497629479586796, -0.487751771570675, 
    -0.477893385772881, -0.467933317658109, -0.457927251227132, 
    -0.448091004208667, -0.438077462739041, -0.42822506272886, 
    -0.418182894985559, -0.408379487647169, -0.39838760621012, 
    -0.388513346123537, -0.378746569653267, -0.36880593088788, 
    -0.358893401212143, -0.349016389409073, -0.339012772359341, 
    -0.329186814716671, -0.319461280825844, -0.309416485704597, 
    -0.299593048121151, -0.289808767649663, -0.279922716079631, 
    -0.270089030953387, -0.260357967453311, -0.250468323335924, 
    -0.240553115022658, -0.230747915433919, -0.2209361522366, 
    -0.211092966456632, -0.201289755902449, -0.191284029150291, 
    -0.181539366892418, -0.171878061946726, -0.161997594128141, 
    -0.152111415897382, -0.14219759703672, -0.132676904755942, 
    -0.122694949110275, -0.112884073778839, -0.103029982497415, 
    -0.0931092770551616, -0.0833606528820154, -0.0733276388607167, 
    -0.0637584245094983, -0.0537775395957463, -0.0441027425153438, 
    -0.0342489635629441, -0.0245082997109253, -0.014608765268722, 
    -0.0050371893579197, 0.00481956623393169, 0.0147196355905571, 
    0.0245868649831837, 0.0343759742327581, 0.0441972302536048, 
    0.0539453224933923, 0.0638286213519449, 0.0737110381845632, 
    0.0833635770593505, 0.0932845134238733, 0.10296297187008, 
    0.112648269405858, 0.122632678422835, 0.132498992812101, 
    0.142125254376619, 0.151981922561905, 0.161631011943247, 
    0.171737712221275, 0.18153392218389, 0.191261958894408, 
    0.201182079608993, 0.211097075072209, 0.221104964956296, 
    0.23060745360006, 0.240686257422712, 0.2504579529287, 0.260205895564967, 
    0.270113709072038, 0.279867522220314, 0.289879215517758, 
    0.299654411056213, 0.309372214826541, 0.319295735349344, 
    0.329300087644066, 0.339140552501705, 0.348957484465756, 
    0.35893193008782, 0.36872652213799, 0.37877858372952, 0.388585509492218, 
    0.398347853687892, 0.408312661753852, 0.418111588323929, 
    0.428227610431515, 0.438025817496282, 0.447931154297961, 
    0.458066285316457, 0.46798055114172, 0.477645072755499, 
    0.487702431156225, 0.497851952412664, 0.507636409370793, 
    0.517434199301946, 0.527645887572147, 0.537547897938443, 
    0.547486552756825, 0.557496252006596, 0.56750994580713, 
    0.577516608328793, 0.587513381643578, 0.59752915424229, 
    0.607511421901266, 0.617475660003778, 0.62771161326947, 
    0.637598125482994, 0.647665001816274, 0.657618597944583, 
    0.667810306628985, 0.677837708515305, 0.687934541368609, 
    0.698056288525676, 0.708138072348196, 0.718242767484332, 
    0.728432913139573, 0.73843987587851, 0.748590904761887, 
    0.758755297350241, 0.768939091625949, 0.779037443687406, 
    0.789216187397952, 0.799410596390982, 0.80957999984041, 
    0.819782847086682, 0.830035207821155, 0.840184028870013, 
    0.850451275131526, 0.860665787253713, 0.870911543372882, 
    0.881196095021928, 0.891430887146812, 0.901722819497326, 
    0.912065219068925, 0.922341566865461, 0.932663409107543, 
    0.942971901368606, 0.953324072419761, 0.963660362974191, 
    0.974040801465008, 0.984410342917171, 0.99480143273287,
  -0.994820515679115, -0.984469818436296, -0.974127776485577, 
    -0.963802367546424, -0.953505767503069, -0.943164001734184, 
    -0.932907270724607, -0.922624892630645, -0.912299552750109, 
    -0.902046006222436, -0.891816784567183, -0.881563387729318, 
    -0.871324537387645, -0.861103903113358, -0.850938155932769, 
    -0.840718632273764, -0.830475590913017, -0.820243335915016, 
    -0.810161574062437, -0.799973522797401, -0.789860536915488, 
    -0.779650677041529, -0.769553810448037, -0.759356794121191, 
    -0.749304731097679, -0.739066556501393, -0.728970932622756, 
    -0.718877726794835, -0.708815926361929, -0.698752200085373, 
    -0.688634336110253, -0.678584056226358, -0.668516911521046, 
    -0.658459133438432, -0.648431552729741, -0.63836660173524, 
    -0.628306310735288, -0.618357137543319, -0.608234762589394, 
    -0.598370123351621, -0.588176051935754, -0.578181622990902, 
    -0.568300170736481, -0.558099589824255, -0.548282547134812, 
    -0.538374025534617, -0.528190607153301, -0.518303683801915, 
    -0.508478480049902, -0.498499205010614, -0.488424477391581, 
    -0.4785157921255, -0.468541949376022, -0.458473655160028, 
    -0.44873277999162, -0.438688634337889, -0.428847231128082, 
    -0.418950029890678, -0.409081682882423, -0.399081394248747, 
    -0.389194894911945, -0.379323305602947, -0.369451722424112, 
    -0.359336233887183, -0.34962593968621, -0.339695925425467, 
    -0.329687030190934, -0.31997415327298, -0.309920695717186, 
    -0.300181519910546, -0.290218445234005, -0.280495051673291, 
    -0.270630089547453, -0.2607080081685, -0.25086046429136, 
    -0.241000657398851, -0.231111860976393, -0.221458468798566, 
    -0.211438902756363, -0.201676608748381, -0.191926625424158, 
    -0.181915724881603, -0.17191392037288, -0.162286401174435, 
    -0.1524708305409, -0.142555535110346, -0.132775033030402, 
    -0.122883452204822, -0.112945791853318, -0.103218041078609, 
    -0.0933982745685819, -0.083704088796223, -0.0735727300441927, 
    -0.0637780779844809, -0.0540372764940887, -0.0442901417314782, 
    -0.0345426106263208, -0.0245738593483934, -0.0148703532225334, 
    -0.00466546082744832, 0.00484288310579304, 0.0148027114795735, 
    0.0245628151347185, 0.0342673170807692, 0.0442895523781737, 
    0.054166085885025, 0.0636156889674471, 0.0736060571647462, 
    0.0834588738912711, 0.0932109341172675, 0.103233559169171, 
    0.113165233499963, 0.122819138264997, 0.132688789968513, 
    0.142376127322684, 0.152551135295008, 0.162169590625845, 
    0.17180508581458, 0.181989281398488, 0.191543124076463, 
    0.201417549051675, 0.211460540417925, 0.221486262798927, 
    0.231306621068021, 0.241045247899838, 0.251034168465793, 
    0.260528491150193, 0.270452273876007, 0.280368261468382, 
    0.290234407128257, 0.299993922583426, 0.310018106876027, 
    0.319910260433589, 0.329833993870587, 0.339720507531785, 
    0.349761263201073, 0.359532243254665, 0.36927098786695, 
    0.379347220975655, 0.389284745233179, 0.399129564494383, 0.4089576867211, 
    0.418986719969502, 0.428736499266605, 0.438849683436844, 
    0.448725407712449, 0.458530154582448, 0.468521995338013, 
    0.478464343439436, 0.488444189912942, 0.498380928457659, 
    0.508365520713536, 0.518321500309958, 0.528375991407925, 
    0.538243497188615, 0.548310940982012, 0.558289007043661, 
    0.568199809114568, 0.578356338241752, 0.588175273135904, 
    0.598216496091174, 0.608278648697089, 0.6183289961317, 0.628385595458955, 
    0.638396127525036, 0.648323951343414, 0.65839939666191, 
    0.668405502537226, 0.678607978603145, 0.688671711140137, 
    0.698741144698678, 0.708751133959714, 0.718932743910462, 
    0.729136423294121, 0.739170785407747, 0.749264054817531, 
    0.759316556906265, 0.769512634937564, 0.779687643030587, 
    0.789823908754227, 0.799945714507524, 0.810173935228218, 
    0.820328301987532, 0.830493766834885, 0.840741902450177, 
    0.850920289021957, 0.861091936011362, 0.871349039690304, 
    0.881592381659248, 0.891823225579628, 0.902022078845994, 
    0.912317865435811, 0.922579607935993, 0.93291043519451, 
    0.943183971511401, 0.95350226328517, 0.963801905651335, 
    0.974135124558356, 0.984471581739587, 0.99482227437698 ;

 alpha =
  0.941971411979642, 0.890372174189576, 0.855457936440095, 0.827648539850122, 
    0.801040898409193, 0.778370250756263, 0.75741266981186, 
    0.738870967721304, 0.719792602794716, 0.699799215798082, 
    0.68462041040326, 0.667453632253247, 0.65109731116906, 0.637942182644103, 
    0.621366827664438, 0.60471685655616, 0.591744795838105, 
    0.577979103797105, 0.56471100777747, 0.551111401035758, 
    0.536099410207298, 0.524908946957505, 0.511821824488495, 
    0.497593768509651, 0.486729739087715, 0.47782818538474, 
    0.460430646876392, 0.449774090656099, 0.437843165761436, 
    0.428228758341013, 0.418653855693251, 0.402823408390624, 
    0.39378254853699, 0.383272692222386, 0.372050222200181, 
    0.359020494099934, 0.350039626427997, 0.341971804677645, 0.3303919664145, 
    0.318743998733199, 0.305728630903301, 0.299678905828266, 
    0.291539454229683, 0.282387649208999, 0.271374432593072, 
    0.264649372895653, 0.253489154954366, 0.245121975963024, 
    0.23600565405276, 0.226183501231076, 0.218754882799658, 
    0.211729164695445, 0.204411496975853, 0.192824188219401, 
    0.18758497079937, 0.180495451427352, 0.168493153120849, 
    0.164987295846107, 0.155692875505351, 0.147157424972915, 
    0.142535765778468, 0.136812813908736, 0.127611662209296, 
    0.122245106975645, 0.115489811986656, 0.110479120145545, 
    0.103046906748027, 0.0971016372859742, 0.0898007350529342, 
    0.0857007968608833, 0.083105462966314, 0.0763348257035983, 
    0.070420849627699, 0.0654980006344216, 0.0616776120150308, 
    0.0563977801899388, 0.0511195096830455, 0.0482936589713996, 
    0.0425287535923744, 0.038957594914545, 0.0369521843566832, 
    0.0324915577115838, 0.0287672826747158, 0.0266984985708136, 
    0.0221989982564453, 0.0206213104860163, 0.0177447883280264, 
    0.0152724494574059, 0.0118671507570594, 0.0108769828594946, 
    0.00911046508744617, 0.00709593909471686, 0.00546961764767395, 
    0.00375183020293232, 0.00280867347721329, 0.00223438367788693, 
    0.00108503889809188, 0.000671165628046408, 0.000287474315095419, 
    2.49054139325047e-05, 2.81376986922422e-05, 0.000267609392590756, 
    0.000602810181254535, 0.00127990728369986, 0.00201424503631129, 
    0.00258772556279946, 0.00458745790028635, 0.00545198665595981, 
    0.00690819587414125, 0.00851483970667737, 0.0108535961938689, 
    0.0127331432715305, 0.0145068325784506, 0.0169240186585914, 
    0.0203329688655853, 0.0225627905795494, 0.025866529461559, 
    0.0284699403601827, 0.0311396318357604, 0.0354768229204748, 
    0.0392469061972291, 0.0423204503195557, 0.0469424326836949, 
    0.0509815725006884, 0.0562818413213769, 0.061058557040707, 
    0.0662537024752682, 0.0712369844854457, 0.0771824572219134, 
    0.0809118844685321, 0.0861146366154782, 0.0936622082353179, 
    0.0966515714171497, 0.104054021704001, 0.111098457655426, 
    0.116290017716938, 0.122408116558254, 0.13030941675394, 
    0.135972417560166, 0.14156493950507, 0.14863342667366, 0.157951906556004, 
    0.166821491554412, 0.172112627685093, 0.178788428122975, 
    0.188075217821636, 0.193866331250586, 0.204803244262765, 
    0.210763177031335, 0.221327533744105, 0.225833314523656, 
    0.235938111705536, 0.247835847474225, 0.254027135914529, 
    0.264438332352001, 0.274696204779882, 0.283191442536686, 
    0.29089664476864, 0.303144822461248, 0.308754906860808, 
    0.323571795416045, 0.330485776693124, 0.339685169009913, 
    0.350913435383466, 0.357863812859743, 0.37181270976081, 
    0.383345692630838, 0.393404989245694, 0.403470502786035, 
    0.413629059531547, 0.426301027105689, 0.436644442409969, 
    0.44833806165474, 0.460464287666772, 0.473423560145414, 
    0.486640823296576, 0.489969859372795, 0.513593700965976, 
    0.524812584569409, 0.536715733251959, 0.549209936354771, 
    0.564946573300357, 0.577001167085799, 0.590534564132847, 
    0.604497216978491, 0.620208572154406, 0.635600175356967, 
    0.651899759779916, 0.668287502797153, 0.686304753175652, 
    0.702737063030184, 0.719856499690872, 0.738313820777173, 
    0.758884776921388, 0.780457022697666, 0.802393495352851, 
    0.826403806326829, 0.855448534333266, 0.890173927613311, 0.942380034933993,
  0.979501040899984, 0.950726505933569, 0.928266417161119, 0.908322187041686, 
    0.89009944442857, 0.872780947706181, 0.856580911479208, 
    0.841477227143122, 0.827195309889691, 0.811404203442365, 
    0.797681065639475, 0.783673416848928, 0.769975565845272, 
    0.757086757043869, 0.743858338085241, 0.731747686248755, 
    0.718978298742539, 0.706364494427921, 0.693032231253437, 
    0.680540472734594, 0.66971600693672, 0.654980481038675, 
    0.644718058964097, 0.63265318862909, 0.620237398341047, 
    0.607033536203212, 0.59560230650014, 0.582447999993776, 
    0.569769899807917, 0.559990286529947, 0.550121466885555, 
    0.533501114782263, 0.525849973303723, 0.512776132504931, 
    0.50213133114004, 0.489638829237088, 0.478603319648348, 
    0.467892647722723, 0.454165147667577, 0.442349549362215, 
    0.432289679546919, 0.424112774813692, 0.410454151842396, 0.3997264899472, 
    0.38760852047686, 0.375125688666296, 0.36387977312129, 0.353572327541557, 
    0.34466791543429, 0.333784251120176, 0.323233550171395, 
    0.308241985075636, 0.300267425269652, 0.289443711915357, 
    0.279107703244583, 0.26827018938847, 0.261719923200379, 
    0.250238505342526, 0.239608168276601, 0.230323373065706, 
    0.219840385753618, 0.208313449240947, 0.200873730456899, 
    0.189671151396118, 0.183533625987249, 0.171678643947949, 
    0.165619780987501, 0.15542409181543, 0.146650101143022, 
    0.136738479572638, 0.127483154696351, 0.12054012704935, 
    0.113527849447266, 0.106030348347296, 0.0991097664676841, 
    0.0889134599768556, 0.0845440197412274, 0.0767081868386003, 
    0.069958800720344, 0.0650436031665829, 0.0589952179080345, 
    0.0533382435466026, 0.0474493770886694, 0.0430058927930528, 
    0.0369327718159463, 0.0332739936207679, 0.0288536708847983, 
    0.0240574318397213, 0.0214274217813009, 0.017250214898168, 
    0.0142727640402949, 0.0121474074053256, 0.00911821639296565, 
    0.00687923730243646, 0.0050020230575756, 0.00326245908824322, 
    0.00201200329534115, 0.000887975454823172, 0.000413222312827284, 
    1.26307235871681e-05, 5.69730257972558e-05, 0.000376579531332325, 
    0.0010446012477404, 0.0017805465600725, 0.0031211741550189, 
    0.00501798821026709, 0.00659664855638742, 0.00879460708907441, 
    0.011075537635831, 0.0148061106959316, 0.0170575148825207, 
    0.0215010957135247, 0.0250182325521378, 0.028488353909651, 
    0.0328881999903532, 0.0378892552662653, 0.0431845655574967, 
    0.04757031050165, 0.0521684549171392, 0.0592125404385253, 
    0.0637792013309591, 0.0711386899304746, 0.0777345131066138, 
    0.0833759112710289, 0.0919786324117245, 0.0972533764308887, 
    0.105331947355772, 0.113188598965716, 0.120933830835353, 
    0.127121151722602, 0.137644445456766, 0.145086230438086, 
    0.156694175000553, 0.164494496126493, 0.17100725072112, 
    0.180896802686845, 0.188945899002542, 0.199566838902591, 
    0.20842395796099, 0.220908863443533, 0.229603359993515, 
    0.237896082208552, 0.248460959960073, 0.257340688276849, 
    0.269106734220672, 0.27964647095725, 0.292849241021656, 
    0.300062610354874, 0.311233045850827, 0.321647812977146, 
    0.333766192746806, 0.345861117448926, 0.353258836256032, 
    0.36706270432868, 0.375181811337002, 0.390502758007296, 0.401545838178, 
    0.409700700012194, 0.42210489674881, 0.433774712847055, 0.44347376686565, 
    0.456631284802164, 0.468024751762533, 0.481360837743467, 
    0.490127420470193, 0.501347109817842, 0.514020015565743, 
    0.525786494077836, 0.535575080096428, 0.548857090838415, 
    0.558681784158194, 0.571958781057693, 0.584134908844709, 
    0.595601532495695, 0.608161892878119, 0.620370506819888, 
    0.63098597034493, 0.646055347722015, 0.655792887473987, 
    0.668258491221032, 0.681122316485172, 0.694428343335321, 
    0.706115451994681, 0.719163195294308, 0.732101071005943, 
    0.744460654358231, 0.756361093445139, 0.770233281003129, 
    0.78352623936475, 0.797197137216119, 0.812024985717482, 
    0.825932090728021, 0.840178732696211, 0.85630546786722, 
    0.873108167261289, 0.889792568344144, 0.908529803571236, 
    0.927819554358463, 0.950704989411347, 0.979256050973262,
  0.990382428585975, 0.973478032791684, 0.958615175743594, 0.94502282157381, 
    0.931721292893005, 0.918623107571302, 0.906703596505137, 
    0.894782282572614, 0.882779296463836, 0.871595674058275, 
    0.859694767746939, 0.84929871650206, 0.836731654392462, 
    0.826979487218991, 0.815543625980948, 0.804763454293029, 
    0.793511239149882, 0.782922134125972, 0.772069843756601, 
    0.761234615515719, 0.750355218042746, 0.740659986949899, 0.7280958667103, 
    0.718566186858279, 0.707276995057246, 0.697608826988401, 
    0.686352094314261, 0.674614700144991, 0.663291132528349, 
    0.652002455610202, 0.640887896011799, 0.630733512527774, 
    0.619089085145405, 0.608359956317207, 0.595814585085433, 
    0.585604465704845, 0.571815434400719, 0.562105765751231, 
    0.550167593784241, 0.539770767559323, 0.52707873458026, 
    0.515496894963391, 0.503885561457873, 0.493413850895221, 
    0.480512338291444, 0.468926791143535, 0.456685578919174, 
    0.44529267557412, 0.431904245291833, 0.420180207615755, 
    0.408569690446684, 0.397979271371129, 0.384678920751179, 
    0.374835338552738, 0.361691416931281, 0.34880874523284, 
    0.338342345511548, 0.326917123175221, 0.313849828686517, 
    0.300650960151625, 0.29164871089203, 0.277196414895284, 
    0.266786893094064, 0.254286345948517, 0.243946906146723, 
    0.23281739002213, 0.221599884925874, 0.212231591730368, 
    0.199260647102884, 0.18878261688302, 0.178391939467056, 
    0.166722290423127, 0.155795082001702, 0.146525612596314, 
    0.137132468842552, 0.127368685078316, 0.116065901105936, 
    0.10868878250164, 0.101483778438068, 0.0925401762891319, 
    0.0841553594551581, 0.0764768216321232, 0.0692117884002018, 
    0.060657661931992, 0.0544396823339413, 0.0474720331763457, 
    0.0415385274120335, 0.0360219578462947, 0.0300532917483822, 
    0.024842062831488, 0.0209288385080132, 0.0165842497726198, 
    0.0132117812849521, 0.00974618631020462, 0.00689582166946991, 
    0.00479710449442765, 0.00275132644981613, 0.00141808364773303, 
    0.000652053029822953, 6.73903131642684e-05, 5.66308206872188e-05, 
    0.000497504739455376, 0.00158013431320378, 0.00296244124037001, 
    0.00492897926585323, 0.00719681487757224, 0.0104227569516562, 
    0.0132369996047642, 0.016709966893775, 0.0203265595812056, 
    0.0244256121816096, 0.0295002522499522, 0.03498816436606, 
    0.0415058266772976, 0.047893108748542, 0.0541634232360703, 
    0.0603937581062475, 0.0669252629604866, 0.0765014854043647, 
    0.0835626419230927, 0.0928001807129507, 0.101164535411745, 
    0.110286314038273, 0.11764694338415, 0.128122982196118, 
    0.137298291679198, 0.147297881830559, 0.15681592521238, 
    0.167840578753071, 0.177955375911239, 0.18756469282723, 
    0.199309390406525, 0.211453803460708, 0.220246780245188, 
    0.230679669580981, 0.242788372658455, 0.253795170195133, 
    0.26791843014327, 0.277623121397233, 0.291773414156589, 
    0.302187165958286, 0.313770306702792, 0.324252397478334, 
    0.338012409871106, 0.348729871797754, 0.362336534551584, 
    0.37354218104762, 0.383861740556842, 0.397264760566254, 
    0.410152937479324, 0.420125007648025, 0.433759146252798, 
    0.446274880232529, 0.457160071999176, 0.469163309724955, 
    0.47997166048273, 0.493484521795038, 0.505117526426922, 
    0.517473043956345, 0.527874008269682, 0.538514511724119, 
    0.550476525525113, 0.562357108322109, 0.574876089290276, 
    0.586863754612094, 0.596316865335379, 0.607725262329926, 
    0.619326405035974, 0.630365679250831, 0.643259272570455, 
    0.652907570682112, 0.664843617531786, 0.674981755742561, 
    0.68464871494494, 0.697968221198984, 0.708148989165462, 
    0.718332698961813, 0.72939621915326, 0.739833483767568, 
    0.751045834027705, 0.762213584913685, 0.773675151513281, 
    0.783028310049665, 0.794500412358986, 0.805315667766405, 
    0.815269427609734, 0.826267285178441, 0.837968936545095, 
    0.849317474577955, 0.860533571283943, 0.871432112965855, 
    0.882497765156909, 0.894374305567538, 0.906214272448227, 
    0.919192181357352, 0.931242436725531, 0.944646629988121, 
    0.958616101937595, 0.973557725159042, 0.990411899990964,
  0.99439416767213, 0.983479861698002, 0.972985534772607, 0.962869665053517, 
    0.953186855110061, 0.943566209477211, 0.934298355751344, 
    0.924912417829641, 0.915631898482098, 0.906542769982959, 
    0.897563017220892, 0.887884328771816, 0.878802663993163, 0.8697359213876, 
    0.860271417344794, 0.851251498009766, 0.842771253725378, 
    0.833542954872561, 0.823459912711613, 0.814839456692611, 
    0.805432882426279, 0.795990577427771, 0.787107424026371, 
    0.777080282700362, 0.768129924668169, 0.757889007402457, 
    0.747647699003621, 0.737816344187736, 0.727440511145021, 
    0.718612531576175, 0.708580006303424, 0.697659973339449, 
    0.687464907624043, 0.677617558668486, 0.666869412051231, 
    0.654963599348566, 0.645617559138597, 0.634279526366896, 
    0.622760937373988, 0.612374628278445, 0.600761817150999, 
    0.589235541138461, 0.576548158219662, 0.566235684442701, 
    0.553273800182146, 0.542156924364679, 0.529711045801822, 
    0.517569459995147, 0.507769605617164, 0.494212966695051, 
    0.47994494486202, 0.467512945718966, 0.454874649948325, 
    0.442192976670765, 0.429474395796213, 0.4159355218171, 0.405754951798126, 
    0.392136240387084, 0.380312585957498, 0.365822547168256, 
    0.353650363849259, 0.341214596292093, 0.325740680663126, 
    0.312048012569151, 0.300789408079208, 0.286532389678321, 
    0.274841448542575, 0.262113976131335, 0.249218086208497, 
    0.238168577261509, 0.222567596113641, 0.211136353540832, 
    0.198242732993826, 0.186966452984051, 0.174932089687838, 
    0.162016442806723, 0.151700044984874, 0.140086645659231, 
    0.128336790511605, 0.117908029177737, 0.108655590080391, 
    0.0993163379846448, 0.0883535260361063, 0.0797850499316422, 
    0.0703290547488824, 0.0615995566613737, 0.0535469643962979, 
    0.0461616091243902, 0.0401509247038084, 0.0342778062799574, 
    0.0273377276106038, 0.0224916778238337, 0.0172945860858936, 
    0.0131421158679454, 0.00968212284214999, 0.00620697241930806, 
    0.00399598382223491, 0.001954965150926, 0.00064027924553933, 
    8.98833453632539e-06, 0.000102406905294891, 0.000575253398211186, 
    0.00210654340741691, 0.00388031149452692, 0.00645238953047512, 
    0.00894689176787957, 0.012925419050181, 0.0174956187347099, 
    0.0218576109581398, 0.0276851307077551, 0.032862313000642, 
    0.040508866057588, 0.0465215501802278, 0.0533875698904913, 
    0.0617430888547224, 0.0703336827421395, 0.0793934221076244, 
    0.0874649205682143, 0.0994691623747366, 0.110461635156191, 
    0.118987873744721, 0.130915329408719, 0.139210112293216, 
    0.151298308719143, 0.16387720333537, 0.175350718491482, 
    0.186313763114245, 0.199080740734673, 0.211206003297234, 
    0.221199747372914, 0.23571154414562, 0.250568189290857, 
    0.260579235925716, 0.276174189095071, 0.288617313361069, 
    0.303859255081365, 0.313989878526973, 0.328214548704553, 
    0.340196369541985, 0.351075315947219, 0.368933384737675, 
    0.379600582410322, 0.39198050820149, 0.404642336023242, 
    0.418389952505333, 0.432358156650778, 0.44290284134643, 
    0.455789074845753, 0.468311956696271, 0.480112106368804, 
    0.493253652030061, 0.504112661196767, 0.520108434929751, 
    0.532159704156322, 0.544358086275982, 0.552921834620558, 
    0.56651996406632, 0.576566160815805, 0.588990744811661, 
    0.600644587499202, 0.610352935623216, 0.622052979832262, 
    0.632325106610149, 0.643070447673489, 0.655609567865045, 
    0.667109720794916, 0.677398615862908, 0.688277163871653, 
    0.697762055405025, 0.706883144710971, 0.718662455436109, 
    0.727923496895398, 0.737710276092395, 0.748762399343741, 
    0.757433382793929, 0.767270665349109, 0.776536197322049, 
    0.786736563401236, 0.796260623795304, 0.805652127677219, 
    0.814882964722273, 0.823973472025679, 0.833604063681312, 
    0.842629496459145, 0.851784386599754, 0.860287214856407, 
    0.870005204676763, 0.879277447534784, 0.888378241931235, 
    0.897388632681794, 0.906258667532911, 0.915261619211529, 
    0.924746835167486, 0.933933041118969, 0.943685222396597, 0.9533322962944, 
    0.963172460970086, 0.973013185851533, 0.983516883452454, 0.994367128987061,
  0.996185743012186, 0.988487314612445, 0.980866643121551, 0.973198946346812, 
    0.965768631932266, 0.958223058270813, 0.950570417282883, 
    0.943327842527345, 0.935427347832001, 0.928113639692221, 
    0.920950296569484, 0.912818363162851, 0.905565024271732, 
    0.898199588359247, 0.889784551946136, 0.882240317358648, 
    0.874586321529065, 0.866595709450644, 0.858677559159813, 
    0.850442035045042, 0.842577499272411, 0.834777651864656, 
    0.82621951374056, 0.818032877854088, 0.809519582109149, 
    0.800231435591438, 0.792088509275569, 0.78270382939766, 
    0.774085600264913, 0.76444991591643, 0.756597565128786, 
    0.746300338737422, 0.737623674809078, 0.727250888535597, 
    0.717917355139711, 0.70860789004962, 0.698451532577725, 
    0.688083855687421, 0.677575183721375, 0.667134940591668, 
    0.65667924993397, 0.645378635251782, 0.634599438970639, 0.62411147927815, 
    0.613057053299455, 0.601097384209987, 0.588705562319632, 
    0.576777934470638, 0.565195906121191, 0.552809433959289, 
    0.541420477904436, 0.528137436756389, 0.516766156866957, 
    0.500981112613645, 0.489507081144197, 0.477042551834201, 
    0.464568180388328, 0.450425459219206, 0.435484568467969, 
    0.42230830530972, 0.408466377384038, 0.394644160981079, 
    0.380511232030855, 0.364551778428404, 0.35233831593364, 
    0.340244013143403, 0.324572246403537, 0.310220831452401, 
    0.294221570417551, 0.280399815321418, 0.266286869135619, 
    0.252811238276822, 0.23800553439436, 0.22491289486877, 0.212395889518457, 
    0.196959575740402, 0.184762776543643, 0.171371186596963, 
    0.15793540627981, 0.144608175971075, 0.132180942025947, 0.12219203572586, 
    0.110352506834563, 0.0983778928540792, 0.0878028751879061, 
    0.0774525098684183, 0.0676086174425767, 0.058068001619212, 
    0.0498827892088696, 0.0417364492695667, 0.0344329376271555, 
    0.027266696776454, 0.0219799308540136, 0.0169196248019973, 
    0.0117301680195427, 0.00778989309327862, 0.00463576547368951, 
    0.00247879462196894, 0.000931035094092071, 6.99394035968935e-05, 
    0.000112349593638275, 0.000725059670386912, 0.00254992621287358, 
    0.00468234497631924, 0.00794638535642454, 0.0115681065888769, 
    0.0161318272171734, 0.0220965328797405, 0.0279619361272965, 
    0.0342275141148572, 0.042388615415147, 0.0486100124095784, 
    0.0579660716930058, 0.0674987931228397, 0.0771424113159448, 
    0.0871926517226648, 0.0976518806954927, 0.109899429701798, 
    0.12178943171954, 0.133446201569158, 0.147216077582771, 
    0.159730012057334, 0.172269338593607, 0.183058385823754, 
    0.198603599901942, 0.212203723446085, 0.224471747779648, 
    0.238798015032457, 0.252635368058205, 0.266805136437406, 
    0.281401775781566, 0.294485149474816, 0.307371112501372, 
    0.323323305299665, 0.337300998918854, 0.352564888160764, 
    0.366880175605299, 0.378466659412313, 0.393268507508617, 
    0.409305374705159, 0.423193762596887, 0.436181052153661, 
    0.448436545943272, 0.461561929310659, 0.476971695717007, 
    0.488511628657023, 0.503479509342903, 0.514665890021176, 
    0.527803014169442, 0.540339335863535, 0.552664052719651, 
    0.565783910795515, 0.576202804565107, 0.588675549320949, 
    0.599862511127348, 0.612184391384187, 0.622128965076211, 
    0.635127822048256, 0.645704876681103, 0.657728717781243, 
    0.666033433724872, 0.676349069065988, 0.689149804933245, 
    0.698339298878469, 0.708029978824949, 0.718642913985803, 
    0.728771444560458, 0.737340989152363, 0.746831436509027, 
    0.755950057959623, 0.766226886361387, 0.774180290912784, 
    0.783413018621444, 0.791420176657404, 0.800744499707193, 
    0.80885020903278, 0.818482705523795, 0.826054958634335, 
    0.834323541353894, 0.842937137689985, 0.851347849543883, 
    0.858727051125479, 0.867219205929811, 0.874486532091399, 
    0.88240130647469, 0.890182909104335, 0.897211860140321, 
    0.905425465894417, 0.913309537643014, 0.920697764894495, 
    0.928423259948961, 0.935588193925884, 0.943325130522421, 
    0.950816078131792, 0.958171193551981, 0.965635272161037, 
    0.973265607433865, 0.980910617190242, 0.988519454195895, 0.996209478155432,
  0.997165747676666, 0.991368079370216, 0.985485138882363, 0.979422379691914, 
    0.973405219011164, 0.96729332702691, 0.961170109645585, 
    0.955082100379624, 0.94877156300158, 0.942631975218178, 
    0.936397425244506, 0.929948549995264, 0.923645515213365, 
    0.917059080120445, 0.910518438166212, 0.904008709767467, 
    0.897071462740343, 0.89099320907767, 0.88323500382219, 0.876570480320019, 
    0.869605807697683, 0.862614358890374, 0.854658122674626, 
    0.84793753588321, 0.839976199534265, 0.832498458736809, 
    0.825219270847463, 0.816592431080683, 0.809733085036262, 
    0.800804144882801, 0.792835479174667, 0.784055476230635, 
    0.775063109012075, 0.766932753403996, 0.7579446385924, 0.749589819745418, 
    0.740004928621682, 0.729833873108708, 0.721028245231699, 
    0.710847849497188, 0.702075477483456, 0.690698374136752, 0.6804287833882, 
    0.669024002092734, 0.657439744996919, 0.646830884997623, 
    0.637239952298458, 0.625353182891206, 0.614141273159098, 
    0.600766842553944, 0.590056182881406, 0.577843687827748, 
    0.563709359345008, 0.551240809682449, 0.53884475181582, 
    0.524815980464991, 0.511037040539314, 0.498806292439164, 
    0.483963917204013, 0.471578594747164, 0.456704726839799, 
    0.44196265522054, 0.425934051851018, 0.413021836989822, 
    0.400285456079941, 0.384364466460344, 0.367919673388837, 
    0.353398352006896, 0.338724913688919, 0.323044258508507, 
    0.308409516462936, 0.292188716818457, 0.276640234049683, 
    0.262618488344717, 0.245426838459751, 0.230815857962323, 
    0.214581827770746, 0.200362770929543, 0.185619661588744, 
    0.170678306681875, 0.158655501558169, 0.144027968148634, 
    0.128984695498812, 0.117344854174227, 0.103915025828028, 
    0.0902142359817706, 0.0811868445742816, 0.0704072981508174, 
    0.0608274239665222, 0.0489371116313748, 0.0423033293647834, 
    0.0336363394096253, 0.0256397381614369, 0.0197413536581337, 
    0.0145806689340377, 0.00945591788928205, 0.00547293154991279, 
    0.0031194000116517, 0.00115257952957689, 9.06246296002065e-05, 
    9.07626755580423e-05, 0.00114264551484167, 0.00267999487315226, 
    0.0064119002860716, 0.00932364046800005, 0.0146847067315019, 
    0.0194898378192499, 0.0266126333382193, 0.0338996773373391, 
    0.0414876605211369, 0.0504186150051803, 0.0606317364981513, 
    0.069919062157367, 0.0807220950182465, 0.0930007594463095, 
    0.106791620990048, 0.118247178080219, 0.130128255315042, 
    0.143531310186262, 0.156213597608613, 0.170248654974049, 
    0.185714699747735, 0.199714493441275, 0.214455341683816, 
    0.229761927979253, 0.245282922488731, 0.260134715540481, 
    0.274256359604936, 0.294177765921782, 0.305702345504835, 
    0.321633086071888, 0.338142357082823, 0.35279465197396, 
    0.368547952066792, 0.384147287967628, 0.397416818990123, 
    0.410279318423594, 0.426567195699148, 0.441117065773165, 
    0.457191976616242, 0.472093981294294, 0.485370980916711, 
    0.498993206801353, 0.513213489857703, 0.526581197911642, 
    0.538704261142963, 0.552156929072985, 0.56384285985494, 
    0.576034387532064, 0.59067649033341, 0.601812456512774, 0.61432541164178, 
    0.624588638684064, 0.636767954801067, 0.64824175785756, 
    0.658919533233543, 0.67030057624771, 0.6792871861905, 0.690550369079031, 
    0.700106512487215, 0.711203574334463, 0.720599249027313, 
    0.729359460891135, 0.739802435682788, 0.749372364840991, 
    0.757591894926422, 0.766725320234139, 0.775521968247974, 
    0.784599643771953, 0.792283134566766, 0.800459517551008, 
    0.809776809184622, 0.816928361281692, 0.82521695261579, 
    0.832636859579922, 0.840234208305668, 0.847929507090345, 
    0.855486531896794, 0.862809028795458, 0.869607676311863, 
    0.876901272587837, 0.883384911050089, 0.890582495895725, 
    0.897376555501291, 0.903922885574687, 0.910306882570641, 
    0.917075130594721, 0.92364753644698, 0.929850433924344, 
    0.936446032135801, 0.942562601659008, 0.948936863929396, 
    0.955017561942668, 0.96109865504553, 0.967256274616128, 
    0.973448918206983, 0.979505601042495, 0.985426672257704, 
    0.99136725703104, 0.997162469333754,
  0.998130814989526, 0.994325227711479, 0.990354636801337, 0.986265405234609, 
    0.982110291812041, 0.977742751297831, 0.973450181680316, 
    0.969216688211726, 0.964559756396445, 0.960188120731208, 
    0.955198099568627, 0.950905339517399, 0.945970150356002, 
    0.941088015108032, 0.936096068379213, 0.930968149064449, 
    0.925930885236925, 0.920811463417786, 0.915524482638056, 
    0.909842652489306, 0.903928125348342, 0.898614270602162, 
    0.892918271295551, 0.886628285524953, 0.881054874817378, 
    0.874986257002581, 0.868486199024734, 0.862611984214189, 
    0.856395033880948, 0.849278014634934, 0.842060081167904, 
    0.835201397103627, 0.828287618965731, 0.820423317513852, 
    0.813622534547717, 0.805492400069173, 0.797637294670553, 
    0.790362533761666, 0.781453311638318, 0.773307502921436, 
    0.763736955553361, 0.755165056239946, 0.746315018208803, 
    0.737723335135613, 0.726060224853057, 0.71750290254199, 
    0.708087220618689, 0.696713673444697, 0.685009878999168, 
    0.676579534595739, 0.664546511884542, 0.65419797169496, 
    0.639620262981516, 0.629058702008082, 0.616420932289393, 
    0.604886089559675, 0.592348124318033, 0.575634920537109, 
    0.564027541358008, 0.5494985511042, 0.535893377277878, 0.52064993751751, 
    0.50561617412059, 0.491361487489398, 0.476117908946724, 
    0.460943034501261, 0.444230802893406, 0.427962173065859, 
    0.411226606056846, 0.392639387639948, 0.378816820701553, 
    0.359983314779186, 0.343864429117731, 0.327232077733907, 
    0.307083837724734, 0.29071459995198, 0.272832686891818, 
    0.255572006355461, 0.238630888908999, 0.2210826693645, 0.203645805227056, 
    0.186117448321109, 0.169449377669476, 0.153625975164666, 
    0.136492461493608, 0.122369218606824, 0.106445255960478, 
    0.0934469734496163, 0.0801709202126546, 0.0676281611153137, 
    0.0576654991071268, 0.0459941258254143, 0.0361657141504203, 
    0.0271532506075979, 0.0193782689090998, 0.0131768402737291, 
    0.00805290380147484, 0.00418914000692347, 0.00138471729243034, 
    0.000123677565250761, 0.000173830471483917, 0.00133952356546791, 
    0.00422346134813588, 0.0080481380670123, 0.0135457677372491, 
    0.0193286714450919, 0.0259781900517693, 0.0344410605993792, 
    0.0460206562106134, 0.0561144530201083, 0.0673329225802757, 
    0.0789009039264016, 0.0935116448734731, 0.107611433421964, 
    0.122279857213858, 0.13737069952841, 0.151121355136655, 
    0.168091572805954, 0.186283674234933, 0.203738225518282, 
    0.22073163307482, 0.238203079811857, 0.253802404692057, 
    0.273757263430906, 0.291129261916337, 0.310130064500884, 
    0.32515735262408, 0.344476108381769, 0.359643122898453, 0.37824694642657, 
    0.395889813841049, 0.412256422788562, 0.427683691935362, 
    0.44284369925524, 0.459187603332512, 0.477540448701963, 
    0.492567641308053, 0.505821171487941, 0.521505197658978, 
    0.534492048776394, 0.549973582257258, 0.563663170273153, 
    0.577354212956387, 0.592345504653517, 0.604207946558462, 
    0.615727703395521, 0.629571450907487, 0.640317147742531, 
    0.651539541514857, 0.663714513891731, 0.674895781668857, 
    0.686243586047881, 0.696197472371028, 0.707145021030777, 
    0.717145741779088, 0.727763447585123, 0.736767308420342, 
    0.746190483583696, 0.756142846767972, 0.763638313639142, 
    0.773234120518755, 0.781629359111786, 0.790528040654712, 
    0.797637690920898, 0.805116374375834, 0.81358402673857, 0.82041253908393, 
    0.828349359741684, 0.835368192560903, 0.841722807055211, 
    0.849007149548562, 0.855457143320393, 0.862321879314636, 
    0.868588621777541, 0.874659186598269, 0.881160452449298, 
    0.886802208804914, 0.892478461598338, 0.898895786343303, 
    0.904132874877097, 0.909926179416717, 0.915041665175875, 
    0.92089220263272, 0.925813769279522, 0.931084805534425, 
    0.936121071637125, 0.941122195745124, 0.945822503866658, 
    0.950638980828216, 0.955411720017112, 0.959991907816993, 
    0.964690018626767, 0.968982915242343, 0.973397634276898, 
    0.977809140320148, 0.982163795058843, 0.986309189308784, 
    0.990369392043113, 0.994322708028094, 0.99812721876231,
  0.998620486543181, 0.995798107755665, 0.992858807264233, 0.989807440993649, 
    0.986627247724068, 0.983406661725766, 0.980138759689752, 
    0.976759668986537, 0.97334126311775, 0.96984712827724, 0.966038960256553, 
    0.962534541733702, 0.958860802461258, 0.954908212336856, 
    0.95099148015138, 0.947088571462402, 0.94272998071171, 0.938828222675758, 
    0.93434961552127, 0.929937527024046, 0.925400192408, 0.920633932974429, 
    0.915961369840287, 0.911204399944653, 0.906380596361615, 
    0.900796586203622, 0.896045634470509, 0.890563831273031, 
    0.885544255956052, 0.879654216316817, 0.874136696536657, 
    0.867889803287436, 0.862083655956364, 0.855775475661712, 
    0.849425168221312, 0.842906092494614, 0.836053552845936, 
    0.828922676513041, 0.822204369312836, 0.81494887694019, 
    0.807133260608541, 0.799558363709094, 0.791011928791385, 
    0.782458367521972, 0.774846470698406, 0.765936182900326, 
    0.756148060473708, 0.747169382289939, 0.738736702286915, 
    0.727690192061693, 0.717470553110704, 0.707266662779288, 
    0.695643721650191, 0.68493325290232, 0.674886891918941, 
    0.662085703604891, 0.649117691035388, 0.637538848198812, 
    0.623840925175041, 0.610204779457385, 0.597173133243262, 
    0.583015727796743, 0.567257146304406, 0.553232651470794, 
    0.536936233286077, 0.521744519249508, 0.50649849082887, 
    0.489131098062139, 0.473029046399148, 0.455172076704929, 
    0.437345425048836, 0.420326408064812, 0.401254537948218, 
    0.381957768969345, 0.363005721095979, 0.345020909379978, 
    0.323167332016149, 0.304787229136324, 0.28609690367003, 
    0.265319353116204, 0.247970848025915, 0.22724418606514, 
    0.207762060496393, 0.189280902359439, 0.168988041498004, 
    0.150206303142637, 0.132747922123041, 0.115561597279887, 
    0.0999441233017441, 0.0843442810989759, 0.0704701093077229, 
    0.0574676060218118, 0.0445927644939868, 0.0343786344393682, 
    0.0249327428368402, 0.0166708102168646, 0.0102390453009109, 
    0.00525551126728013, 0.00180355097300272, 0.000219836338784457, 
    0.000177823667514864, 0.00173447850781187, 0.00542664244614094, 
    0.0100287406999326, 0.0172583446567066, 0.0253327584985927, 
    0.0336976030793839, 0.0456602946255008, 0.057635779487418, 
    0.0709446629191043, 0.082888854847564, 0.0988784741810798, 
    0.116466767886954, 0.133272203428362, 0.150248799609163, 
    0.169060936991327, 0.189278384286101, 0.207157582665659, 
    0.225448089120174, 0.244088194351096, 0.26316209860933, 
    0.284590880167989, 0.304250179664117, 0.325265564191917, 
    0.345251009822954, 0.363078225150509, 0.383994812706251, 
    0.401379967050579, 0.418358992732303, 0.438037873233191, 
    0.454211603813995, 0.472164606068182, 0.490592295841651, 
    0.505817235965557, 0.524402743946502, 0.538999480619705, 
    0.551791412295194, 0.570007298678507, 0.583250920264697, 
    0.597512397218644, 0.609301301068601, 0.623014459087405, 
    0.63775002363771, 0.649034113825682, 0.662801641350495, 
    0.673023051811323, 0.685435394681583, 0.696066782424659, 
    0.708408603334291, 0.716313091492823, 0.72842085738261, 
    0.737738599221403, 0.747955293896081, 0.757239011844492, 
    0.765737504027432, 0.77469638615687, 0.782586785169918, 
    0.790674559221354, 0.799648585894773, 0.807512364044838, 
    0.814413482257966, 0.821975606453969, 0.828730033089798, 
    0.836656823428544, 0.843043935642396, 0.849241301101473, 
    0.85590239942532, 0.862228934864497, 0.867973332326405, 
    0.873673290812887, 0.879605535286552, 0.885208049884984, 
    0.890845426692001, 0.896170407956616, 0.901679838286683, 
    0.906277953558263, 0.911211208588887, 0.916123145175575, 
    0.920722068030271, 0.925439963757138, 0.929619190280326, 
    0.934018493706021, 0.938511900795548, 0.942753735562124, 
    0.946852336410459, 0.950899977598915, 0.954789376881393, 
    0.958610242267681, 0.962478663428727, 0.966116991400782, 
    0.969724294498234, 0.973303761140133, 0.976747216795566, 
    0.980100394147996, 0.983415789514796, 0.986653041534866, 
    0.989798532734426, 0.992842246541878, 0.995792881259154, 0.99861862374056,
  0.998778599046271, 0.996274733457679, 0.993710012824724, 0.990993685055853, 
    0.988218322323338, 0.985387193713416, 0.982427872891801, 
    0.979324085576475, 0.976245851625279, 0.973168233953604, 
    0.969910335156288, 0.966487235763925, 0.963272517446514, 
    0.959743235260279, 0.955943897175278, 0.952738492264491, 
    0.948727384658585, 0.944994488909806, 0.941117937725034, 
    0.937166172588778, 0.932967006887398, 0.928904908953113, 
    0.924458722012608, 0.920355687257625, 0.915598948994879, 
    0.911042786481527, 0.906076353996933, 0.901300216017168, 
    0.896380134901697, 0.891395823557809, 0.885978845733847, 
    0.880455334401865, 0.874884644663818, 0.869247150966172, 
    0.862623463836852, 0.857245520812833, 0.85072229473465, 
    0.844221702698593, 0.837716459334212, 0.830612228232157, 
    0.823859776112909, 0.81708786030396, 0.808916777188917, 
    0.800328198511732, 0.793298548574069, 0.78497804655361, 
    0.776602626434809, 0.766813875352452, 0.757979101299489, 
    0.749111812315433, 0.738937152480732, 0.730115415927825, 
    0.718177711168301, 0.709033019414173, 0.696783809294862, 
    0.685173780475499, 0.674550993558714, 0.662299397772925, 
    0.649327647182605, 0.637237603420453, 0.623241588720765, 
    0.609100128869966, 0.593478177827085, 0.579892443824733, 
    0.564557370172745, 0.549143053954469, 0.533336164817788, 
    0.515861381708779, 0.499953534477888, 0.482454317624718, 
    0.462390549302479, 0.446536404457675, 0.428078481155464, 
    0.408204813445672, 0.389120773145621, 0.367600351299486, 
    0.34520200206173, 0.325792240476955, 0.306112596005114, 
    0.286008054269605, 0.265123451088498, 0.244773931924377, 
    0.223935461894075, 0.204617287561474, 0.1833096029263, 0.167105320512018, 
    0.146368880518247, 0.128571283685632, 0.110528546764816, 
    0.0942850674678974, 0.0777514016032248, 0.0625876307387251, 
    0.0487811280045375, 0.0379918488678619, 0.0275648689791325, 
    0.0182693002966395, 0.0112044737629205, 0.00574313532553657, 
    0.00195184783127583, 0.000247783771410977, 0.000255395676704853, 
    0.00204693624469943, 0.00629276402853702, 0.011107294427802, 
    0.018965910626154, 0.0269814477507346, 0.0381220267331434, 
    0.049912350241807, 0.0626479601101414, 0.0772940226304573, 
    0.0938854145639922, 0.109981887628472, 0.128606630751784, 
    0.147156031864283, 0.163785838765444, 0.185412560480408, 
    0.202777142750285, 0.225605300272973, 0.245608004653665, 
    0.266040927757859, 0.286907489979198, 0.308016180609089, 
    0.328276666683754, 0.347597904446802, 0.368292349889307, 
    0.386971485121606, 0.4088968140222, 0.42644671251956, 0.445789139990347, 
    0.466249682434395, 0.480158351443781, 0.49821752633137, 0.51584454440247, 
    0.533059426054137, 0.549304480809543, 0.565279357865705, 
    0.580557961794368, 0.594247184451275, 0.609692992464269, 
    0.621121271240229, 0.63593705316736, 0.648334320244069, 
    0.661382345053721, 0.673197340090292, 0.684743897929873, 
    0.695537483257681, 0.707623226512955, 0.718725266394271, 
    0.729874530849974, 0.739982588468886, 0.748793223674029, 
    0.759174153697227, 0.766916145831267, 0.776280125162668, 
    0.784527872819671, 0.793168705974551, 0.800704552398761, 
    0.808755940769377, 0.815897200342893, 0.823765941856324, 
    0.830620500995798, 0.837500735712558, 0.844568823120938, 
    0.850906457210731, 0.856657789603047, 0.862715745543479, 
    0.868476721716401, 0.874789603135756, 0.880549524926419, 
    0.885763100628273, 0.891271327537877, 0.896553097021395, 
    0.901466421991019, 0.9061574641517, 0.911111906819739, 0.91575827469481, 
    0.920111490615869, 0.924429506327917, 0.929074348000948, 
    0.932762353876303, 0.937174951751174, 0.940857183173784, 
    0.944970969681575, 0.948667361135901, 0.952540721275515, 0.9563044975466, 
    0.959596861306932, 0.96317269773295, 0.96655923128845, 0.969866029807437, 
    0.973220318290502, 0.976373177211956, 0.979447079955702, 
    0.98241470303239, 0.985354821496025, 0.988231856514896, 
    0.990970914422807, 0.993700386053839, 0.996301546169151, 0.998779545459298,
  0.998900136653537, 0.996665864176002, 0.994327448046302, 0.991955489466112, 
    0.989425746070923, 0.986830460063615, 0.984237696289428, 
    0.981566245104066, 0.97871946879726, 0.975894869757984, 
    0.972921732014535, 0.9699629072461, 0.966779320340236, 0.963679049696698, 
    0.96047140816149, 0.957205934191983, 0.953650078599754, 
    0.950228678644546, 0.946720244231987, 0.943059324427352, 
    0.939324263502894, 0.935506563794094, 0.931551716736025, 
    0.927322222162755, 0.923439281592724, 0.91881830390475, 
    0.914687144757817, 0.909964492445661, 0.905800064354607, 
    0.900593844528779, 0.895771571565224, 0.890675444052702, 
    0.885888163348937, 0.880040303683711, 0.87530965269329, 
    0.869272949465707, 0.863361323122075, 0.857031143408317, 
    0.851096448029843, 0.844041934837538, 0.837825321010583, 
    0.830919855059678, 0.82403304511649, 0.817307828281869, 
    0.808931098695221, 0.801205201856668, 0.792621607450702, 
    0.784084165771576, 0.776698828666517, 0.767554034650588, 
    0.75744414571883, 0.747759112579753, 0.737959126439338, 
    0.727315041220656, 0.717677557389621, 0.70798689063068, 
    0.695035979520451, 0.682678169933418, 0.669870864806337, 
    0.658248079830834, 0.645100573687094, 0.63130846045988, 
    0.617566761635708, 0.603914486261381, 0.587496338754827, 
    0.573477481544091, 0.556457707134455, 0.538763518993168, 
    0.523341910318116, 0.505168300721553, 0.486155689633336, 
    0.468887830548732, 0.447780884726896, 0.430865898257123, 
    0.411173642120319, 0.391262480816428, 0.370303757191134, 
    0.349828312746381, 0.328241550967753, 0.307065205704644, 
    0.285547186515161, 0.264590809731524, 0.241819372739912, 
    0.220210262820597, 0.199429777166176, 0.178844737318698, 
    0.158098881963903, 0.138582312053364, 0.119093673797902, 
    0.100903545751669, 0.085347744644426, 0.0685839926910951, 
    0.0549029646972995, 0.0418643540362049, 0.0302740102337264, 
    0.0197786016343756, 0.0124109879539676, 0.0060964212027756, 
    0.0024615774449537, 0.000202371495313487, 0.000273608769906642, 
    0.00223319190127867, 0.00578903041186027, 0.0126100098986408, 
    0.0195816114417461, 0.0294059603792516, 0.0412303027489332, 
    0.0554105946710857, 0.0692616679545127, 0.0851458333944715, 
    0.102054967557503, 0.11989738411239, 0.140255581947716, 
    0.158004750706358, 0.17880322943499, 0.199184071070802, 
    0.219001770209206, 0.241434982137302, 0.262154351913874, 
    0.283682037732307, 0.306218860544261, 0.327906838227942, 
    0.350432800038761, 0.371326931722734, 0.390393380821844, 
    0.411334667368911, 0.431832480945549, 0.450547447754663, 
    0.468774133901123, 0.488199618375965, 0.50373894414038, 
    0.523088460800454, 0.540207853759937, 0.555677117431939, 
    0.572024394473514, 0.588270427590232, 0.601470947747097, 
    0.616918044897907, 0.632478304593113, 0.643951140007518, 
    0.65841402211537, 0.670650295197151, 0.682720313605879, 0.6941621970869, 
    0.707032323701081, 0.717066016587233, 0.728421507546051, 
    0.738291696573793, 0.747935123297862, 0.757563422820454, 
    0.766807018761637, 0.77667373655166, 0.784831163656514, 
    0.793738786637344, 0.801364785702393, 0.809181275656411, 
    0.816403806340259, 0.823955858724538, 0.830898567265794, 
    0.837706562891939, 0.844216836892033, 0.851071579514199, 
    0.857227894384588, 0.863044723493272, 0.868695900699787, 
    0.87442027879477, 0.88013212606195, 0.885430758953404, 0.890301780121058, 
    0.895574751831779, 0.901017998337048, 0.905234482724332, 
    0.91019092788919, 0.914859614014888, 0.9192225506837, 0.923550616805455, 
    0.92771334200536, 0.931595865140241, 0.935445656517242, 
    0.939351401525166, 0.943167085680158, 0.946590824157712, 
    0.950234052029279, 0.953642179398619, 0.957154398608781, 
    0.96040513086275, 0.963813192372516, 0.966837611221, 0.969864120727595, 
    0.972947259751321, 0.975804723219217, 0.978671975521405, 
    0.981565857326285, 0.984255061716605, 0.986910676582415, 
    0.989462665025746, 0.991943061305174, 0.994325593600446, 
    0.996674762755693, 0.998901597809231,
  0.999096386336031, 0.997248719705735, 0.995336590287022, 0.993345931521051, 
    0.991301559485817, 0.989132530523894, 0.986972109141045, 
    0.98474306297177, 0.982338119633783, 0.980008738647176, 
    0.977624406781224, 0.974982586213337, 0.97237885732136, 
    0.969666100173655, 0.966967112745809, 0.964150080806941, 
    0.961239680162186, 0.958459912369279, 0.955205668314446, 
    0.952286431178852, 0.948891863532219, 0.945786430673317, 
    0.942475190084452, 0.938947655714815, 0.93547853673802, 
    0.931752667895925, 0.927880151046155, 0.923919141886397, 
    0.920168804549142, 0.915667485735793, 0.911820509206031, 
    0.90690229009796, 0.902389902871381, 0.897999424111815, 
    0.893216313580705, 0.88829623164542, 0.882912922066582, 
    0.877650666713212, 0.872197286861368, 0.865802159640854, 
    0.860378562461711, 0.854007436314298, 0.847574088986958, 
    0.841231981686811, 0.83444173118948, 0.827591201538672, 
    0.820051667396059, 0.81307739705966, 0.805210009649852, 
    0.796643702248915, 0.788160715083668, 0.779264690303372, 
    0.771515968741643, 0.760307802854106, 0.751302941310739, 
    0.740347542968712, 0.731046789543833, 0.719778931775223, 
    0.707965334587236, 0.694755763883343, 0.683747723210442, 
    0.669781583650596, 0.657019926013976, 0.644048454863421, 
    0.629158837430921, 0.613365781517955, 0.598098453148183, 
    0.58352551040502, 0.565401270310945, 0.548105205639679, 
    0.531314587217963, 0.512510110883474, 0.49382118869888, 
    0.473252601139053, 0.452637572795343, 0.432420548651418, 
    0.411166625708033, 0.390304503487523, 0.36536075202137, 
    0.344824607591489, 0.322857149977263, 0.297816277175968, 
    0.275276728515006, 0.25315581013973, 0.228184057880866, 
    0.205833454423338, 0.181789902744052, 0.162628713236936, 
    0.138683742187767, 0.117728634516661, 0.0980849378527524, 
    0.0818064825141491, 0.0635093187987495, 0.0481159389935149, 
    0.0351678248110907, 0.0233744169126689, 0.014221186033705, 
    0.00764736135247905, 0.00279709369991324, 0.000260157792099835, 
    0.00029305487130239, 0.002630267972568, 0.00752188139060934, 
    0.0143945018212351, 0.0237817389737315, 0.0352757058654693, 
    0.0480516358138974, 0.0643072046153464, 0.0803677401282377, 
    0.0987957455528354, 0.119846860632393, 0.139755345312363, 
    0.16053041049196, 0.18363421783791, 0.204868428424458, 0.226596402526406, 
    0.250141256565284, 0.274195171766261, 0.297343120804141, 
    0.321441150997402, 0.344197203410878, 0.364771431103224, 
    0.388362676208601, 0.412449903405722, 0.433038274251586, 
    0.453049385116054, 0.471922551576142, 0.49315361751497, 
    0.512855463951804, 0.53110887136747, 0.548095005503688, 
    0.565238644449871, 0.582028425353124, 0.59791104182462, 0.61494330480054, 
    0.627754025254362, 0.64260378017244, 0.656794660518141, 
    0.670425385554236, 0.684519654374114, 0.695537303705836, 
    0.707338372003037, 0.720551002591844, 0.730533451774626, 
    0.740942286130072, 0.751341430789751, 0.760434281560887, 
    0.770315855813676, 0.77917362901376, 0.789020462562655, 
    0.796600520347006, 0.804908821488832, 0.812617256192862, 
    0.819759575800869, 0.82775936773495, 0.834466461213194, 
    0.841761534748407, 0.847560742452836, 0.854023526140034, 
    0.860507084716184, 0.866530001790141, 0.872039894391187, 
    0.877846443922768, 0.882899670563553, 0.887683934108601, 
    0.893044818095576, 0.897772944104695, 0.902613818687646, 
    0.906928972729799, 0.911568339544831, 0.915770872474195, 
    0.920001197132769, 0.923985755076171, 0.927921356904989, 
    0.931694644315096, 0.935354466732695, 0.938884827331407, 
    0.942164591110615, 0.945864973873913, 0.949119073987958, 
    0.952219464774281, 0.955346133236671, 0.958414257397861, 
    0.961396069532391, 0.964225805111823, 0.967067792452486, 
    0.969707551442567, 0.972410196467178, 0.975084158505581, 
    0.977422322527534, 0.979966905567048, 0.982429828974745, 
    0.984674860301032, 0.986963202423196, 0.989161557101146, 
    0.991277027826559, 0.993329840765105, 0.995345562914318, 
    0.997250860150465, 0.999091465083693,
  0.999225053475532, 0.997661070878073, 0.996031016491253, 0.994344654299014, 
    0.992581385967659, 0.990767686772001, 0.988894495943554, 
    0.986969108453899, 0.98498227384871, 0.982895872966238, 
    0.980851856740909, 0.978670120523833, 0.976429687224343, 
    0.974114276983188, 0.971936246816699, 0.969297417594975, 
    0.966962299251645, 0.964452080607788, 0.961689849193037, 
    0.958830018427333, 0.956355809946042, 0.95342692546526, 
    0.950333556125921, 0.947344690116889, 0.944055531321466, 
    0.940967955193819, 0.937709969562842, 0.93437183531219, 
    0.930705371291828, 0.926778453245114, 0.923318004563025, 
    0.91915469372285, 0.915496107579367, 0.911371768258761, 
    0.907039786264048, 0.902657173805789, 0.897734889447773, 
    0.893167602040174, 0.888219793958491, 0.88329612896224, 0.87781801264874, 
    0.872586787053267, 0.866396825187987, 0.860120484788229, 
    0.854386448970186, 0.848513055579539, 0.841630756796809, 
    0.834531446219084, 0.827165401055634, 0.820028468611842, 
    0.812238655889825, 0.80397069986332, 0.796458651553578, 
    0.786501819111345, 0.778684505025736, 0.76846741116606, 
    0.757485788317233, 0.748533532169104, 0.737629930752212, 
    0.725959839400793, 0.714839210710246, 0.701612221548224, 
    0.690637041959969, 0.676477593437099, 0.662971714090097, 
    0.647327193977354, 0.632745761482111, 0.617476037669569, 
    0.600745334339147, 0.58497295836845, 0.566218231906097, 
    0.549001067486319, 0.528576815608727, 0.511451738327976, 
    0.487253009734777, 0.468149741878839, 0.445102955752263, 
    0.425082751725054, 0.403022240214376, 0.378314712101912, 
    0.353546803950659, 0.328189722285688, 0.306773304186924, 
    0.280032311933331, 0.255426594905292, 0.229768572455311, 
    0.204474945164455, 0.181643171888788, 0.156713375309216, 
    0.134886680615878, 0.112523630500355, 0.0911024144414605, 
    0.0732823111756263, 0.0567160625977494, 0.0406139823583485, 
    0.0282547899516449, 0.0166073836158078, 0.00827698940703026, 
    0.00316333024876121, 0.000416670036749072, 0.000409139603770569, 
    0.0032046637093002, 0.00850934034244689, 0.0162530985217861, 
    0.0266757248446504, 0.0403220205102863, 0.0562652887478083, 
    0.0729656158357921, 0.0914775628026107, 0.112794509103454, 
    0.136038124030853, 0.156633991658623, 0.180326336877182, 
    0.204725020152059, 0.229810672817692, 0.256642220049274, 
    0.280878191941152, 0.303798755102426, 0.32969793271688, 
    0.353601562887507, 0.376398289176845, 0.40045424469285, 
    0.425706323520315, 0.447491869461377, 0.468901462349868, 
    0.489800115507529, 0.50861260972565, 0.530975813136521, 
    0.547923331008237, 0.566292903882429, 0.583707098835576, 
    0.60176485369425, 0.61717893939474, 0.633386811067284, 0.649086915996787, 
    0.662580082300176, 0.67605566462064, 0.688853919345827, 
    0.702435275232414, 0.714937973694406, 0.726803693650319, 
    0.737351014289467, 0.748653421884862, 0.758670624129419, 
    0.769002553143734, 0.779088569719189, 0.786953086727781, 
    0.795530365447374, 0.804553421457494, 0.812670138395229, 
    0.819794720722114, 0.827293396121113, 0.834377217050674, 
    0.842037882770417, 0.848645830520802, 0.854585559472507, 
    0.860632436187332, 0.865898382366025, 0.872175109062718, 
    0.877965505313886, 0.882937181907143, 0.888370037841274, 
    0.892877464448169, 0.897891085544385, 0.902429690246376, 
    0.906739264614968, 0.911292860248461, 0.9151561200343, 0.91903968454319, 
    0.923312890728908, 0.927166181445121, 0.930622206004617, 
    0.934299836568759, 0.937689341781325, 0.941020062967474, 
    0.944042642615947, 0.947311438975909, 0.950209728821425, 
    0.953308960464558, 0.956225051505776, 0.959231501729177, 
    0.961516707668639, 0.964375962146893, 0.966787436290518, 
    0.969401303726138, 0.971848149049499, 0.974140241090633, 
    0.976554990519584, 0.97861069601356, 0.980778390347582, 
    0.982920570809113, 0.984983796466624, 0.986973505028751, 
    0.988859930000853, 0.990745804881192, 0.992581060874908, 
    0.994324981254073, 0.996040453799765, 0.997651882826916, 0.999225631165327,
  0.999325191133185, 0.997959971206817, 0.996545009352335, 0.995067498855179, 
    0.993557938884241, 0.99197908703488, 0.990333428550764, 
    0.988625382748517, 0.986953417220766, 0.985145956280023, 
    0.983296494175784, 0.981491786296862, 0.97941040884984, 
    0.977454780690364, 0.97543873789271, 0.973276624043817, 
    0.971073109546047, 0.968808403217121, 0.96653968258304, 
    0.964072898820285, 0.961527309768856, 0.959224920267265, 
    0.956375660099636, 0.953837567512599, 0.951096518068303, 
    0.948220901179321, 0.945168086280709, 0.942060443245833, 
    0.938966701750235, 0.935784263699093, 0.932533334990639, 
    0.928936925249494, 0.925153434213716, 0.92161433998919, 
    0.917855258480133, 0.913633576887538, 0.909832894565513, 
    0.905339707389178, 0.900747489149007, 0.896240957592231, 
    0.891388341477318, 0.886506467149822, 0.881388835864116, 
    0.875766694845289, 0.870289781676703, 0.864821278058506, 
    0.859076116581783, 0.852155423242305, 0.84550629944939, 
    0.838578545993551, 0.832469669763405, 0.82398768620635, 
    0.816840968573051, 0.808191492861431, 0.799848383777265, 
    0.79098803763056, 0.781658310725312, 0.772758483660887, 0.76206001480879, 
    0.752051023321047, 0.739746865309026, 0.729819889463929, 
    0.717611962952242, 0.703927361577621, 0.69168545059798, 
    0.678046485654464, 0.662560294334, 0.647244179989643, 0.632451918131306, 
    0.615903690262198, 0.599031150213653, 0.580956334523164, 
    0.562371694179413, 0.541275908104256, 0.521660629197763, 
    0.501704626732817, 0.477600886553868, 0.457153107663456, 
    0.432993619641428, 0.407856186531981, 0.3845476762255, 0.360245642491092, 
    0.333358893018564, 0.307515442754483, 0.280549443484659, 
    0.25335956783031, 0.229227158393316, 0.201709917110489, 
    0.174731619009002, 0.14924687713199, 0.124656527136514, 
    0.104700651890074, 0.0827438121961541, 0.0631928433742707, 
    0.0461471261552441, 0.0308624461396743, 0.0195710684489054, 
    0.00936239853986585, 0.00359709172954459, 0.000487752762393072, 
    0.000473151004262376, 0.00354571004904306, 0.00992450622711253, 
    0.0196510434230395, 0.0317844507760946, 0.0457421232404903, 
    0.0636771702368584, 0.0824965703242619, 0.103271601681857, 
    0.124517404771632, 0.148884154666996, 0.17505302646864, 
    0.199660032333378, 0.226136937805156, 0.253620286238737, 
    0.280928789789837, 0.306578284525561, 0.334134517740212, 
    0.357894731895361, 0.385466464637613, 0.406837531711567, 
    0.432125549989518, 0.455589266536104, 0.477111748745087, 
    0.501198238958689, 0.523103419851748, 0.541686656152131, 
    0.56092729633486, 0.58083657595368, 0.597721224276537, 0.616349296801723, 
    0.632653988508088, 0.648920527471153, 0.663410283872762, 
    0.67886846573778, 0.690621048331742, 0.704986034374847, 
    0.716806903798795, 0.728013624747961, 0.740572318494357, 
    0.75088172748798, 0.762550292163567, 0.771756804006788, 
    0.782097189750556, 0.791331145809204, 0.800536099343564, 
    0.808265255910429, 0.81647467025186, 0.823953555497471, 
    0.831227554408769, 0.839292191046754, 0.846004691180169, 
    0.852429856826439, 0.858499390229735, 0.864430678370798, 
    0.870185587942319, 0.876268406249984, 0.881190839376933, 
    0.886581786952865, 0.891201648500624, 0.896533530135128, 
    0.900844408027468, 0.904975911748333, 0.909700716184238, 
    0.91389209136978, 0.917508689791649, 0.921784965510292, 
    0.925365049141592, 0.928710544617015, 0.932317484779666, 
    0.935627243334693, 0.938685301174429, 0.942105409504087, 
    0.945468375983001, 0.947994094970816, 0.951190576593789, 
    0.953768411941747, 0.956596191550296, 0.959287705436385, 
    0.961597097946996, 0.964093588918851, 0.966456802255174, 
    0.968944101986825, 0.971229852320402, 0.973259466726509, 
    0.975478211113115, 0.977504617206848, 0.979455459418007, 
    0.981452180064002, 0.983291940147442, 0.985182005289769, 
    0.986898455415241, 0.988626161123298, 0.990329976839967, 
    0.991976094392946, 0.993544467696033, 0.995066281172367, 
    0.996539488938722, 0.997956728980933, 0.999322652451704,
  0.999401681446108, 0.998196357625579, 0.99693988038956, 0.995639609749115, 
    0.994290639804333, 0.992921120645425, 0.991469573903631, 
    0.989989505458044, 0.988484935176767, 0.986851575354239, 
    0.985237488664802, 0.983576957502617, 0.981779038019016, 
    0.980086261888638, 0.978271226651035, 0.976356213223139, 
    0.974391635426275, 0.972350879808032, 0.970346765971636, 
    0.968102009373793, 0.965894149871618, 0.963814895620497, 
    0.961372645430722, 0.958849983286016, 0.956450223153517, 
    0.953777958709617, 0.951214687631169, 0.948355397223593, 
    0.945561612452993, 0.942550738391183, 0.939640566288537, 
    0.936421576841007, 0.933124603546232, 0.930011214398361, 
    0.926153188113285, 0.922673215713171, 0.919004497912475, 
    0.915162541120376, 0.910813544535093, 0.906691593237808, 
    0.902636603296318, 0.897963620848334, 0.893388398016363, 
    0.888137580750827, 0.88313433765777, 0.877885523451273, 
    0.872195852631643, 0.866851267847907, 0.860259365306843, 
    0.853978483917244, 0.847408417349041, 0.840837536532036, 
    0.833305436754504, 0.826053536651937, 0.817817670387501, 
    0.809713588391443, 0.80096261181025, 0.791536551652101, 
    0.782389838521687, 0.773122920744277, 0.762049027120479, 
    0.751729995990308, 0.739902569234195, 0.728041989508036, 
    0.715380997677559, 0.702338148691922, 0.688499457517361, 
    0.672897442773021, 0.658521196869367, 0.6415620313158, 0.626416763218687, 
    0.609694722992481, 0.589683327066807, 0.569955212356602, 
    0.550562702428218, 0.528498725639773, 0.50713699147899, 
    0.485588957139066, 0.461597342532412, 0.437006672689333, 
    0.411593353377869, 0.387003606102103, 0.359918652493706, 
    0.331456092262702, 0.304734273109642, 0.277022753247281, 
    0.248642104169652, 0.21961369713169, 0.192947645357843, 
    0.165375839093002, 0.139060914084237, 0.114061864060696, 
    0.0909150302302075, 0.0708334560395052, 0.0517437538905028, 
    0.0354504240300702, 0.0219109775091991, 0.0103921864579152, 
    0.0042968363348528, 0.000491945234003377, 0.000503395016585338, 
    0.00418977956729249, 0.0103214624208384, 0.0216881886308747, 
    0.0349358247103771, 0.0514564533596203, 0.0712362615966918, 
    0.0911766746025369, 0.112967605878911, 0.139279738577513, 
    0.164358629167006, 0.193484196044875, 0.22047447947666, 
    0.248095494782922, 0.277458304598493, 0.305767395696139, 
    0.33253199274061, 0.358426099511018, 0.385848210624282, 
    0.412028433617835, 0.435925443816548, 0.461308339624467, 
    0.485237145809912, 0.508191614627101, 0.528298186356544, 
    0.55042102449476, 0.570003098291472, 0.589877312883371, 
    0.608083044078536, 0.6257120524345, 0.643156953393799, 0.658426120861637, 
    0.674131955959028, 0.688465570058219, 0.702717401205915, 
    0.71643683853439, 0.727687059828177, 0.740547523630387, 
    0.751511279809722, 0.763669915713313, 0.772132714984115, 
    0.782846979674917, 0.79224642680954, 0.801273899185625, 0.80954664017127, 
    0.81816352983057, 0.825844307411249, 0.83317451027145, 0.840275669262587, 
    0.847748616353196, 0.854121269547367, 0.860502502497907, 
    0.866443524678405, 0.872013305263532, 0.877518865075737, 
    0.882897495404425, 0.888297788835002, 0.893463023929235, 
    0.897741987268209, 0.902013442335388, 0.906733005515611, 
    0.911003824768756, 0.914784161774274, 0.919123246895613, 
    0.922803974592148, 0.926544375853471, 0.929865287477201, 
    0.933122571312146, 0.936362594079076, 0.939550965626181, 
    0.942899142215452, 0.945658198908642, 0.948284947353666, 
    0.951297101185768, 0.953823512989744, 0.956579290427724, 
    0.959023853567236, 0.961318940701502, 0.96357594414842, 
    0.965931015046381, 0.968121296433947, 0.970225626463391, 
    0.972352567689223, 0.974405420215758, 0.97625832538395, 
    0.978252278344766, 0.98008324624318, 0.981732985475452, 
    0.983581606762626, 0.98522829760313, 0.986841018845005, 
    0.988482531381353, 0.990002227251741, 0.991469864238436, 
    0.992922786031215, 0.994291722463167, 0.995640684717162, 
    0.996943945739272, 0.998194630867356, 0.999400912554302,
  0.999511555597172, 0.998530471198875, 0.997514918510425, 0.9964785441698, 
    0.995371330127478, 0.994231067187108, 0.993062687961038, 
    0.991880508071866, 0.990621227001225, 0.989341190007835, 
    0.988050947264536, 0.986637168549056, 0.985204682099716, 
    0.983795434001956, 0.982253198923467, 0.980847134569711, 
    0.979137927779963, 0.977482125802053, 0.975803556230993, 
    0.974003705067804, 0.972243263340927, 0.970358618291619, 
    0.968391718190155, 0.966404822216143, 0.964306933114142, 
    0.962284012487882, 0.959956296207302, 0.957616962538758, 
    0.95527091275642, 0.952914642732446, 0.950318053332808, 0.947778500862, 
    0.944987564112738, 0.941945549209709, 0.93929390464931, 
    0.935963276885362, 0.932750783233445, 0.929675100557218, 
    0.926014338450585, 0.92249368991809, 0.91918575737551, 0.914760767473221, 
    0.911377192121115, 0.906900117613279, 0.90259543248925, 
    0.898059388070929, 0.893101125276603, 0.888256521567095, 
    0.883391938068884, 0.877476086168226, 0.871881535620955, 
    0.86584634927612, 0.859813867805626, 0.852307740776201, 
    0.845676821339547, 0.838733097311117, 0.830688362215207, 
    0.823165935829422, 0.815015124710327, 0.806437133530777, 
    0.796236116198785, 0.787581404100709, 0.776485196514998, 
    0.766336653018147, 0.754513065331252, 0.742289077432886, 
    0.729744662627621, 0.715330622524231, 0.702399685410478, 
    0.686851521450439, 0.67171294046127, 0.653817521698609, 
    0.637449819508026, 0.617569515296334, 0.600848082297132, 
    0.578047504518968, 0.5572332908589, 0.536533185657292, 0.510491607004015, 
    0.487170147557164, 0.460934912969355, 0.435953323996151, 
    0.404229720525716, 0.376490045715459, 0.347558758354622, 
    0.317335251683958, 0.286133551568865, 0.255671164550969, 
    0.226025728994494, 0.19462774539296, 0.164221740563476, 
    0.137006920021784, 0.108984903823894, 0.0855740183095384, 
    0.0621795413267412, 0.0423771039668855, 0.0263536042767572, 
    0.0127699405532655, 0.00479366592929175, 0.000530086210127526, 
    0.000512345037934598, 0.00471121567557174, 0.0134708785108288, 
    0.0273244242542281, 0.0422960440884222, 0.0635242860145595, 
    0.083754272696432, 0.10905278981556, 0.137512531556367, 
    0.166127533130336, 0.192603636305045, 0.22356078210125, 
    0.257556576685202, 0.285901591581954, 0.319366580870897, 
    0.348696947747505, 0.377639643049738, 0.407143342274959, 
    0.43398848919732, 0.459808529812245, 0.485838555647771, 
    0.512158528163856, 0.533373931680156, 0.5591589609149, 0.577079759146805, 
    0.599518883668011, 0.619130011966847, 0.636755029979226, 
    0.654204688147436, 0.671234687603053, 0.687053431334011, 
    0.701650385199867, 0.716285269004103, 0.72940544595742, 
    0.742121498806402, 0.754570510050918, 0.76592279756777, 
    0.776612207328873, 0.786445765013737, 0.796638864913239, 
    0.806617472043361, 0.814575800745051, 0.823550514250361, 
    0.831518409500918, 0.838884425032048, 0.846206766904705, 
    0.853139937627567, 0.859931667998949, 0.866389932736602, 
    0.871668501217444, 0.87760345927745, 0.882597918579042, 
    0.888030069333809, 0.892808192842032, 0.897882947078482, 
    0.902616378711633, 0.906958196273796, 0.91104058967038, 
    0.915219019489811, 0.918797603868666, 0.922752292888712, 
    0.926255008336993, 0.930087757162468, 0.93290796079836, 
    0.936301817692619, 0.939179830002915, 0.942139554252361, 
    0.945011107850528, 0.947755407254271, 0.95036186154359, 
    0.952878279063695, 0.955452228131326, 0.957471055485327, 
    0.959965676585688, 0.962350150379015, 0.96431948283707, 
    0.966534119654071, 0.96828550123534, 0.970355691632119, 
    0.972186959166609, 0.973969282109519, 0.975738665295802, 
    0.977508732149986, 0.979129489071271, 0.980648541561997, 
    0.982233335569141, 0.983791875994556, 0.985275043472947, 
    0.986691903544346, 0.988053420072425, 0.989352203675839, 
    0.99062065552392, 0.991859588092555, 0.993062577910144, 
    0.994243154021983, 0.995381918021406, 0.996454113072526, 
    0.997514663084217, 0.998534002418199, 0.99951102855103,
  0.999552556032763, 0.998664237403988, 0.997734052919512, 0.996767605380649, 
    0.995779358147247, 0.994739438958981, 0.993669933931236, 
    0.992590262249443, 0.991411568681888, 0.990256148361176, 
    0.989092819138164, 0.987763923906088, 0.986512607695646, 
    0.985238432933453, 0.98375367626249, 0.98240484508503, 0.980940830792323, 
    0.979361568481206, 0.977821820701579, 0.976283135437828, 
    0.97458309204445, 0.972937632258513, 0.970933645240718, 
    0.969169874239569, 0.96732227487211, 0.965234146257331, 0.96316008285924, 
    0.961260303000261, 0.959139076920285, 0.956902352760269, 
    0.954421934025717, 0.95201569108646, 0.949368124025605, 
    0.946873915731439, 0.944400759209841, 0.941622430637446, 
    0.938532269720793, 0.935340867361241, 0.932009399893178, 
    0.928682112611921, 0.92523190143567, 0.921916641990432, 
    0.918031421536603, 0.914175618823299, 0.909897188246424, 
    0.905726854822336, 0.901343720567198, 0.896421587012845, 
    0.891586204719685, 0.886519157005374, 0.881236901311375, 
    0.876311620923418, 0.869905007308707, 0.863768456208518, 
    0.857262118866135, 0.850189278777757, 0.843281398143493, 
    0.835110170316503, 0.827747726198147, 0.819454469909181, 
    0.810645749442631, 0.801062106850608, 0.791750482435362, 
    0.781081005261728, 0.770208019195686, 0.758010232288088, 
    0.746407207499814, 0.733564268079381, 0.720516544677963, 
    0.705345971811406, 0.690468761538135, 0.674493250668913, 
    0.656145951333807, 0.639170634712597, 0.619841290008341, 
    0.599353295180159, 0.578252881530105, 0.555032273064457, 
    0.531473519144651, 0.507225034127612, 0.479353518809876, 
    0.453781697996496, 0.426992192591972, 0.396264462503104, 
    0.368128806779064, 0.337325650594135, 0.305667772523385, 
    0.272386944211333, 0.240747973864796, 0.209119300532558, 
    0.176740733842632, 0.146703654671055, 0.118649268401476, 
    0.0903146214381478, 0.0666357577747068, 0.0462478164894057, 
    0.0280374695017512, 0.0144122276021484, 0.00587730991054476, 
    0.000651846014758622, 0.000598617332930131, 0.00574112229484655, 
    0.0146590801647587, 0.0277850967471567, 0.0452563208929056, 
    0.0667540519066202, 0.0904403389425741, 0.116915430423038, 
    0.14681219717982, 0.17642263829788, 0.206997281561772, 0.240889903035202, 
    0.273705995075537, 0.306502888921535, 0.33607571809534, 
    0.366238617885336, 0.397336999110125, 0.425689405585357, 
    0.45390544664359, 0.482913160498556, 0.50905961344626, 0.533706104630588, 
    0.555476146745024, 0.578546938147196, 0.600425551294662, 
    0.620176673435056, 0.638865422695121, 0.656951125957899, 
    0.67456778060948, 0.689700153583888, 0.704732660942183, 
    0.719811205573813, 0.733666392595357, 0.745590795865563, 
    0.759233571406526, 0.770703177249962, 0.780789361004097, 
    0.791665454940194, 0.801527906318693, 0.810477280453433, 
    0.818756670185855, 0.827304429528845, 0.835562995399687, 
    0.843207304130485, 0.850376421439691, 0.857431344011066, 
    0.864045205084318, 0.870144342637663, 0.875772803626189, 
    0.881721192059241, 0.886883777366793, 0.891768865670189, 
    0.896431923639634, 0.901183580355801, 0.905941184122293, 
    0.910337950861421, 0.914489835321055, 0.918106221861389, 
    0.921647158492681, 0.925504135267818, 0.928802760155025, 
    0.932335148183069, 0.935321557067216, 0.938418746012833, 
    0.941316178432919, 0.944069014025506, 0.946725652060003, 
    0.949491598895241, 0.952073925760468, 0.954439230631908, 
    0.956965845781433, 0.95909429245794, 0.961093608830369, 
    0.963335435505265, 0.965455622636131, 0.967319237316138, 
    0.96920087770796, 0.971117568235566, 0.972853034944645, 
    0.974604806411347, 0.976278062020964, 0.977912439597297, 
    0.979416230712489, 0.980973024057353, 0.98237066748235, 
    0.983844937345941, 0.985186504598878, 0.986497977432322, 
    0.987814358522261, 0.989064996532264, 0.990282180782801, 
    0.991429527596655, 0.992574623457503, 0.993680817176211, 
    0.99475291480225, 0.995763883408587, 0.996766916078352, 
    0.997736229607611, 0.998658313265702, 0.999552038708569,
  0.999586558160188, 0.998765929399203, 0.997910065838087, 0.997024731182463, 
    0.996101603178214, 0.995152031086055, 0.994172929073752, 
    0.993192472609877, 0.992112783103677, 0.991017392896383, 
    0.989915271583215, 0.988825086629382, 0.987595809806362, 
    0.986426272962975, 0.985151069619223, 0.983741989649964, 
    0.982433166802549, 0.981034602018028, 0.979574280843836, 
    0.978170375252548, 0.976489005593397, 0.9750208483334, 0.97332839020249, 
    0.971602565394141, 0.96988066239882, 0.968022002611769, 0.9660121958982, 
    0.964126877283987, 0.962313542184672, 0.960021345446957, 
    0.957850370826845, 0.955597224968226, 0.953454460493241, 
    0.950864920542217, 0.948516149189442, 0.945680356076154, 
    0.94304138327242, 0.940332611136987, 0.937267877986673, 
    0.934081452278545, 0.930878923446048, 0.927838752623266, 
    0.924365732148819, 0.920686617421787, 0.916761579608172, 
    0.912598417094406, 0.908435728795135, 0.903667238404399, 
    0.899576270492935, 0.894623315534048, 0.889493621385125, 
    0.884381343113333, 0.87864950675275, 0.873043435984157, 0.86705450069689, 
    0.860179119743439, 0.853649227402378, 0.846568266108176, 
    0.838820520855845, 0.83135885665796, 0.821894622620497, 0.81307556557704, 
    0.804395645026032, 0.79488229033762, 0.784175049866593, 
    0.773532127594979, 0.761848442592614, 0.749439302674714, 
    0.735500380632493, 0.722344260516595, 0.706813605707435, 
    0.691633331511653, 0.674828232125846, 0.657058005769118, 
    0.638044376517689, 0.618624385566869, 0.599353579920295, 
    0.575096933043131, 0.552848057474801, 0.527602357220057, 
    0.501906974775652, 0.474247237879724, 0.446875121325636, 
    0.41712470566328, 0.384717713151884, 0.354161921129044, 0.32122599505667, 
    0.288324199630918, 0.255879963227501, 0.221730648477116, 
    0.189664141968571, 0.156173314344004, 0.127688245485291, 
    0.0981757782899249, 0.0720026920637535, 0.049566760412275, 
    0.0303867095011105, 0.0160461014568184, 0.00580970093459081, 
    0.000621384035380759, 0.000715193643010153, 0.00576157271973431, 
    0.0152517484300939, 0.0314273847673242, 0.0507644494623752, 
    0.0718671078802238, 0.0980153951563979, 0.126710839517573, 
    0.156657467914907, 0.189219071124423, 0.222404376906384, 
    0.255870483150484, 0.289185313320123, 0.321035983092349, 
    0.355958679685827, 0.387632328640932, 0.416551356576806, 
    0.447151043000039, 0.475224704162037, 0.502378974414701, 
    0.529027187325386, 0.552919922558784, 0.575434256525435, 
    0.596730651644033, 0.61976155467104, 0.637640076621165, 
    0.658237521462711, 0.67518290727891, 0.692228730690324, 
    0.707060841276468, 0.721344790459159, 0.736019875288166, 
    0.749382260385868, 0.761989803070766, 0.772538406446264, 
    0.784327267705842, 0.794421920060089, 0.804522317993832, 
    0.813544904676425, 0.823248923815225, 0.831544509299746, 
    0.83900053914395, 0.846346527863966, 0.853326527187771, 
    0.860593951049262, 0.86687391499589, 0.872977603488431, 
    0.878980541664682, 0.884461972958719, 0.88967884138462, 
    0.894866190847826, 0.899282141770383, 0.904353740458241, 
    0.908602046297435, 0.912566884478242, 0.916534298171517, 
    0.920386014822974, 0.924171574957428, 0.927468692290413, 
    0.930909870814632, 0.93414756106286, 0.937138668057615, 
    0.940146995793445, 0.942966699876198, 0.945792198523662, 
    0.948240086592505, 0.950768875699028, 0.953229797667574, 
    0.955534482984647, 0.95794663605218, 0.960170789159103, 
    0.962071192849772, 0.964108711221324, 0.966299287179516, 
    0.968051071315541, 0.969918705216317, 0.97165108234553, 
    0.973347188101043, 0.974968740428315, 0.976524559660347, 
    0.97808127443482, 0.979585002497311, 0.981020189091464, 
    0.982431618294111, 0.983746028500883, 0.985099790757343, 
    0.986351317149169, 0.987611453092337, 0.98875789282426, 
    0.989928347550347, 0.991053823928322, 0.9921440751714, 0.993175596422648, 
    0.994187676000341, 0.995158820936158, 0.996105705304883, 
    0.997022557990565, 0.997906055513116, 0.998762507548517, 0.999589157697216,
  0.999641498919789, 0.998928851706107, 0.998198075436508, 0.997434896838605, 
    0.996641954116397, 0.995819324598597, 0.99498435390972, 
    0.994094102984598, 0.99319760810178, 0.992272978450407, 
    0.991310211780352, 0.99034052482914, 0.989258734723814, 
    0.988221767734635, 0.98714366141142, 0.985997782912717, 
    0.984792752153367, 0.983660687979417, 0.982370644812787, 
    0.980996231935074, 0.979697939484052, 0.978404485035343, 
    0.976916524372817, 0.975364475330184, 0.973927806586021, 
    0.972289536454383, 0.970720133097775, 0.969038119364594, 
    0.967237581912117, 0.965549254323153, 0.963588861395666, 
    0.961441838562987, 0.959559119472832, 0.957204351744494, 
    0.955143556385223, 0.952871266668625, 0.950451346540524, 
    0.94785529105516, 0.945530676004917, 0.942528103122422, 
    0.939574588385084, 0.936932352302386, 0.933887820025724, 
    0.930318064807532, 0.927212240652156, 0.923609380990342, 
    0.920002769096036, 0.915664478242391, 0.912020815421721, 
    0.907828427654825, 0.903336386868047, 0.898764164642312, 
    0.893416080849411, 0.888091033872545, 0.882417801631435, 
    0.877263278268091, 0.870886373632478, 0.864343645711193, 
    0.857480620649671, 0.85039359975844, 0.842264107294384, 
    0.834257886226718, 0.825802696750693, 0.817377150911884, 
    0.80719895173037, 0.797409954320647, 0.787636346204749, 0.77464534461475, 
    0.761886500876789, 0.749379813547301, 0.73693116853895, 
    0.721680059941846, 0.705771785199522, 0.689302986708689, 
    0.669988707368817, 0.651580552385999, 0.632368252639233, 
    0.610876170526999, 0.587905257542861, 0.56464106118381, 
    0.538272208872317, 0.50948723651921, 0.481344358394086, 
    0.450130902542373, 0.420959944287004, 0.387444687557058, 
    0.354022164899428, 0.318945561238459, 0.284104986536803, 
    0.246797534882755, 0.212481290859532, 0.177642257072369, 
    0.142103919424527, 0.11086327487153, 0.0822324416371782, 
    0.0569457252415102, 0.0353013643845588, 0.0178921061854488, 
    0.0063809855963998, 0.000804044588343946, 0.000693029001315955, 
    0.00662022754278715, 0.0181505507179673, 0.034801370548946, 
    0.0572031269314853, 0.0816679322050754, 0.112274247968829, 
    0.141989670231988, 0.176707258293592, 0.211562762878877, 
    0.24686292422278, 0.283622673317714, 0.319262801988025, 
    0.355009664021917, 0.388411409859405, 0.420189213827913, 
    0.453189676739361, 0.479727899349635, 0.509873341932213, 
    0.536973316087847, 0.563272011704384, 0.587246488195438, 
    0.609683285747881, 0.631248922604389, 0.653461243706161, 
    0.670790751421353, 0.689170547614956, 0.705966698313855, 
    0.720638198581117, 0.735849625360921, 0.749431790548346, 
    0.762718008707612, 0.774052517053051, 0.786980578404629, 
    0.797398984252463, 0.807562769630862, 0.816308911284279, 
    0.826362976749969, 0.834430843255487, 0.84285093545578, 
    0.850292156980778, 0.857566407694839, 0.864444828158511, 
    0.870845672110321, 0.87715317468308, 0.8828831759104, 0.888136215524575, 
    0.893380198314355, 0.898498628248392, 0.903614713638076, 
    0.907365653172563, 0.911814148074697, 0.915888682360836, 
    0.919806210175911, 0.923491209818524, 0.927097668212797, 
    0.930440288824319, 0.933899312214747, 0.93677167304582, 0.93993661866745, 
    0.942637970282277, 0.94547977635884, 0.947991765623612, 
    0.950681304474504, 0.952818449084427, 0.955119135509145, 
    0.957444098108374, 0.959531287095747, 0.961465785023939, 
    0.963491337882114, 0.965337037542468, 0.967191844477612, 
    0.968994612433238, 0.970695774405579, 0.972276272109056, 
    0.973889783357661, 0.975475255999946, 0.976933964828134, 
    0.97841881694499, 0.979798810481283, 0.981099882398301, 
    0.982407433257485, 0.98358692057262, 0.984860073973219, 
    0.985968880931549, 0.98709087278558, 0.988192159645307, 
    0.989294668672367, 0.990303803458819, 0.991286272599575, 
    0.992282504861151, 0.993200300773301, 0.994109683281812, 
    0.99498536909867, 0.995815416160705, 0.99665094415861, 0.997423844453339, 
    0.998187750162734, 0.998927594407766, 0.999641678036809,
  0.999684785702764, 0.999057640463813, 0.998403705387892, 0.997740614410753, 
    0.997057675558794, 0.996330981428619, 0.995579820638635, 
    0.994830000456381, 0.994028598797716, 0.9932230591699, 0.992386429514226, 
    0.991502623098097, 0.990626542926452, 0.989660851481749, 
    0.988674085951244, 0.987713750338665, 0.986682528598359, 
    0.985613398256277, 0.984498919606254, 0.983318644956531, 
    0.982201135003489, 0.98101212844083, 0.979723256856011, 
    0.978401878921677, 0.977040040192943, 0.975627284862613, 
    0.974183046804259, 0.972797501921567, 0.971135323093824, 
    0.969539037297683, 0.967774193478124, 0.965999085550136, 
    0.964197287950694, 0.962387759975234, 0.960215162433231, 
    0.958352210914607, 0.956202876943391, 0.953834506864599, 
    0.951793289756909, 0.949117082817865, 0.946592728467793, 
    0.943990921118149, 0.941134466660337, 0.938501771332479, 
    0.93552959991358, 0.93239396657548, 0.928916808220323, 0.925165207193339, 
    0.921671828243458, 0.917706997510946, 0.913693814878176, 
    0.909359330971658, 0.90526906940253, 0.900646580008796, 
    0.895237170421872, 0.890238304472158, 0.8843688524539, 0.878427398738849, 
    0.872477130770962, 0.866387080653873, 0.859239568005662, 
    0.851540313372463, 0.843887078945484, 0.835974888432386, 
    0.826204879362086, 0.816894558525645, 0.807546208233264, 
    0.795791664134495, 0.785028277222824, 0.772803003885339, 
    0.760231181687642, 0.745810548858009, 0.73186010705303, 
    0.714918347322911, 0.697101356706791, 0.681062458886012, 
    0.660974304816937, 0.640965197310791, 0.617439756719093, 
    0.594098646640667, 0.568628781523747, 0.542383335050907, 
    0.513917737434086, 0.483461632605034, 0.450097316154547, 
    0.41741901351711, 0.382519781994107, 0.347322415515192, 
    0.310197014012906, 0.270718487883133, 0.23288110927774, 
    0.196184136272342, 0.160823742506943, 0.122325741550826, 
    0.0938466091377307, 0.0627866556227013, 0.0389535222102849, 
    0.0202972723591231, 0.00758506038099968, 0.000937059190545454, 
    0.000851444929450195, 0.00786970583223504, 0.0206749040752202, 
    0.0402095289165446, 0.0634820883358193, 0.0919531055233731, 
    0.12434967280517, 0.158754441371951, 0.195747481576604, 0.23270109457117, 
    0.272705375937607, 0.309533123515114, 0.346329688733236, 
    0.383381910095993, 0.418582038509166, 0.450633846990409, 
    0.484189695760135, 0.512130817305172, 0.542600826949863, 
    0.568396106777548, 0.592992411733701, 0.61787575291912, 
    0.639565012517507, 0.660733870694876, 0.680061440289097, 
    0.698274131074342, 0.715090782266247, 0.73240272960282, 0.74667942873915, 
    0.759849308363716, 0.772663101926145, 0.784789226614044, 
    0.79679781530802, 0.8069414054707, 0.816538400612277, 0.826485308830482, 
    0.835096197211827, 0.843292674065345, 0.851034454162721, 
    0.859206263581404, 0.86611338178357, 0.872704072446011, 
    0.878646990404737, 0.884469747496936, 0.889948898502895, 
    0.895264723580068, 0.900332021781976, 0.904998902935141, 
    0.909536775373185, 0.913782565995874, 0.917899852775019, 
    0.921686882176889, 0.925628014283565, 0.928607991835006, 
    0.932333972396738, 0.935166780148294, 0.938434929612238, 
    0.941369329289894, 0.943796038547894, 0.946782300044622, 
    0.949343465096961, 0.951680792887117, 0.953994536446067, 
    0.956098026301299, 0.958344944433349, 0.960289047894975, 
    0.96235709777472, 0.964262253564519, 0.966027351355327, 
    0.967665778615557, 0.969495607802767, 0.971163137058894, 
    0.972671627007468, 0.97408149557871, 0.975708324080973, 0.97705010943564, 
    0.978521889654139, 0.979792483614441, 0.981032623073671, 
    0.982193447460636, 0.983309037482177, 0.98448548698028, 
    0.985597620041729, 0.986690637555168, 0.987675157185679, 
    0.98872614812811, 0.989694494621027, 0.990620566543615, 
    0.991518698654776, 0.992367158829835, 0.993226207439359, 
    0.994034726065226, 0.994829207410768, 0.995578247851546, 
    0.996332968680328, 0.997045513070161, 0.997738972763329, 
    0.998409505478076, 0.999062343889637, 0.999685035343276,
  0.999716701576306, 0.999155967322368, 0.998580113753384, 0.997982743045717, 
    0.997375581596014, 0.996722677359579, 0.99605674698873, 
    0.995414821576001, 0.994678440086203, 0.993957631125354, 
    0.993206768847996, 0.992402461777497, 0.991597888031457, 
    0.990781672309437, 0.989928147497282, 0.989004608169651, 
    0.988116705420429, 0.987148252600572, 0.98621941358529, 
    0.985157188817154, 0.984066952464678, 0.983032907558304, 
    0.981901357622653, 0.980757816501025, 0.979538546584727, 
    0.978311967745566, 0.976989077444051, 0.975551483827848, 
    0.974161233259438, 0.972740565531088, 0.971173764528019, 
    0.969587379564867, 0.96808460988693, 0.966376657045013, 0.96451703759326, 
    0.962662035547796, 0.960854328352722, 0.958699267475326, 
    0.95674450541666, 0.954435301912407, 0.952149977036773, 
    0.949764962792036, 0.947228757498362, 0.944603913897756, 
    0.941847805196577, 0.938968540085108, 0.935844222310863, 
    0.932921015101452, 0.929698112728934, 0.925927601453179, 
    0.922169172146554, 0.918529040061211, 0.914253980640565, 
    0.910136420222473, 0.905564836588166, 0.900488190645552, 
    0.89574487577743, 0.890540595159659, 0.884287035136631, 
    0.878654135498766, 0.872416147366452, 0.865074187953089, 
    0.85819658544419, 0.850237825453036, 0.841543765610795, 
    0.833678409606679, 0.823341846416935, 0.813136007133386, 
    0.802688021290855, 0.791243740911662, 0.779692618713679, 
    0.767440984023945, 0.752442083151974, 0.737356755867357, 
    0.720716202026052, 0.703925070441419, 0.685365094850152, 
    0.664715751623147, 0.643557073279478, 0.620976587642904, 
    0.596371696115636, 0.569394551524605, 0.542383686014675, 
    0.511804650716199, 0.478293436750115, 0.44610702530386, 
    0.408550155190651, 0.372648696685601, 0.334197595702763, 
    0.29216285579354, 0.254598466842738, 0.212757844348929, 
    0.174805728404862, 0.139068267863412, 0.101284335200309, 
    0.0701623208486062, 0.0433676352821954, 0.0230688770077151, 
    0.00826615510489354, 0.000862628313351811, 0.000816970216553045, 
    0.00824900775658228, 0.0223075871758849, 0.043931709156172, 
    0.071694348541377, 0.101517889521192, 0.136601395443179, 
    0.174175492685723, 0.213511798116339, 0.253982817010077, 
    0.293330276179029, 0.334775391405517, 0.37126478556414, 
    0.408203330935834, 0.446060789472681, 0.479075688772403, 
    0.511158728100278, 0.540224386921188, 0.566239663158145, 
    0.595422698863591, 0.620403709465654, 0.644815179968758, 
    0.664059396836281, 0.68528230567721, 0.704280503754034, 
    0.720265710581662, 0.736770396129806, 0.752435926841882, 
    0.766473705760969, 0.780064375118811, 0.791971912725755, 
    0.803578721014676, 0.813725796746732, 0.82385045396431, 
    0.833157911963059, 0.841113104116475, 0.849519504782995, 
    0.857701231804319, 0.864894823859029, 0.871722711764083, 
    0.87859907002506, 0.884594064425965, 0.890202015874039, 
    0.895326537000249, 0.901092014899778, 0.905383478721901, 
    0.909920225267102, 0.914527535065426, 0.918128526817571, 
    0.922410379750883, 0.925869174336237, 0.929491059788781, 
    0.933053072854465, 0.936070565981635, 0.939021087590308, 
    0.941929990927247, 0.944592472068648, 0.947275310238494, 
    0.949823881270189, 0.952262843168138, 0.954462543266435, 
    0.956584071738911, 0.95864708968772, 0.960884629779989, 
    0.962638736468296, 0.964445193882513, 0.966184332859442, 
    0.967959561904257, 0.969696674736533, 0.971110750842712, 
    0.972643217021123, 0.974247717840069, 0.975626325361495, 
    0.976914442579653, 0.978251608310982, 0.979476386753499, 
    0.980691481106043, 0.981914034858524, 0.982967951422977, 
    0.984083625080935, 0.985125946278741, 0.9862113705085, 0.987209412489685, 
    0.988153069149822, 0.989043333769923, 0.989913337497325, 
    0.990747991223311, 0.991598501785933, 0.992415331947024, 
    0.993216564382322, 0.99394999417832, 0.994673919429863, 
    0.995359405544305, 0.996068640696288, 0.996724117673852, 
    0.997363668755621, 0.997984891601347, 0.998581772078221, 
    0.999159494774627, 0.999717272562097,
  0.999745056758972, 0.999239782321485, 0.998722676895225, 0.998182426258991, 
    0.997617954456703, 0.997056593338915, 0.996458844048359, 
    0.995842083206856, 0.995214404091863, 0.994535770402685, 
    0.993871739081546, 0.99314680516298, 0.992418574817361, 
    0.991661305520832, 0.990901240327081, 0.990112856701659, 
    0.989249101700193, 0.988429506673276, 0.987536493772015, 
    0.98661778199578, 0.985651062965257, 0.984627127210279, 
    0.983605961536722, 0.982629882738158, 0.981494503376625, 
    0.980401167586432, 0.979190133300797, 0.977956880245007, 
    0.976681469821708, 0.975438126737008, 0.973992759776283, 
    0.972469465254578, 0.971050483325796, 0.969568169292063, 
    0.967951440674314, 0.96610337914766, 0.964490875167232, 
    0.962704967112666, 0.960713074036862, 0.958687218458989, 
    0.956606575769934, 0.95443733931172, 0.952269116396355, 
    0.949788664314029, 0.947242400593532, 0.944642957951843, 
    0.941804223179538, 0.939217650220746, 0.935830246863021, 
    0.932639507085029, 0.929352853687179, 0.925949548041357, 
    0.921837764558206, 0.917934742566324, 0.913899100287094, 
    0.909486341819303, 0.904563116074557, 0.899660798364644, 
    0.894574630589329, 0.889210122802296, 0.88298242971215, 0.87656046256033, 
    0.870056916997657, 0.863236681729992, 0.854402263730829, 
    0.846956682245969, 0.838610631332931, 0.829201492206559, 
    0.818411277206575, 0.808829448391153, 0.795753056212234, 
    0.783882956456405, 0.770658618534656, 0.755704914790809, 
    0.741704218214145, 0.724548045287491, 0.707042458260291, 
    0.687735014246038, 0.667354253772731, 0.644451923372162, 
    0.618896886160335, 0.596150380358236, 0.566964223076232, 
    0.535554036159635, 0.503345736953625, 0.470969262837178, 
    0.433515341336778, 0.396698498947303, 0.356227700931172, 
    0.315530665749245, 0.275266820524516, 0.229584634772837, 
    0.187663444358651, 0.148469553489207, 0.11220031987249, 
    0.0779082221313826, 0.0482478616994463, 0.0252745135723694, 
    0.00935071915915743, 0.00102284674660367, 0.00110564220549593, 
    0.00949599584300527, 0.0256274152267887, 0.0482640359992445, 
    0.0773688305826944, 0.112357851363557, 0.150930952395744, 
    0.189487245552967, 0.231714779947021, 0.272982842432727, 
    0.316205781069247, 0.356410643296211, 0.395583813527103, 
    0.434380856300395, 0.469010961424327, 0.504711814125009, 
    0.535105915491432, 0.565914461167236, 0.594368279830139, 
    0.619961856631762, 0.644793359283316, 0.666438224308853, 
    0.687852843698647, 0.706099928944301, 0.723962830896769, 
    0.742067482744319, 0.755979802294334, 0.770796857390187, 
    0.783660232261301, 0.796629973393682, 0.808038609275009, 
    0.818410552585796, 0.828390654941281, 0.838570434046366, 
    0.847029885040728, 0.854993619711817, 0.862611033754936, 
    0.870215994606712, 0.876689720508755, 0.882944166374794, 
    0.888418443421338, 0.894462333269211, 0.899833444386805, 
    0.904551022431704, 0.909441136474112, 0.913605304962935, 
    0.917764723603541, 0.921737257298923, 0.925842764099254, 
    0.929295097296953, 0.932520330648682, 0.935910807422742, 
    0.938981702232376, 0.941756959226911, 0.944853689772466, 
    0.947246565584667, 0.94979154029304, 0.952099424271745, 
    0.954326305498788, 0.956579014292898, 0.958627780613742, 
    0.960824143553944, 0.962627333636993, 0.964426469631545, 
    0.966293796191603, 0.967894360950865, 0.969565926788519, 
    0.970997370748774, 0.972493068991015, 0.973910113600346, 
    0.975385099574866, 0.976737104427774, 0.977960751255974, 
    0.979124331931443, 0.980378070926626, 0.98144412856829, 
    0.982587662004958, 0.983615214938399, 0.98464630527738, 
    0.985716683749416, 0.986617155932202, 0.987490896830045, 
    0.988418920926958, 0.989235744582863, 0.990090483144911, 
    0.990883465858961, 0.991675697898346, 0.992445828282869, 
    0.993171208129478, 0.993869611890549, 0.994555271246258, 
    0.995205436356245, 0.995831735641631, 0.996453321815425, 
    0.997040026474532, 0.9976277744922, 0.99818220526528, 0.998721558745277, 
    0.999240364163306, 0.99974289191095,
  0.999749728256862, 0.999258589825262, 0.998748992013169, 0.998223704116802, 
    0.99767726208251, 0.997109436037908, 0.996527349188895, 
    0.995948870882216, 0.995332779717778, 0.994676602007682, 
    0.994026003606772, 0.993305338528606, 0.992602085671751, 
    0.991887606530744, 0.991110284302859, 0.990346670267085, 
    0.98956914137476, 0.98873235200515, 0.987826112820402, 0.986906663444151, 
    0.985935580114485, 0.985051362217822, 0.984054025108515, 
    0.982992038383354, 0.981959935048972, 0.98084778008311, 
    0.979535307441172, 0.978460761052229, 0.977208809220423, 
    0.975928645897669, 0.974550645213876, 0.973167048486115, 
    0.971778618487119, 0.970146389705226, 0.968696536528267, 
    0.966992767352426, 0.96527241625155, 0.963443012137933, 
    0.961665863678694, 0.959864506816378, 0.957692472964574, 
    0.955457226330647, 0.953325522716475, 0.950967592892612, 
    0.948279626517884, 0.946008031727249, 0.943133719628415, 
    0.940189833226265, 0.937413415462351, 0.934281989516517, 
    0.931051247021122, 0.927526648107161, 0.923658817782183, 
    0.919650579864043, 0.915393619653839, 0.911350737597871, 
    0.906844762128231, 0.902076292889989, 0.896595000853274, 
    0.891406927900565, 0.88538814764058, 0.878754185687264, 
    0.872948602444952, 0.865191681283119, 0.857668341084436, 
    0.850108463044583, 0.841240875472825, 0.831725228892177, 
    0.822159017398895, 0.811383937384216, 0.800244380889623, 
    0.787908448840651, 0.775148329461496, 0.761144926391284, 
    0.745788724242636, 0.729036504881457, 0.71240221534712, 
    0.692649648050276, 0.6722177182108, 0.649429814002617, 0.624819710427854, 
    0.598300130365538, 0.571772396274124, 0.540002848731839, 
    0.511961876701559, 0.475559718834913, 0.438867219791746, 
    0.402922270858304, 0.361542071565656, 0.321085224750741, 
    0.278324714515694, 0.236832335469908, 0.193790089441213, 
    0.153492330006324, 0.113605894471238, 0.07969878971358, 
    0.0504080488002694, 0.0253714538662893, 0.00936542208992971, 
    0.00103848061847609, 0.00118168642981441, 0.00931884588419745, 
    0.025972220036343, 0.0496802030096172, 0.0800051076499589, 
    0.113648383700702, 0.152174589969416, 0.194098575011979, 
    0.236227414281099, 0.277414502346752, 0.322425303223266, 
    0.361264899806123, 0.40226110274495, 0.440212503327497, 
    0.476291074609391, 0.511012857876803, 0.542059161640542, 
    0.570772496136829, 0.599547095018775, 0.625268289262769, 
    0.648899357999573, 0.670850012574007, 0.691097619764652, 
    0.711673393888159, 0.72975007615958, 0.745434184069415, 
    0.761517489984331, 0.77513814903672, 0.788440616928489, 
    0.799698475342775, 0.811873556320753, 0.822282592523055, 
    0.832342792566485, 0.840881696991423, 0.849536205594388, 
    0.857932709247287, 0.865128182153545, 0.872455846592336, 
    0.879344611961607, 0.885557036530687, 0.89087075997929, 
    0.896717392209553, 0.901895893877931, 0.906820736496772, 
    0.91128953617305, 0.915792021058803, 0.920014126268513, 
    0.923857289129562, 0.92737304355264, 0.931025724242832, 
    0.934451834351566, 0.937129064697588, 0.940407326535602, 
    0.943345142621239, 0.945734448202863, 0.948292608689802, 
    0.950764300432951, 0.953159902890643, 0.955417375321919, 
    0.957731701242964, 0.959711783357512, 0.96143928794094, 
    0.963402064693399, 0.965358524163279, 0.966893275998205, 
    0.968559316236298, 0.970236916160505, 0.971636006410224, 
    0.973071275152874, 0.974531448374338, 0.976049936647345, 
    0.977209980156388, 0.978457156642408, 0.979604740092108, 
    0.980871611228634, 0.981890648352094, 0.982975615441496, 
    0.984021452501248, 0.984975646029971, 0.986004939226325, 
    0.986968781787747, 0.98784362044579, 0.988686248381267, 
    0.989508490361821, 0.990334426663781, 0.991136829902235, 
    0.991875376513504, 0.99263712040265, 0.993305742432269, 
    0.994014629958751, 0.994677500569451, 0.995317718349466, 
    0.995937260295239, 0.996531183666525, 0.997111674472876, 
    0.997677619038449, 0.998223459150115, 0.998750232617179, 
    0.999258234075324, 0.999749229617448,
  0.999754615794338, 0.99927577162449, 0.998773525129233, 0.998260297637948, 
    0.997739223168597, 0.997178359053438, 0.996611354520341, 
    0.996025616221107, 0.995429924496558, 0.994802857256655, 
    0.994142434326866, 0.993489820007489, 0.99277423425032, 
    0.992064979342153, 0.991331618699233, 0.990631408280385, 
    0.989729964976427, 0.989012406213694, 0.988084442793767, 
    0.987237633232216, 0.986354154180701, 0.985390455061457, 
    0.984387969420968, 0.983382642335008, 0.9822967268595, 0.981287064864582, 
    0.980085356986551, 0.978981490231773, 0.977794662308997, 
    0.97654815247387, 0.975139641591096, 0.973769605336837, 
    0.972379872982814, 0.970805190114398, 0.969349867463507, 
    0.967736571295498, 0.96617105883226, 0.964363779927639, 
    0.962544940320739, 0.960521994393496, 0.958650026857333, 
    0.956695742276747, 0.954380402743925, 0.951848258765234, 
    0.949407420012358, 0.947027683506959, 0.944457122881116, 
    0.941678440329919, 0.938740828473476, 0.935786137231541, 
    0.932377401619835, 0.92895262386922, 0.925336407106464, 
    0.921444983926673, 0.917501889510062, 0.913085533438791, 
    0.908916650765149, 0.903910665146264, 0.898778220711554, 
    0.89320315855457, 0.88766462768238, 0.881768895419224, 0.874940300457866, 
    0.868379826336684, 0.861209310913739, 0.852790791716183, 
    0.84410008641971, 0.835565885825426, 0.825790974218036, 
    0.815367570412467, 0.804252450751307, 0.791375639225732, 
    0.778851150577334, 0.765486134021974, 0.748689891722588, 
    0.733607899736366, 0.715148658538484, 0.696445367480779, 
    0.67739200459199, 0.654738333645857, 0.630379352183558, 
    0.605436666979198, 0.577518741955491, 0.548113841304892, 
    0.516364188148559, 0.482459262184042, 0.44443216544238, 
    0.407988620279961, 0.36743594220518, 0.3263009247319, 0.283038113231729, 
    0.241789948873217, 0.196162204801886, 0.155478301671026, 
    0.115244128503688, 0.0810328367687401, 0.0499418805792907, 
    0.0262029151076208, 0.00977253884735651, 0.00101820694859385, 
    0.00105838006997085, 0.00977883040695859, 0.0263187850247883, 
    0.0511910857306298, 0.0805304351115091, 0.11658682177036, 
    0.15505558628633, 0.197403062694529, 0.240206614715953, 
    0.282322330580854, 0.324532427243793, 0.366597012822122, 
    0.40791322338002, 0.445519592966921, 0.482587072199042, 
    0.516583118492006, 0.548515234547526, 0.577566893634513, 
    0.604946702697276, 0.630422740671034, 0.654459490813352, 
    0.676890573563661, 0.697531112732869, 0.716496007513551, 
    0.733809753302004, 0.750173354265828, 0.764085608836087, 
    0.778978035887011, 0.791442121615499, 0.804077501899613, 
    0.815599462794571, 0.825787989496467, 0.83561731752793, 
    0.844041816318981, 0.852617390414055, 0.86082155665642, 
    0.868353982756975, 0.874870603141658, 0.881668384871959, 
    0.887497214170589, 0.893509084409306, 0.898651790781539, 
    0.903724542393177, 0.908606440818681, 0.913263163499301, 
    0.917744783503842, 0.921553357592322, 0.925606378645456, 
    0.929046798504823, 0.93234905276972, 0.935616509286501, 
    0.938644911649004, 0.94161084202438, 0.944397368746958, 0.94717747073039, 
    0.949416424405087, 0.951982505144317, 0.95447563374935, 
    0.956442335499092, 0.958355053543943, 0.960574948626566, 
    0.962496356336443, 0.964227480906813, 0.96604699409729, 
    0.967675949183686, 0.969364501004265, 0.970941516336677, 
    0.972369927893304, 0.97377416144037, 0.97511117879222, 0.976550809290422, 
    0.977737794939871, 0.97890270849027, 0.98008411374248, 0.981258773286364, 
    0.982291600355259, 0.983393334889097, 0.98440355032813, 
    0.985384346491522, 0.986258063385462, 0.987272427914515, 
    0.988095235885627, 0.988972202045963, 0.989739607331163, 
    0.990599305111881, 0.991290397779312, 0.992068162520858, 
    0.992777312243214, 0.993472232660357, 0.994156256413526, 
    0.994796893727907, 0.995425223214302, 0.996027977485068, 
    0.996625167880742, 0.997183655461356, 0.997734449882112, 
    0.998269617588451, 0.998776997407467, 0.999278278697531, 0.999755391479848,
  0.99976673428062, 0.99930559623191, 0.998831689477739, 0.998346419089402, 
    0.997841834782092, 0.997312837289353, 0.996762903593534, 
    0.99620365048507, 0.995629050542641, 0.995041099541048, 
    0.994410594726201, 0.993771468279849, 0.993099184270033, 
    0.99240926588464, 0.991712049981225, 0.990986912189674, 
    0.990228010301243, 0.989451970574327, 0.988621693156869, 0.9877784642102, 
    0.986917305471706, 0.986012511467412, 0.985040307021778, 
    0.984113892351427, 0.983093862025386, 0.98208712894924, 
    0.980982366273411, 0.979861056974631, 0.978701599049359, 
    0.977504208129299, 0.976314289278007, 0.974972588023441, 
    0.973593267170594, 0.972143578250408, 0.970631067559479, 
    0.969207595346418, 0.967593316940197, 0.965937209435185, 
    0.964029735928439, 0.962120927234346, 0.960442667140555, 
    0.95833547626414, 0.956159551176324, 0.95415003294943, 0.951896358971206, 
    0.949293120077828, 0.946668555487922, 0.944245868013283, 
    0.941288706447497, 0.938404682017817, 0.935175030903398, 
    0.931985672275016, 0.928627833241472, 0.924796118059523, 
    0.92085847012631, 0.916877607446366, 0.913037796017993, 
    0.907777818323743, 0.902716026544023, 0.897402181018452, 
    0.892072426000091, 0.886296390994106, 0.880131454740711, 
    0.873320710656888, 0.865880511934624, 0.857945196696411, 
    0.85023991339563, 0.841406130604323, 0.831607121257559, 
    0.821165456693773, 0.81109508572362, 0.79959124929625, 0.786963877335949, 
    0.773405914166525, 0.758137655190393, 0.741747988061736, 
    0.725195486558481, 0.707131612004459, 0.687470360392035, 
    0.664608639888647, 0.641758121591917, 0.616599879914203, 
    0.588869759354888, 0.559456597153417, 0.527014044588026, 
    0.492388870721759, 0.454931381166354, 0.417986986340384, 
    0.377705754666347, 0.33851495201652, 0.293125442959569, 
    0.247960797066311, 0.204767248398804, 0.161702047297636, 
    0.120671101569895, 0.0833562317679306, 0.0535831929450022, 
    0.0276431545227692, 0.0101213942681174, 0.00114467071742554, 
    0.00103445619155282, 0.0103357168112965, 0.0287305872854773, 
    0.0532294037086977, 0.083659868519079, 0.121233440670671, 
    0.161732401487639, 0.204541804650441, 0.247859750478673, 
    0.291878711109161, 0.33619892649995, 0.378806908599605, 0.41805993520787, 
    0.455322145284171, 0.491231532981761, 0.525908289968927, 
    0.559288229986958, 0.588062237250336, 0.616165322360218, 
    0.641199074133808, 0.664611591202396, 0.685950400297542, 
    0.70660799517541, 0.724039820546518, 0.742251576083357, 
    0.759008584574581, 0.773318992017819, 0.786355305212389, 
    0.799537885261725, 0.810988746929882, 0.821678134393885, 
    0.832083001409703, 0.841381140552576, 0.850143862619286, 
    0.857926740629119, 0.866496657407963, 0.873494585217268, 
    0.879707055297955, 0.885990112320038, 0.89247800262511, 
    0.897575438858186, 0.902829821542182, 0.908098446431471, 
    0.912471881202982, 0.916732706250475, 0.921059854948823, 
    0.924736656634052, 0.928539220089314, 0.932097848936068, 
    0.935245028489836, 0.938535491686779, 0.941120580615206, 
    0.944233371841561, 0.946712244281535, 0.949441930204658, 
    0.951605056985329, 0.953962906180967, 0.956245543806643, 
    0.958254940585544, 0.960380874958454, 0.962279427007092, 
    0.964138996948429, 0.965797789931181, 0.967545531386574, 
    0.969146764285664, 0.970801176735505, 0.972158880696172, 
    0.973481310151345, 0.975024145554748, 0.976148044147384, 
    0.977575784679424, 0.978819278396573, 0.979940767106067, 
    0.98101860156576, 0.982131103666409, 0.98312850487079, 0.984108381844602, 
    0.985132796853215, 0.98608678378803, 0.986912715857179, 
    0.987778660889995, 0.988604396286039, 0.989445170798773, 
    0.990241055572417, 0.99100506084035, 0.991704944227478, 
    0.992415297920824, 0.993116418763443, 0.993791129747842, 
    0.994406330956783, 0.995020460775758, 0.995618113865267, 
    0.996202006023885, 0.996764581124918, 0.9973036079676, 0.997831455519525, 
    0.998342103441473, 0.998832189583407, 0.999309244190239, 0.99976672644068,
  0.999784479224028, 0.999364347024858, 0.998925421709953, 0.998477324902955, 
    0.998015698801182, 0.997534500655101, 0.99702899015647, 0.99651156575347, 
    0.995985382624618, 0.995428006639918, 0.994877623090588, 
    0.994276376445849, 0.993676891733425, 0.993033229365589, 
    0.99240153542025, 0.991713125454777, 0.991017194607951, 
    0.990310970202699, 0.989553367917421, 0.988799826352283, 
    0.987977111211647, 0.987203443677991, 0.98624531176087, 
    0.985413251478204, 0.984501926289147, 0.983594479114347, 
    0.982461575229632, 0.981521446244197, 0.980451972719884, 
    0.979326298797808, 0.978196933271379, 0.977053254490559, 
    0.97563352136175, 0.974341677259021, 0.973100144737026, 0.97173403052913, 
    0.970169944309407, 0.9685691558418, 0.96695110931072, 0.9652880456789, 
    0.963421085528664, 0.961624071863917, 0.959737784047066, 
    0.95759966779102, 0.955580297158202, 0.953313277291769, 
    0.950939648935224, 0.948344486472188, 0.945954663304452, 
    0.943031304609622, 0.94011219236137, 0.937045228030667, 
    0.934142478589239, 0.930520425531468, 0.926915615628321, 
    0.923303555782416, 0.919148012637194, 0.914747014729241, 
    0.910132815576493, 0.905373958987918, 0.89999947118542, 
    0.894343290444669, 0.888815609391203, 0.881878960748415, 
    0.875674134439308, 0.868318669779891, 0.860546224662168, 
    0.852168559047713, 0.843397405863405, 0.833556325138952, 
    0.823765600042655, 0.81260401760796, 0.801263784980834, 
    0.787856230271217, 0.773722481023931, 0.75769768234791, 
    0.741796663064061, 0.723709833622068, 0.703699453633346, 
    0.683334348921845, 0.661078745406871, 0.635657428739632, 
    0.60692448291575, 0.580213728127373, 0.548228244213276, 
    0.514733354152636, 0.475966236472651, 0.440018078578917, 
    0.398539553924074, 0.354616736308775, 0.309887299584172, 
    0.262262377066798, 0.217009448993895, 0.172790673385415, 
    0.130855620473845, 0.0901273237975842, 0.0559916048890359, 
    0.0292558566809694, 0.0112392570375796, 0.00125769243981883, 
    0.00117237317614749, 0.0109884731158543, 0.029932303399003, 
    0.0569340525474968, 0.0907540268289777, 0.131513310823865, 
    0.172438418356259, 0.21956115302556, 0.26480041565827, 0.309873098288966, 
    0.354951835314063, 0.398137098370095, 0.440292691877007, 
    0.47849903209261, 0.514234250546574, 0.548510436277265, 
    0.578316258895228, 0.608160956224783, 0.635609952298406, 
    0.660729736340193, 0.681972555701499, 0.70550205373526, 
    0.723938115836903, 0.742030686519695, 0.75747145991452, 
    0.772705212502835, 0.78729562565501, 0.800761288396688, 
    0.812491690324143, 0.823662358927837, 0.833713912734426, 
    0.843530604399056, 0.8527850932941, 0.860727562087291, 0.868521426051161, 
    0.875651134740757, 0.881858765118041, 0.888430950890622, 
    0.894476855145831, 0.899900904214311, 0.905417367601548, 
    0.909870215015334, 0.914582685470346, 0.918902506363256, 
    0.922958810751507, 0.926821663623285, 0.930636062411205, 
    0.933812019768272, 0.937234361628245, 0.940211485665713, 
    0.943033052801319, 0.945818413197364, 0.948271177401255, 
    0.951039101588972, 0.953185159625391, 0.955555353206696, 
    0.957706879210764, 0.95967768611086, 0.961666882651854, 
    0.963568984353913, 0.965212595063531, 0.967012180769044, 
    0.968626530573716, 0.969997323113212, 0.97161730770022, 
    0.972967627545747, 0.974422227097121, 0.975659771257357, 
    0.977007133937071, 0.978128598214251, 0.979293695618268, 
    0.980441364885181, 0.981519453964862, 0.982513317404138, 
    0.983534364277392, 0.984458229209041, 0.985407116287369, 
    0.986331642951449, 0.987185770678657, 0.988020914166502, 
    0.988800840229199, 0.989635145765722, 0.990290767345711, 
    0.991054066142094, 0.991711927793217, 0.992407870235365, 
    0.993017824453883, 0.993675858231565, 0.994263918573671, 
    0.994866292790462, 0.995424999236948, 0.995987231905805, 
    0.996509777961354, 0.997023745526167, 0.997532542824115, 
    0.998014459121368, 0.998481727268139, 0.998929237424962, 
    0.99936227239731, 0.999783823633901,
  0.999800213267002, 0.999410191496412, 0.999005029633776, 0.998586276589386, 
    0.998163650070628, 0.997708768020743, 0.997251825982251, 
    0.996780068651906, 0.996276162494164, 0.99578523165081, 
    0.995248780261852, 0.99471480420693, 0.994169906686228, 
    0.993585047059325, 0.992973133651912, 0.992348230367695, 
    0.991717020362079, 0.991059896130367, 0.990306039731665, 
    0.989653898155826, 0.988903170767518, 0.988121118382884, 
    0.987354507624041, 0.986488713308645, 0.985659576552717, 
    0.984817444180849, 0.983886830445823, 0.982902193868926, 
    0.981865211951498, 0.980872384769113, 0.979825065558588, 
    0.978702279275308, 0.977572034593698, 0.976344082053229, 
    0.975002710602399, 0.973736977593503, 0.972334454964699, 
    0.970835588775078, 0.969263061127826, 0.967770081134718, 
    0.966121616108181, 0.964496375226884, 0.96263898803853, 
    0.960734770710306, 0.958718732824837, 0.956632277347923, 
    0.954483960081499, 0.952184489617909, 0.949844730171345, 
    0.94715750323799, 0.944545593567794, 0.941494443629972, 
    0.938627912039862, 0.935620014999714, 0.931917472568837, 
    0.928267191802892, 0.924837278723421, 0.920451002624266, 
    0.916179876704106, 0.911605033815676, 0.906838363656617, 
    0.901465667876519, 0.895981730705593, 0.890281829932352, 
    0.883862973513407, 0.877006914141919, 0.869538522239885, 
    0.862041996576856, 0.853460017977484, 0.844754383932286, 
    0.83438197671823, 0.823592793254753, 0.812948887616031, 
    0.799580598681949, 0.78667630356836, 0.772195097374983, 
    0.756717329566358, 0.739084101193461, 0.719073625244126, 
    0.699034853265929, 0.677121300461102, 0.653701737375243, 
    0.626090325915516, 0.59750350808334, 0.565764607260232, 
    0.532973055714968, 0.496917228080609, 0.459912288308609, 
    0.417431272470817, 0.372187246006695, 0.325561575963778, 
    0.279875124914425, 0.230141420029572, 0.183700782318772, 
    0.140346479115986, 0.0968501793631125, 0.0614924725018473, 
    0.0316746874390985, 0.0119877314318341, 0.0012540967457764, 
    0.00130949185367423, 0.0116872352229263, 0.0320584093678236, 
    0.060994207213525, 0.0971920654640601, 0.138222322454755, 
    0.184563040902091, 0.232146633577522, 0.279106730482671, 
    0.327575211889747, 0.374137364767858, 0.41650784728829, 
    0.459229072752675, 0.497074711800552, 0.533611432945055, 
    0.567815689296909, 0.597351380544917, 0.627317787280513, 
    0.654054466305183, 0.677548320275379, 0.698972256142459, 
    0.720321685677123, 0.739138722523859, 0.756240086597596, 
    0.772650427515771, 0.786518198071861, 0.799718560142126, 
    0.812034523044492, 0.824071871882072, 0.834513970483862, 
    0.843409501849916, 0.853373986214292, 0.862024160415469, 
    0.869914969333785, 0.877088529411132, 0.883932609102385, 
    0.890131782959629, 0.896329822608343, 0.901370122511245, 
    0.906809098212654, 0.911786332785732, 0.916099086849186, 
    0.920507294894582, 0.924755981321553, 0.92843577401767, 0.93199115097465, 
    0.93539636788088, 0.938417955452574, 0.941697479272314, 
    0.944516347491453, 0.94717026955694, 0.949631264617452, 
    0.952193555978674, 0.954494418832307, 0.956565168399234, 
    0.958819294531934, 0.960733435400927, 0.962575362273132, 
    0.96448207812968, 0.966237951903493, 0.967805844246185, 
    0.969399819104683, 0.970836764493848, 0.972344077373124, 
    0.973719293426033, 0.975075161723149, 0.976292420873899, 
    0.977432067202108, 0.978678746953595, 0.979880932936653, 
    0.98090125034645, 0.981930615004237, 0.982880607824501, 
    0.983921577972653, 0.984788263003048, 0.985645443328548, 
    0.986488731404246, 0.987383201318177, 0.988156307681377, 
    0.988930840696019, 0.989649951975611, 0.990417618204016, 
    0.991071610464771, 0.99169512489146, 0.992324531377569, 
    0.992984875312787, 0.993578094327314, 0.994163500087246, 
    0.994702369941558, 0.995255840340198, 0.995773649160547, 
    0.99628132810171, 0.996780485999929, 0.997261913734634, 
    0.997713217417321, 0.998159838018006, 0.998588481299699, 
    0.999007670101421, 0.999410377788252, 0.999798559169073,
  0.999813597137324, 0.999450516507485, 0.999075730396681, 0.998694767569164, 
    0.998286971443393, 0.997881036346444, 0.997444362664677, 
    0.997006753276966, 0.996548879944282, 0.996073952677641, 
    0.99559595771928, 0.99509788017769, 0.994574909104819, 0.994013144296605, 
    0.993464934994348, 0.99288934360086, 0.992298883535707, 0.99165552739523, 
    0.991027314201579, 0.990377074450822, 0.989685558496454, 
    0.988981308410402, 0.988232904206664, 0.987495340043397, 
    0.986689391930984, 0.985815187938729, 0.984982836791428, 
    0.984134620960189, 0.983206786078288, 0.982227327667932, 
    0.981150190483168, 0.980175514046995, 0.979027066747693, 
    0.97791420334884, 0.976850791931011, 0.975539975222955, 
    0.974297608654393, 0.972979396002572, 0.971522608881529, 
    0.969961525657562, 0.968437460028582, 0.966759147833484, 
    0.965211978918654, 0.963425583404181, 0.961538556538281, 0.9596118712972, 
    0.957500848374974, 0.955519234086875, 0.953011616809557, 
    0.950607267320195, 0.94819279090376, 0.945458183571616, 
    0.942560135884979, 0.939565870136157, 0.936476366887364, 
    0.933102553944834, 0.929651225454658, 0.925913478431166, 
    0.921682523575639, 0.917331093253941, 0.912773108313677, 
    0.907756611443307, 0.902836597149354, 0.896824458630257, 
    0.890936100932351, 0.884926251206453, 0.877831430191088, 
    0.87048502621058, 0.862524045259934, 0.853888164176577, 0.84402884455457, 
    0.834582416257334, 0.823411102717044, 0.811749837267336, 
    0.798099839637859, 0.783908160457815, 0.770501002292118, 
    0.752572019663231, 0.734501931898178, 0.713825907680918, 
    0.692875651160901, 0.668765546850795, 0.643537490633295, 
    0.614779606538422, 0.583908129610694, 0.55138821335381, 
    0.515397821546786, 0.477054091764604, 0.435955215882263, 
    0.389045387651815, 0.342173675096715, 0.293957063128478, 
    0.246708740244291, 0.195939743719265, 0.147568064697612, 
    0.105333377888551, 0.0669248963979039, 0.0345147563337198, 
    0.0136259115701329, 0.00160966169869747, 0.0015523940130181, 
    0.0121297772209065, 0.0342706882558623, 0.0659596418380213, 
    0.104479104265243, 0.147875765736785, 0.196276679369965, 
    0.244377138505915, 0.294301386680081, 0.345128195488196, 
    0.38910144944281, 0.43420976911249, 0.476215113340742, 0.514205370410016, 
    0.552057755515452, 0.585006674810443, 0.615097836556127, 
    0.644604667514059, 0.669000911030623, 0.693440201514927, 
    0.714342962669118, 0.733473476910601, 0.751834566063143, 
    0.769122406946591, 0.784323980236166, 0.799196136362551, 
    0.811079702721208, 0.823559799350667, 0.834126123265194, 
    0.844617009387557, 0.853420670400306, 0.862325495366719, 
    0.870426018674182, 0.877704103605469, 0.885307572194772, 
    0.891258380074526, 0.897188565971315, 0.902874708030653, 
    0.907850668202715, 0.9127744979974, 0.917352898790239, 0.92196258772597, 
    0.925807873190379, 0.92943660537721, 0.932999476463184, 
    0.936272946796082, 0.939429598612286, 0.942549898344693, 
    0.945406933907377, 0.948114142400764, 0.950750768321671, 
    0.953225132726522, 0.955218884191944, 0.957531556750443, 
    0.959626318333238, 0.961500266970287, 0.963341506242655, 
    0.965114186137685, 0.966880017868515, 0.968453229010013, 
    0.970042687506981, 0.971569992061323, 0.972914192147685, 
    0.974245156624555, 0.975516526165501, 0.976798484433398, 
    0.977982231554549, 0.979183052484157, 0.98013260248008, 
    0.981161256246776, 0.98221106328603, 0.983180754009001, 
    0.984130441057561, 0.984976986596863, 0.985840972373534, 
    0.986684746132183, 0.987480146627836, 0.98825074823205, 
    0.988960529804102, 0.989696413269992, 0.990348264674656, 
    0.991043882942095, 0.991638310004021, 0.992300060378698, 
    0.992894515161808, 0.99344874421457, 0.994049698823112, 
    0.994563527695559, 0.995093570042028, 0.995589743317854, 
    0.996068632917673, 0.996538834112769, 0.997014473882979, 
    0.997454476372092, 0.997877364113356, 0.998287996974264, 
    0.998689078664417, 0.999074584065117, 0.999451305339559, 0.99981289032071,
  0.999830486069399, 0.999502054933313, 0.999163361144473, 0.998812172443848, 
    0.998451180595549, 0.998081651274563, 0.997689045839372, 
    0.997287928641368, 0.996877617979101, 0.996446977456054, 
    0.996021287316817, 0.995560326901323, 0.995084774100557, 
    0.994605269399345, 0.994104448580012, 0.993580175391184, 
    0.993022469133496, 0.992474819879988, 0.991906033665287, 
    0.991313389252635, 0.990686763215418, 0.990033709920489, 
    0.989372436260251, 0.988677598711847, 0.987961826849481, 
    0.987153175632172, 0.986405475111691, 0.985598101891804, 
    0.984829316649925, 0.983898973142642, 0.982994496877239, 
    0.982077501324844, 0.981054105114093, 0.980026593323306, 
    0.97890102225401, 0.977921796135221, 0.976581526427547, 
    0.975394329367104, 0.974194079699568, 0.972839896949741, 
    0.97137361798772, 0.969978012025225, 0.968475723281091, 
    0.966758520797716, 0.965052709772945, 0.963355622271415, 
    0.961425163706977, 0.959568597582157, 0.957347670540338, 
    0.955200831525697, 0.953035593827387, 0.950551449663637, 
    0.947811083504021, 0.945046556002715, 0.942256823043243, 
    0.938979583868353, 0.935583149523288, 0.932520981642976, 
    0.928767081523293, 0.924631250258357, 0.920734627264157, 
    0.915869221345589, 0.911211317108503, 0.905880694877705, 
    0.900867163906559, 0.894367672376405, 0.887836996178685, 
    0.881409591281708, 0.873836836453833, 0.865576219117493, 
    0.857138839274409, 0.847742947936289, 0.837414539391947, 
    0.826790244252838, 0.813568447238988, 0.800767536991321, 
    0.78589361028741, 0.770519187036025, 0.753248943435176, 
    0.734377528076593, 0.713635161845612, 0.690969233922328, 
    0.665146140540028, 0.640239037216329, 0.609551478504366, 
    0.575330313836517, 0.539713320755002, 0.500684542146499, 
    0.458795299983947, 0.41471501278445, 0.366189475539671, 
    0.315742300240559, 0.263739435468679, 0.211840984226033, 
    0.160790646945028, 0.113926725165864, 0.0709409481393507, 
    0.0376380305860472, 0.0141296077386317, 0.00146854799999999, 
    0.00166464986092317, 0.0142813182682996, 0.0380339952036456, 
    0.0721372517999656, 0.113681751295793, 0.161845562274279, 
    0.211587054532439, 0.263736335249154, 0.315610945957775, 
    0.366433947162058, 0.412920768289453, 0.45894266628891, 0.50059336433775, 
    0.540251724390553, 0.575109129820732, 0.608959235891507, 
    0.638827380122858, 0.666103654468164, 0.692635885857086, 
    0.713615939813804, 0.735281393601945, 0.752577622098637, 
    0.770065109866516, 0.786464116781383, 0.800651247261116, 
    0.813637376100435, 0.826330316771001, 0.837174190945088, 
    0.847757489157062, 0.857063483115133, 0.865905333534456, 
    0.87390306642997, 0.881129744813623, 0.887896925158847, 0.89456939271922, 
    0.900771787719944, 0.905850167563144, 0.910848482281525, 
    0.915991582099372, 0.920700792542809, 0.924615723290018, 
    0.928467350072453, 0.932154001463421, 0.935860152080075, 
    0.939072710068674, 0.942273773323872, 0.944994007219102, 
    0.947965497839995, 0.950341633194103, 0.952980384652007, 
    0.954986541671118, 0.957358020991228, 0.959453336594313, 
    0.961450043483684, 0.963344434470815, 0.965118951040782, 
    0.966752011868033, 0.968292048399592, 0.969906194673455, 
    0.971491336890873, 0.97280868762911, 0.974122435815066, 
    0.975381935495615, 0.976661380990296, 0.977798479397326, 
    0.978927422891518, 0.979927930931588, 0.981073491131044, 
    0.982036718356109, 0.982924920918903, 0.983900812735859, 
    0.984782707099902, 0.985662582554806, 0.986430361640967, 
    0.987193089811044, 0.987898713365709, 0.988650216235888, 
    0.989361465568905, 0.990050351522122, 0.990632300438889, 
    0.991301006326473, 0.991915751606894, 0.992488080582745, 
    0.99302589202357, 0.993567099895393, 0.994094527988759, 0.99459469349315, 
    0.995075487329501, 0.995555706290006, 0.996024979016867, 
    0.996452116692731, 0.996885119137505, 0.997296297960698, 
    0.997697890958082, 0.998072444884019, 0.998449164376005, 
    0.998807259606963, 0.999162254571905, 0.999502903795111, 0.999829754301444,
  0.999835036663103, 0.999518311383696, 0.999189765758987, 0.998852820362082, 
    0.998500739989166, 0.998137044130024, 0.997759569727673, 
    0.997370236158762, 0.996975920860562, 0.996551469958802, 
    0.996130261497096, 0.995678230286804, 0.995261137438959, 
    0.994783227035972, 0.994266887930742, 0.993779650200158, 
    0.993240895283686, 0.992704451679726, 0.992145175420043, 
    0.991540300766204, 0.990939232221303, 0.990325097960637, 
    0.989696593158595, 0.98903425639523, 0.98828041209546, 0.987583266715425, 
    0.986893369315328, 0.986120896233011, 0.985274135274587, 
    0.984349986193072, 0.983473385506211, 0.982570526444331, 
    0.981589629637504, 0.980607069203768, 0.979598622269122, 
    0.978528112003751, 0.977407806503073, 0.97622138227091, 
    0.974987149682672, 0.973611521441493, 0.972302664203314, 
    0.970832616577078, 0.969442731497842, 0.967795279798234, 
    0.966085593180221, 0.96452334028368, 0.96265987376218, 0.960548680354404, 
    0.958504085233815, 0.956489212318163, 0.954399302824939, 
    0.951824166418487, 0.949295178345047, 0.946642551810418, 
    0.943819126765293, 0.940935747970304, 0.937712207674797, 
    0.934402073810531, 0.930870169684098, 0.926958445242911, 
    0.92270715453918, 0.918676416545695, 0.913703643094006, 
    0.908667250580382, 0.903016492400318, 0.897488126931091, 
    0.890448094561002, 0.88389105736906, 0.876934684341701, 0.86963345443989, 
    0.860734334298766, 0.852164625017673, 0.841434191166475, 
    0.830855506125643, 0.818511836826866, 0.806243053077744, 
    0.791877384849326, 0.776253569650713, 0.759907927545518, 
    0.740309308689509, 0.719229560374978, 0.696993894795285, 
    0.672754022559444, 0.645593649986281, 0.61621963418309, 
    0.584186855320007, 0.547938170341024, 0.507518814820895, 
    0.467571625740236, 0.419658511244658, 0.374355702931415, 
    0.321717001284091, 0.267254327139382, 0.217109923138337, 
    0.165919532217935, 0.117098099108785, 0.0747840884357537, 
    0.0388198415971236, 0.0137041325924116, 0.00140923492412752, 
    0.00150118990476102, 0.0149913791462447, 0.0398696141051295, 
    0.074280838435771, 0.118158203025197, 0.165654394662254, 
    0.216326273687192, 0.268735067932545, 0.321862967193871, 
    0.373158321503619, 0.419357680177684, 0.466820926794579, 
    0.50757529465038, 0.548089545271633, 0.581276975764711, 
    0.616020204017479, 0.646265524733194, 0.672327296822946, 
    0.697497272426606, 0.719970137131044, 0.739905491020456, 
    0.758400069303026, 0.77604657176284, 0.792341296200573, 
    0.805650797247962, 0.818831006014102, 0.830656550998918, 
    0.841851773515114, 0.85172683132099, 0.861008987204312, 
    0.869369567866685, 0.877447361532587, 0.885078047093789, 
    0.891077545964124, 0.897385468670967, 0.903219550057539, 0.9084327656975, 
    0.913642091614971, 0.918453319177628, 0.922864364370702, 
    0.926908714670658, 0.930622380518873, 0.934147045510464, 
    0.937582773070789, 0.940895915959037, 0.943944829743995, 
    0.946827891041173, 0.949225488025848, 0.951903557134655, 
    0.954269702656261, 0.956500026159604, 0.958724820471176, 
    0.960618123195883, 0.962616772436674, 0.964516424525472, 
    0.966135365602317, 0.967642673599546, 0.969277025486825, 
    0.970854473005586, 0.972270493139287, 0.973650601168536, 
    0.97489858784705, 0.976191216148862, 0.977365913877058, 
    0.978461625894053, 0.979595482488556, 0.980619338979496, 
    0.981624556844702, 0.982555947464858, 0.983507884419877, 
    0.984372321190364, 0.985201133671095, 0.986029806896063, 
    0.986851698102751, 0.987615827858009, 0.988265037410739, 
    0.989042396582881, 0.989673937206315, 0.990315152597463, 
    0.990957701667883, 0.991556590255461, 0.992137697474322, 
    0.992713782712748, 0.993251575591052, 0.993758953350833, 
    0.994289595881197, 0.994772255208059, 0.995234958577928, 
    0.995697394624484, 0.996131819347647, 0.996561068839683, 
    0.99695724718223, 0.997377720612736, 0.997769761255391, 
    0.998129141242661, 0.998499576131379, 0.998851981594645, 
    0.99918803961795, 0.999516463537512, 0.999835470933612,
  0.9998520931025, 0.999569510387439, 0.999276951496407, 0.998969617357508, 
    0.998662091729373, 0.998341417762832, 0.99800590220891, 
    0.997656167224814, 0.997305000526631, 0.99693443427135, 
    0.996565201866492, 0.996168770406809, 0.995760948131241, 
    0.995337782667772, 0.994909317396084, 0.994453662481025, 
    0.994007294379804, 0.993504335391642, 0.992996340936943, 
    0.992528415237164, 0.991930252003566, 0.991402436328722, 
    0.990797451353302, 0.99020005110533, 0.989620112264965, 
    0.988938296723777, 0.988251480512767, 0.987558496049474, 0.9868200164479, 
    0.986074200896746, 0.985288846842008, 0.984460032027094, 
    0.983655523412718, 0.982738412497069, 0.981812275319701, 
    0.98078766270301, 0.979776741219994, 0.978837890336343, 0.97769249714423, 
    0.976523195923638, 0.97538972871691, 0.973882241870923, 
    0.972656066378997, 0.971263537987528, 0.969699657540845, 
    0.968190129449991, 0.966521343954317, 0.964916372567777, 
    0.962993388337719, 0.961111347657621, 0.959203802621544, 
    0.956918750917437, 0.954494021932133, 0.952333728728761, 
    0.94962585000723, 0.947013331877532, 0.944209709402647, 
    0.941048115947228, 0.937880916919636, 0.934447155063585, 
    0.930876433170365, 0.926556288247668, 0.922167941299343, 
    0.917793341562062, 0.913173850729072, 0.907761194504796, 
    0.901904121403403, 0.895721225865289, 0.888753109959439, 
    0.881630530898061, 0.873745251215707, 0.865483122009929, 
    0.856245265668908, 0.845974358833023, 0.835270079550261, 
    0.822580814601272, 0.810057031975062, 0.79561672772733, 
    0.780259467792381, 0.762248082837412, 0.743403233158999, 
    0.721670770011737, 0.698513575837488, 0.672038823839041, 
    0.640873908577111, 0.610048827613166, 0.575731629407096, 
    0.537212350997116, 0.495027652902951, 0.448678912914741, 
    0.400118894909324, 0.347599941964291, 0.292836022708252, 
    0.236604289536866, 0.180818623630054, 0.128949390106606, 
    0.0824621192408451, 0.0440329773069499, 0.016562496319523, 
    0.00205992301400881, 0.0018219331762163, 0.0165743621022615, 
    0.0441035522293675, 0.0820223190608, 0.129468148171452, 
    0.181465951434082, 0.237039129476795, 0.293618599077556, 
    0.34699908838966, 0.400885571602976, 0.448453485346075, 0.49514321666422, 
    0.536504414697305, 0.575191810440681, 0.610636669066585, 
    0.642583887043179, 0.671935677625223, 0.697034525788565, 
    0.721257405357895, 0.743029867498613, 0.761701831026488, 
    0.779921446976349, 0.7957641431725, 0.810133665615021, 0.822929261862322, 
    0.835279125621711, 0.846299631161166, 0.856260378625515, 
    0.865979386234499, 0.873869369094476, 0.882268396328679, 
    0.889342919216074, 0.895306595813293, 0.902100096348342, 
    0.907426505809417, 0.91299036543921, 0.918137189041727, 
    0.922411467326715, 0.92662122873571, 0.930803500601078, 
    0.934370583140992, 0.937681879796472, 0.941175446755905, 
    0.944204597328979, 0.946963436810385, 0.949798353107748, 
    0.952255482409336, 0.95483345772996, 0.956875128439556, 
    0.959090409613605, 0.961143667019743, 0.963097983290399, 
    0.964769296515238, 0.966606332598491, 0.968094077083978, 
    0.96977242928172, 0.971341444971039, 0.972688330337288, 
    0.973878396863896, 0.975304755741018, 0.976409933275943, 
    0.977678040834003, 0.978768871293219, 0.97985860983364, 
    0.980836984015572, 0.981770813615109, 0.982725641810249, 
    0.983629351289944, 0.984494114961579, 0.985292653886901, 
    0.986077591273253, 0.986881275690136, 0.987589921158576, 
    0.988281038345215, 0.988924924937577, 0.989565517603204, 
    0.990195551069998, 0.99083210366097, 0.991387974092411, 0.99194073589206, 
    0.992517343877811, 0.992980706902214, 0.993503141777481, 
    0.993980298515909, 0.994450721246596, 0.994896083341854, 
    0.995329864003137, 0.995766725137485, 0.996159856017358, 
    0.99654972306181, 0.996937710356496, 0.997300491943043, 
    0.997667159184483, 0.998001934641621, 0.998337949891792, 
    0.998660167570412, 0.998970153225269, 0.999277212881406, 
    0.999569421783912, 0.999852377958233,
  0.999859663485878, 0.999592275331203, 0.999312758953375, 0.999030229313516, 
    0.99872944131411, 0.998423747759474, 0.998106358021765, 
    0.997791420099709, 0.997444710110391, 0.997102078889492, 
    0.996728665096296, 0.99635871736829, 0.995973324810036, 
    0.995594066377623, 0.995180051991241, 0.994768277618792, 
    0.994282934831539, 0.993844278904016, 0.993376346337748, 
    0.992872997943911, 0.992375808914008, 0.991857914428361, 
    0.991302625406415, 0.990742055759782, 0.990135758851448, 
    0.989515808650924, 0.988920031932979, 0.988176921990367, 
    0.987551760195759, 0.986772684277498, 0.986083541361624, 
    0.985271191584174, 0.98442553292219, 0.983581051317405, 
    0.982658479947329, 0.98185181069324, 0.980850640627083, 
    0.979815281628463, 0.978794733353374, 0.977608843928988, 
    0.976618795947336, 0.975331246729177, 0.974045823902601, 
    0.972792986971968, 0.971284098011806, 0.969874354738928, 
    0.96815459808266, 0.96668694475646, 0.96486585197795, 0.963078509272094, 
    0.961187812696377, 0.959152641940278, 0.957003329640259, 
    0.954546141564825, 0.952135499891918, 0.949650978792047, 
    0.946986229795426, 0.943990510143283, 0.940802698637821, 
    0.937664966169811, 0.933972707129773, 0.930143657857493, 
    0.926374062788191, 0.921763147354024, 0.917199087924756, 
    0.911570150794461, 0.906480797254664, 0.901061455194642, 
    0.894160540894099, 0.887004137965664, 0.879880481763335, 
    0.871778244638652, 0.862696149781291, 0.852968511227217, 
    0.842714593463347, 0.830703512955263, 0.818143210825219, 
    0.804038248976748, 0.788829833838813, 0.770766789561403, 
    0.753351598978372, 0.731160408151591, 0.70891422255406, 
    0.682956620687695, 0.655212820465747, 0.62341249268537, 
    0.588463597503928, 0.549617859432447, 0.508320829442744, 
    0.462282044993349, 0.412960585456608, 0.359253451452297, 
    0.303466264033157, 0.245720602156686, 0.189697461789869, 
    0.135778251472096, 0.0857337533002099, 0.0465810172624319, 
    0.0169299402543477, 0.00216197253763299, 0.00185543884844859, 
    0.0169040464649596, 0.0467897143348083, 0.0868022273251411, 
    0.134898499787563, 0.189383261311617, 0.247367503052809, 
    0.304179877890816, 0.359243366450448, 0.412504042920783, 
    0.462745976673739, 0.507819033131227, 0.550196680647141, 
    0.588669183536034, 0.623737287097517, 0.654126507284099, 
    0.683564785119768, 0.708151548868317, 0.732354784137994, 
    0.752824267716427, 0.772043744982995, 0.787520594058088, 
    0.804484873408677, 0.818025884267297, 0.83008187057132, 
    0.842675026892697, 0.853409638396575, 0.863406733638947, 
    0.872225828667194, 0.87978246750011, 0.887313552344644, 
    0.894280636157277, 0.900285915637865, 0.906199489805738, 
    0.911954236459067, 0.917033748510524, 0.921775735901472, 
    0.926060691466934, 0.930260758872007, 0.933713360352523, 
    0.937441663054812, 0.941045988913695, 0.944013726710286, 
    0.946852232827943, 0.949583091345139, 0.952245776762192, 
    0.954675033694929, 0.956851438127937, 0.959172123392309, 
    0.960983225665885, 0.963080518558972, 0.964913565364222, 
    0.966602312758394, 0.968294552490217, 0.969784588755657, 
    0.971258548470046, 0.972683181067683, 0.974017374979742, 
    0.975268160034065, 0.976574158668746, 0.977728278555642, 
    0.978811848225145, 0.979916616617771, 0.980992128363298, 
    0.981855464996298, 0.982742729325566, 0.983557351653928, 
    0.984460990373021, 0.985360435649966, 0.986059849476636, 
    0.986712949034395, 0.98754224160576, 0.988220086024933, 
    0.988908752201211, 0.989529062079137, 0.990153884070919, 
    0.990732799066092, 0.991315795596587, 0.991813111482317, 
    0.992369969131067, 0.992885591587321, 0.993359134240779, 
    0.993849953409148, 0.994316337735502, 0.994744975425579, 
    0.995181378495052, 0.995578970074558, 0.995972289080633, 
    0.996368225826667, 0.996730610906256, 0.997096760509823, 
    0.997447774061775, 0.997783221635276, 0.998106920910997, 
    0.998421124237049, 0.99873299023828, 0.999025598151056, 
    0.999314240892197, 0.999591313949866, 0.999859349283015,
  0.999865466584164, 0.999610608435177, 0.999348761718882, 0.999077502201815, 
    0.998794041610005, 0.998507552090267, 0.998208474256043, 
    0.997889459791408, 0.997581217761223, 0.997239721890708, 
    0.996899432054134, 0.996543128162079, 0.996188031918452, 
    0.995812763329446, 0.995414758396667, 0.99500590099088, 
    0.994574340407158, 0.994148437358359, 0.993682946257903, 
    0.993226735607194, 0.992740900857718, 0.992220318509106, 
    0.991716323784523, 0.991179458938975, 0.990607315231553, 
    0.990041158990726, 0.989435371123687, 0.988781528265036, 
    0.988138736829734, 0.987456075674404, 0.986786403472318, 
    0.985972905192826, 0.985140718482192, 0.984397763254311, 
    0.983550750724942, 0.982723097856816, 0.981793925553067, 
    0.980824538773984, 0.979779163767148, 0.978787490721159, 
    0.977634135479916, 0.976463515679215, 0.975231721786953, 
    0.974007060654382, 0.972769785032483, 0.971198265837583, 
    0.969778319990039, 0.968297220251306, 0.966673925720437, 
    0.964839029567402, 0.963123279744506, 0.960970492751085, 
    0.958941358638596, 0.956947102927196, 0.954503476985718, 
    0.952187694116526, 0.949470462033602, 0.946615378941634, 
    0.943577866274029, 0.940252803812298, 0.93710434810483, 
    0.933310968979853, 0.929554256086507, 0.925264238528321, 
    0.920552532456222, 0.915964806133216, 0.910517043796801, 
    0.905102120350804, 0.898953689875171, 0.891689454504403, 
    0.885581495543217, 0.877472563354218, 0.868509158235971, 
    0.859002184200431, 0.84911142507671, 0.837663367288598, 
    0.825333903426159, 0.811885387134956, 0.797627629277805, 
    0.780044407041469, 0.76215953045406, 0.74145516845146, 0.718693476288345, 
    0.69452506066413, 0.666384566960966, 0.63504857926946, 0.601790269734396, 
    0.562573745757766, 0.521700929067618, 0.475173155874219, 
    0.424461968840869, 0.372243759486311, 0.31450161285631, 
    0.257208802412054, 0.196353358783756, 0.141846570230379, 
    0.0905834541097855, 0.0477545056643998, 0.017511500272288, 
    0.00191898134767347, 0.00218620064756123, 0.0181862491811316, 
    0.0488970456232753, 0.0901156357987218, 0.141092041508979, 
    0.198474822553235, 0.25680204029076, 0.313676657671295, 
    0.370321509047684, 0.424125787637882, 0.476840241927574, 
    0.521235940239105, 0.561522365638445, 0.60091769622133, 
    0.635515665569464, 0.666359260560125, 0.693498313961401, 
    0.718691584489521, 0.741782100555639, 0.762312196333675, 
    0.780678791994356, 0.797033069834698, 0.812023654519788, 
    0.825619251351907, 0.838005006521974, 0.848895987262422, 
    0.858641573813743, 0.868546730323296, 0.876900903339697, 
    0.884595472024474, 0.892420690260272, 0.899008854458744, 
    0.904927682646471, 0.91088909056094, 0.915896136456453, 
    0.920665404510218, 0.925232190200002, 0.92961276204297, 
    0.933190539240682, 0.936788137186883, 0.940450949197602, 
    0.943669748166769, 0.946528152992856, 0.949460436213064, 
    0.952012553074835, 0.954512993079774, 0.956913748888052, 
    0.958929744675599, 0.961044822403905, 0.962735803373589, 
    0.964746124309564, 0.966549689256992, 0.968292875590957, 
    0.969742285394312, 0.971288969813273, 0.972722190723838, 
    0.974011623799585, 0.97528360470266, 0.976503129017385, 
    0.977710647738297, 0.97870560303572, 0.979763627257127, 
    0.980849754126599, 0.981808525713644, 0.982711337395085, 
    0.983564790299858, 0.984429381220549, 0.985261573249092, 
    0.98601209274105, 0.986791330671197, 0.987476938153663, 
    0.988146652334657, 0.988766813101644, 0.98943171332314, 
    0.990043403048509, 0.990631882563979, 0.991174923705269, 
    0.991743933836113, 0.992242865447558, 0.992738180535582, 
    0.99323676247326, 0.993682551591733, 0.994151912639783, 
    0.994582752083658, 0.995015641168273, 0.995404707993185, 
    0.99580550859886, 0.996185508652036, 0.996545831674827, 0.99690123779651, 
    0.997244025767289, 0.997569822378678, 0.997904345854401, 
    0.998202073366158, 0.998498363454784, 0.998793899461028, 
    0.999074902701363, 0.999349163842377, 0.999611986187694, 0.999866270721148,
  0.999868397964182, 0.999618836425232, 0.999365066985028, 0.999099191658601, 
    0.998817264514754, 0.998539317824042, 0.998243931558823, 
    0.997946414280561, 0.997629865190784, 0.997306688132856, 
    0.996986647161747, 0.996638208560205, 0.996266340508039, 
    0.995889392098917, 0.995516964202913, 0.995123622206912, 
    0.994712513698133, 0.994290589280757, 0.993837857140603, 
    0.993379496758787, 0.992903954952185, 0.992445219266361, 
    0.991897439006835, 0.991406276282139, 0.990827011647402, 
    0.990278030371502, 0.989694074552683, 0.989084244027146, 
    0.988413396871777, 0.987805781972226, 0.987084286769272, 
    0.986340772509582, 0.985577564380454, 0.984819449337, 0.983944587176416, 
    0.983126466048628, 0.982247293409535, 0.981323536780432, 
    0.980308508299901, 0.979188779146716, 0.978289849959911, 
    0.977121649793707, 0.975853531279622, 0.974629455094327, 
    0.973295146289876, 0.971915345514347, 0.970483592124518, 
    0.96905834185641, 0.967351615161926, 0.96552599607393, 0.963924475631821, 
    0.962022416555081, 0.959877107157356, 0.957709461180107, 
    0.955631498085979, 0.953113752365774, 0.950572777160786, 
    0.94779072673178, 0.944821192129739, 0.94166682915595, 0.938392415255634, 
    0.934962227494142, 0.931067345405277, 0.926873217997304, 
    0.922365954180315, 0.91762215428343, 0.912663638694505, 
    0.907138122526506, 0.900844973567669, 0.894534050207657, 
    0.887089184732762, 0.879607703757872, 0.87145382652833, 
    0.862184872063804, 0.851798995190339, 0.841519410752629, 
    0.829048861980112, 0.81499573930252, 0.80044715908972, 0.784669862552961, 
    0.76730786967763, 0.746272655506394, 0.724116672077889, 
    0.699229638378779, 0.671468156463114, 0.641135024275083, 
    0.606287586799575, 0.568887165603728, 0.527487404694218, 
    0.481225373872934, 0.430957604573876, 0.376642830395709, 
    0.319819621501388, 0.261689207652077, 0.202002810282443, 
    0.144227667097205, 0.0926849199897928, 0.04988989831933, 
    0.018208237230666, 0.00216851484073608, 0.00193353222628366, 
    0.0187819155880043, 0.049613744767073, 0.0923919514357116, 
    0.145540141536351, 0.201719031799745, 0.260390839890375, 
    0.321703651708662, 0.37637607351535, 0.430255704169736, 0.4795128279617, 
    0.529109665819663, 0.569466491265889, 0.607169866472677, 
    0.642109658049499, 0.671861675132795, 0.698016455607407, 
    0.724146707288418, 0.747132546283189, 0.766347998638965, 
    0.784125687644174, 0.800435731144526, 0.815673113481404, 
    0.828961105178988, 0.840465969357672, 0.852058398371744, 
    0.862304233427663, 0.871180342180353, 0.879847540187414, 
    0.887288654053547, 0.894457641798328, 0.901012564273509, 
    0.90679826626251, 0.912506470178694, 0.917888449767781, 
    0.922624037468982, 0.926808030019666, 0.930924433139015, 
    0.934909308549447, 0.938522868363964, 0.941695397920712, 
    0.944852128534615, 0.947763140800038, 0.950588580590428, 
    0.953071407843109, 0.955576922580414, 0.957980459377666, 
    0.959912009994222, 0.961863153943657, 0.963707769163113, 
    0.965610981581854, 0.967217978883658, 0.969016743850495, 
    0.970478556234808, 0.971932787406907, 0.97336377111492, 
    0.974602674868037, 0.975969295363203, 0.977079589015308, 
    0.978257719231051, 0.979328758840013, 0.980448245597267, 
    0.981283520636305, 0.982210000898621, 0.983132725507106, 
    0.983934967040084, 0.984811222256973, 0.985580907446106, 
    0.986325313817734, 0.987075920625539, 0.98776936842952, 
    0.988441591635769, 0.989054673027677, 0.989652538161312, 
    0.990286640133887, 0.990859241959783, 0.99139974746371, 
    0.991903977664604, 0.992459798126047, 0.99292193059796, 
    0.993375579013508, 0.993848754282303, 0.994281157274939, 
    0.994715092462535, 0.995124481114245, 0.99552664817325, 0.99589608098777, 
    0.996280106116539, 0.996625784399303, 0.996979106660761, 
    0.997304387455731, 0.997634189971309, 0.997943764264454, 
    0.998246907226113, 0.998537552719705, 0.998824462514318, 
    0.999097157888666, 0.999362360221718, 0.999620654171869, 0.999869348939569,
  0.999876866130344, 0.999645651655607, 0.999405093809877, 0.999156035850542, 
    0.998906048147321, 0.99864005818026, 0.998363612650162, 
    0.998078544817317, 0.997791907839711, 0.997486028604174, 
    0.997180185995703, 0.996845891709463, 0.996529334353881, 
    0.996178888369285, 0.995816140812528, 0.995439422771976, 
    0.995080921094138, 0.994694594991476, 0.994253043399556, 
    0.99384513512447, 0.993395235866998, 0.992938699366765, 
    0.992442559084464, 0.991991342903538, 0.991447786224934, 
    0.990907312984714, 0.990380512051042, 0.989838747061618, 
    0.989191858803442, 0.988543735479461, 0.987926022869174, 
    0.987276196055982, 0.98654497500534, 0.985844190366545, 
    0.985077483166284, 0.984271955933873, 0.983465404947984, 
    0.982514286527084, 0.981597873418158, 0.980667430641312, 
    0.979646445333061, 0.978546643159653, 0.977454124401742, 
    0.976412894660783, 0.975133748017475, 0.973745758367338, 
    0.97243362513397, 0.971104022685543, 0.969511734213733, 
    0.968031321742156, 0.966165600095958, 0.964463813318704, 
    0.962581592065634, 0.96046652264885, 0.958344389717509, 
    0.955988903392194, 0.95376664766209, 0.951130584762808, 
    0.948544967737231, 0.945606304497468, 0.942276516603073, 
    0.938840632829098, 0.935313262005882, 0.931541085314205, 
    0.927372919523515, 0.922631791660188, 0.918254655744632, 
    0.912960407177402, 0.907059789339378, 0.900957723233261, 
    0.894174892004603, 0.887034081893676, 0.878800470029417, 
    0.870307910796173, 0.860874973269337, 0.850252392189251, 
    0.838463113122134, 0.826162519618323, 0.810951887421341, 
    0.795636323839989, 0.778204524411643, 0.759214544652157, 
    0.737767369405834, 0.712802111707992, 0.686628024563545, 
    0.657068252277344, 0.622672616373809, 0.585334196526642, 
    0.543922561965485, 0.498890019201202, 0.44777824181481, 
    0.394815789662698, 0.335156320719055, 0.276481112782926, 
    0.211710117043384, 0.151426852831484, 0.0984312339121549, 
    0.0526910914136973, 0.0198928914105318, 0.00238770207299147, 
    0.00212510282972675, 0.02006789008782, 0.0515331711738187, 
    0.0994843332792578, 0.153116310318343, 0.212422633489428, 
    0.275155903531948, 0.333597411923303, 0.393506884180255, 
    0.446040457750544, 0.497499722921073, 0.544330328841649, 
    0.586188789919396, 0.623435772247954, 0.656900354311719, 
    0.686486912177561, 0.712482666747613, 0.736889199756196, 
    0.759048760013591, 0.778802281719091, 0.796174289725908, 
    0.812015863380945, 0.825389948246303, 0.838520603729644, 
    0.849850206660958, 0.860646692815728, 0.87042487089478, 
    0.879010061978724, 0.886522227036998, 0.894294074238268, 0.9015588254225, 
    0.907517310485886, 0.912745548424131, 0.917930192071353, 
    0.922989548838838, 0.927531377820913, 0.931587997668593, 
    0.935547750258777, 0.939193835905289, 0.942334420805014, 
    0.945378424484049, 0.948451310324827, 0.951099598143288, 
    0.953708018068226, 0.956274290458388, 0.958496159289516, 
    0.96054984059916, 0.962501639931461, 0.964393026141441, 0.96624678647295, 
    0.967818179061515, 0.969459306741463, 0.971074627690992, 
    0.972470200842973, 0.973770457339763, 0.974983540296922, 
    0.976353979745216, 0.977436145475177, 0.978598496889263, 
    0.979683249306112, 0.980616022298204, 0.981670387844031, 
    0.982519035749217, 0.983402246426611, 0.984208712067351, 
    0.985029530608794, 0.985839746448713, 0.986596217035199, 
    0.987260644004236, 0.987984342614076, 0.98860884104348, 
    0.989192632874116, 0.989781455511375, 0.990404166450232, 
    0.990932895330341, 0.991443050100574, 0.991965582450236, 
    0.992447550532356, 0.992940801687948, 0.993397504750036, 
    0.993816826976419, 0.994268536704808, 0.99467185891433, 
    0.995095701910567, 0.995452467663802, 0.995829779929182, 
    0.996195605623645, 0.996523373259944, 0.996858356516828, 
    0.997173352751363, 0.997491399903959, 0.997793199903244, 
    0.998086141680898, 0.998368402768184, 0.998639354036298, 
    0.998905600922037, 0.999157656476705, 0.999405908223829, 
    0.999646535686924, 0.999877469134928,
  0.999882142726552, 0.999660150724533, 0.999428312088553, 0.999195025038078, 
    0.99895030717009, 0.998693481650468, 0.998433992301237, 
    0.998162861605551, 0.997891068196116, 0.997603347376965, 
    0.997309274985101, 0.996993080291533, 0.996664041846827, 
    0.996343723393677, 0.996005684287534, 0.995651418769686, 
    0.995275083232318, 0.994893438521473, 0.994504632402874, 
    0.994107754173903, 0.99366346093456, 0.993239371541902, 
    0.992818908288568, 0.992307410199454, 0.991826863016836, 
    0.991305886661205, 0.990780975968063, 0.990228793851825, 
    0.989707172735263, 0.989072941716538, 0.98842064530549, 
    0.987792673792796, 0.987151968364461, 0.986403987986911, 
    0.985664117285528, 0.984931413651031, 0.98410056886908, 
    0.983320199805524, 0.982440586997601, 0.981537770472108, 
    0.980497848440831, 0.979479394725619, 0.97841897524047, 
    0.977383205590934, 0.976014712396065, 0.974858596360861, 
    0.973564259132809, 0.972323682625733, 0.970725783899761, 
    0.969253581537539, 0.967661574369348, 0.965978696106809, 
    0.964105579928309, 0.962177882555039, 0.9600685373456, 0.958170864806677, 
    0.955711059695852, 0.953319253966736, 0.950405197795075, 
    0.947780425889512, 0.94472476908189, 0.941528527225338, 
    0.938251537133676, 0.93400689180383, 0.930413321449559, 0.92582044649617, 
    0.921231350254087, 0.916431104352603, 0.910878491071117, 
    0.904733745745911, 0.89833103558643, 0.891452247722923, 
    0.883454729268944, 0.875208718817255, 0.866170250491016, 
    0.856125695968951, 0.844773046028365, 0.832339561899223, 
    0.817729853682851, 0.803173351951242, 0.786114918304713, 
    0.767346188282613, 0.746625272184213, 0.723219437974193, 
    0.696056752961404, 0.666554983559318, 0.632621128134993, 
    0.595655108350425, 0.553801758453382, 0.510446061736278, 
    0.458767790311307, 0.40395089104591, 0.345255025864315, 
    0.283488607837214, 0.222248339140854, 0.158317034474519, 
    0.104325721066803, 0.0556747687186438, 0.0209108957261566, 
    0.00226307913921807, 0.00227298237511963, 0.0201451496518548, 
    0.0560100118390799, 0.103586380055026, 0.159521371297216, 
    0.217594894184287, 0.282468333315627, 0.343081094963945, 
    0.403991550799651, 0.45752545298309, 0.510282184167907, 
    0.555024838728696, 0.597219464935784, 0.633498971688338, 
    0.665775937711618, 0.696170039365329, 0.721156148616413, 
    0.746138719647159, 0.768446135265649, 0.785654979515492, 
    0.802685748560691, 0.818228208872717, 0.832418263146699, 
    0.84433098296431, 0.855684716113908, 0.865635312144339, 
    0.875280757776578, 0.883937633602324, 0.891421490445521, 
    0.898391771495057, 0.904738653290561, 0.910663175400423, 
    0.916419343397012, 0.921117129643443, 0.925904149327172, 
    0.930483861084633, 0.934386538234916, 0.938002066954983, 
    0.941596451914404, 0.944735868421485, 0.947858374157571, 
    0.950534290644908, 0.953105731317847, 0.955641413998221, 
    0.958011809233585, 0.960109561205084, 0.962141696601634, 
    0.964073265600776, 0.965834032767242, 0.967689653443087, 
    0.969083828378237, 0.970690331977045, 0.972281321470175, 
    0.97363894181552, 0.974901820438692, 0.976185142853486, 
    0.977376735926672, 0.978458712106473, 0.979480104639355, 
    0.98057564753598, 0.981485525472568, 0.982428554034115, 
    0.983267397331773, 0.984076135064308, 0.984946759538915, 
    0.985679026712556, 0.986420723937084, 0.987111166826609, 
    0.987735825628065, 0.988524305795225, 0.989073661562182, 
    0.989673801119909, 0.990221482756731, 0.990801509567594, 
    0.991347567511494, 0.991827125865932, 0.992322640812507, 
    0.992791902997017, 0.993259166643725, 0.99367576000033, 
    0.994106134506754, 0.994512375951173, 0.99491283862221, 
    0.995284384375896, 0.995643941553559, 0.996009726060775, 
    0.996325656023342, 0.996669734399733, 0.997000548590794, 
    0.997294498832821, 0.99759525800972, 0.997889650944669, 
    0.998166704484335, 0.998435832550763, 0.998696393951887, 
    0.998948404339882, 0.999194564325167, 0.99942971229421, 
    0.999659729609713, 0.999882260745066,
  0.999901752188654, 0.999718885895073, 0.999529865493523, 0.999335805191204, 
    0.999137544429098, 0.998927662931529, 0.998709116052482, 
    0.998483092920944, 0.998258202364042, 0.998022244613111, 
    0.997774706462896, 0.99752661982193, 0.997265412205485, 
    0.996993041353159, 0.996707006102038, 0.996415339968331, 
    0.996128170761567, 0.995806687644187, 0.995479685423031, 
    0.995139508484755, 0.994798669256951, 0.994443646749342, 
    0.994082275261847, 0.993694888596143, 0.993272756222323, 
    0.992863846320945, 0.992397081735743, 0.991975129494635, 
    0.991482921945936, 0.991031395781325, 0.990511509043984, 
    0.989955898402462, 0.989407447503182, 0.988833496607271, 
    0.988206653596178, 0.98760792252558, 0.986948120732521, 
    0.986313248778938, 0.985467111405895, 0.984740814401316, 
    0.983967033125558, 0.983087345221219, 0.982156121451362, 
    0.981293932415528, 0.980307221604327, 0.979352720283104, 
    0.97822219057345, 0.977018131943222, 0.975946579869176, 
    0.974660952647493, 0.9731959059514, 0.971834677893137, 0.970285703690214, 
    0.968719253555924, 0.966940109083521, 0.965061055953575, 
    0.963276456557822, 0.961305006353235, 0.958923728299532, 
    0.956557034146207, 0.953972494347369, 0.951381846597303, 
    0.948465092041255, 0.945428680912145, 0.942094724780185, 
    0.938155430969639, 0.934069322579274, 0.929979561889388, 
    0.925104929264244, 0.92022620138313, 0.914872882939999, 
    0.908795145820258, 0.9021787245896, 0.895040275742275, 0.886812405993601, 
    0.878639320055109, 0.868226113505929, 0.857432777833447, 
    0.844948233366235, 0.831721768440033, 0.817158839807206, 
    0.800050248986441, 0.781351541992174, 0.7590410030755, 0.736497033896536, 
    0.707896933750107, 0.676004841888311, 0.641059922633978, 
    0.603973896208129, 0.558285004350815, 0.507396694239094, 
    0.451710221365692, 0.389248690708019, 0.323904215191347, 
    0.254955344483887, 0.186757849014746, 0.122451632042482, 
    0.0666061747201185, 0.0252961504947816, 0.00274102946494491, 
    0.0027096735838916, 0.0248380542205255, 0.0663687551567626, 
    0.120679261762286, 0.188120525886886, 0.256076190565536, 
    0.322803368830225, 0.39022192645613, 0.453283187022958, 
    0.506281673472795, 0.557015387605358, 0.603485385963842, 
    0.641528240022288, 0.677848499743819, 0.707516135674196, 
    0.73561956423405, 0.760380237875815, 0.780589974512991, 
    0.800162776962228, 0.816627339516278, 0.831634846987422, 
    0.845055360941258, 0.857401342614342, 0.86827034484423, 0.87775186783526, 
    0.886947204103414, 0.894921621673583, 0.901800663625422, 
    0.908811871318664, 0.914873951261172, 0.920367500610923, 
    0.925450319104259, 0.929979354695679, 0.934322063620258, 
    0.938253831441852, 0.94189792728385, 0.945304142771085, 
    0.948557210652803, 0.95133576548827, 0.954031847911276, 
    0.956518553834437, 0.95885392082811, 0.96110783588334, 0.963348429022389, 
    0.965215283878115, 0.966956153011636, 0.968645582588091, 
    0.97015205359028, 0.971799164450579, 0.973249876297538, 
    0.974573090189775, 0.975854974894335, 0.977053469422843, 
    0.978188634950235, 0.979333832626241, 0.980412129946072, 
    0.98127198657256, 0.982229886204898, 0.983110299694508, 
    0.983929400869235, 0.984778229940843, 0.985499239535079, 
    0.986207927964215, 0.986902634650518, 0.98754859507011, 
    0.988229329227073, 0.988831086830971, 0.989449960991479, 
    0.989938407662971, 0.990486485538826, 0.991016003626146, 
    0.991492501665434, 0.991951528115205, 0.992443668079967, 
    0.992870015872457, 0.993314319329094, 0.993702007053471, 
    0.994062588686914, 0.994439391203369, 0.994824761719346, 
    0.995136340265668, 0.995500407083559, 0.995808619477064, 
    0.996111194657368, 0.996413751406022, 0.996706430606652, 
    0.996984576873445, 0.997264155442507, 0.997531853197844, 
    0.997783573169794, 0.998021630777856, 0.99825758759225, 
    0.998485645789896, 0.998711872410552, 0.998923608542354, 
    0.999134398346899, 0.999333659778582, 0.999530713903384, 
    0.999718575352448, 0.999901311503664,
  0.999915340272951, 0.999759579217283, 0.999599035037202, 0.999433772845281, 
    0.999262644732496, 0.999088096441456, 0.998904944891073, 
    0.998716395854043, 0.99852203103113, 0.9983204160154, 0.998114542039117, 
    0.997896692313789, 0.997676390462448, 0.997447692970683, 
    0.997202519614997, 0.99696168309232, 0.99670875863884, 0.996439823364869, 
    0.996160969770755, 0.995876161087083, 0.995577484846091, 
    0.995282261560968, 0.994958439209701, 0.994634715606865, 
    0.994304842206153, 0.993930482641049, 0.993545730288992, 
    0.993180146433194, 0.992799090151453, 0.992355466081592, 
    0.991897467471271, 0.991484493336814, 0.990999525072897, 
    0.990485586970121, 0.98997850808026, 0.989463555814467, 
    0.988859434281078, 0.988293585208025, 0.987627496156042, 
    0.986969817144559, 0.986325995501906, 0.985625807111959, 
    0.984877495635677, 0.984041721503378, 0.98323237160961, 
    0.982347733881618, 0.981432313719758, 0.980456131326088, 
    0.979388312138409, 0.978358797631285, 0.977154269771398, 
    0.976020709190856, 0.974648417664815, 0.973260793933548, 
    0.971905399577869, 0.970206581481242, 0.968622391096317, 
    0.966825104446233, 0.96477889751267, 0.962752647257018, 
    0.960851300296925, 0.958389794327661, 0.955847402376695, 
    0.953074531872415, 0.950200842705761, 0.947046253213762, 
    0.943438128124295, 0.939830332152598, 0.935939459100664, 
    0.931312294484123, 0.926587928893111, 0.921590764086744, 
    0.915694576630855, 0.908962846755856, 0.902324019933741, 
    0.894669156889957, 0.885749557395698, 0.87620677263399, 
    0.865629231345605, 0.853424878183419, 0.839842635014667, 
    0.824055016497607, 0.807375007522368, 0.787638594760241, 
    0.764953779441653, 0.74014397685712, 0.712428833843773, 
    0.678600005985873, 0.640606553844494, 0.597994384961069, 
    0.549264465240855, 0.490250567362083, 0.430117026709098, 
    0.361190390047433, 0.28670575265912, 0.212652656351315, 
    0.140339473541236, 0.0755842000307551, 0.0290743439522593, 
    0.00363162956908924, 0.0030996975476672, 0.0283284340396093, 
    0.0767678724554838, 0.140973310066624, 0.213000668936952, 
    0.288052444277677, 0.360154898596541, 0.43088051454909, 
    0.491690291317845, 0.548469788573512, 0.596078604344488, 
    0.640523862084266, 0.677697994184721, 0.71260967804216, 0.74106295907846, 
    0.765725186629503, 0.788212436873897, 0.807489505974494, 
    0.825343325589263, 0.839861315620992, 0.853724079404213, 
    0.865216524004695, 0.876350435444256, 0.885529221447114, 
    0.894522517018428, 0.902275839372001, 0.909356968223119, 
    0.915761561578979, 0.921548804880854, 0.926525539611876, 
    0.931476542359265, 0.935837754702424, 0.939767411030701, 
    0.94380230282434, 0.947291452896967, 0.950235284827294, 
    0.953119173057196, 0.955861614236465, 0.958601627403772, 
    0.96071775061271, 0.962864386505195, 0.964912737387403, 0.96679328523365, 
    0.96862365603411, 0.970177893702164, 0.971807146710388, 
    0.973315323638374, 0.974639801961113, 0.975944053063673, 
    0.977157551324463, 0.978401338649396, 0.979403172138288, 
    0.980451934240469, 0.981400362043205, 0.982434262321595, 
    0.983238479690101, 0.984002936385572, 0.98491558307632, 
    0.985594487340791, 0.986351368264198, 0.987035696910785, 
    0.987649057494291, 0.988308339498752, 0.988864596602772, 
    0.989443675487727, 0.989988440059739, 0.990468573858892, 
    0.990971286779401, 0.99145807447573, 0.991923440196787, 
    0.992359649805431, 0.992752067913738, 0.9931851716453, 0.993564601895325, 
    0.993922857836875, 0.994294482448818, 0.994630029568568, 
    0.994960476505526, 0.995268138151556, 0.995607184394319, 
    0.995885896611379, 0.996169561445012, 0.996438213630557, 
    0.996705546604874, 0.996960885243127, 0.997208908472461, 
    0.997445752862476, 0.997675151345988, 0.99790100668566, 
    0.998118135217431, 0.99831962917733, 0.998522445058731, 
    0.998712999825699, 0.998902336610348, 0.99908714714925, 
    0.999261028643692, 0.999433711915183, 0.999600214395976, 
    0.999760517333471, 0.999915253344729,
  0.999924981781433, 0.999790249156954, 0.999651038159634, 0.999507185138351, 
    0.999358349723841, 0.99920803007819, 0.99904628801091, 0.998884072360064, 
    0.998712794315197, 0.998536428024767, 0.998360429790307, 
    0.99816852255783, 0.997978218456356, 0.997779091283135, 
    0.997587062137543, 0.997358376279909, 0.997144656481336, 
    0.996910294432366, 0.996668785467596, 0.996420636174792, 
    0.996169494086247, 0.995897295487445, 0.995627631626964, 
    0.995327518471994, 0.99503877946333, 0.994740582641512, 
    0.994393420767095, 0.994070979756589, 0.993748371471106, 
    0.993357584050992, 0.992955825234348, 0.99258583270463, 0.99214314843598, 
    0.991712025197001, 0.991272747286228, 0.990831553121783, 
    0.990326442772485, 0.989782603063896, 0.98930407595331, 
    0.988700438127163, 0.98804014882106, 0.987485125606062, 
    0.986839452641876, 0.986125174555035, 0.985455066141262, 
    0.984575118044654, 0.983810849565792, 0.982986063975335, 
    0.982046314226874, 0.981126540737271, 0.980071176843487, 
    0.978997532137693, 0.977940303348903, 0.976691236196767, 
    0.975473825863298, 0.974137136835521, 0.972520077910852, 
    0.971098668173438, 0.969252100046964, 0.967525108267731, 
    0.965847843524755, 0.963626792182107, 0.961435654914364, 
    0.958970069673001, 0.956402417960318, 0.953644043969434, 
    0.950679515157133, 0.947624995496557, 0.943941454080427, 
    0.939926465353424, 0.93552332387277, 0.931102361814986, 0.9259076352444, 
    0.920176762964133, 0.913806497715383, 0.906818561735477, 
    0.899323239016405, 0.891030042596504, 0.881180709513565, 0.8694453540701, 
    0.857840585307801, 0.843916274409206, 0.828703253405365, 
    0.810640008178263, 0.79075086946481, 0.765800669272012, 
    0.739488537713985, 0.708110015106318, 0.671841646795617, 
    0.628790430307698, 0.582427490416114, 0.52754443106157, 0.46360954967235, 
    0.392911701619391, 0.317481751974216, 0.236025617961835, 
    0.158178812247233, 0.0874263238522743, 0.0341796812027832, 
    0.00361313421822649, 0.00388267996240891, 0.0338893153977205, 
    0.0868671646441685, 0.1586999210999, 0.236853316416411, 
    0.318032416311497, 0.393475930783313, 0.463873501312453, 
    0.526143652650628, 0.580998580396424, 0.630405367581056, 
    0.672068665022429, 0.707889956713939, 0.73917859591153, 
    0.766531102035146, 0.790356740143733, 0.811026343369154, 
    0.82882842680198, 0.843597271408436, 0.85801319443814, 0.870345429332049, 
    0.880639206712014, 0.890512382340747, 0.899334259387973, 
    0.907018374271551, 0.913847002023516, 0.920125944078177, 
    0.925867076121859, 0.931025613520872, 0.935695879299939, 
    0.940009879210638, 0.943794513693551, 0.947351650072578, 
    0.950649501477653, 0.953596069322228, 0.956412385924854, 
    0.958958872965142, 0.961598035815449, 0.963652217679473, 
    0.965641087569817, 0.967449521918812, 0.969307611489296, 
    0.971026492449756, 0.972619656648421, 0.974080964436009, 
    0.975465483762878, 0.976677932617177, 0.977960679815547, 
    0.979054044861913, 0.980102373724611, 0.981125495757618, 
    0.982106894715365, 0.983002254901624, 0.983787749734451, 
    0.984655927322597, 0.985442770759103, 0.986082496453658, 
    0.986796366922336, 0.987477535475758, 0.98813929617312, 0.98870204670118, 
    0.989269154076845, 0.989835707075977, 0.990304050044709, 
    0.990812481841969, 0.991264858764375, 0.991733097372639, 
    0.992127804683021, 0.992580257782544, 0.9929802456718, 0.993358291261404, 
    0.99371634706413, 0.994052254455942, 0.994401653585871, 
    0.994729055823805, 0.995023915356485, 0.995341895074702, 
    0.995624550655447, 0.995899248350651, 0.996165687971825, 
    0.99642852455539, 0.996670428091206, 0.996904135724194, 
    0.997145693126095, 0.997359441261007, 0.997574161619239, 
    0.997780236947161, 0.997978071044521, 0.998176789749934, 
    0.998352848447458, 0.998538617928744, 0.998714929018578, 
    0.998881690366945, 0.999044957567457, 0.999203168514026, 
    0.999355093897147, 0.999506503370132, 0.999651320199236, 
    0.999789994223189, 0.999924951102624,
  0.999932522099177, 0.999813012589097, 0.999690295097023, 0.99956375810174, 
    0.99943198505607, 0.999295687748085, 0.999156553413254, 
    0.999010115996012, 0.998862588264277, 0.998709249019791, 
    0.998550943611079, 0.998384573649704, 0.998205320740535, 
    0.99803801227802, 0.997853267266659, 0.997670687451587, 0.99746513382583, 
    0.997265848037296, 0.997051116002518, 0.99684031305966, 
    0.996611389431294, 0.996386467099792, 0.996122314220324, 
    0.995874125905439, 0.995616201837118, 0.995326132275246, 
    0.995059463979213, 0.994758774907287, 0.994444797030369, 
    0.994103801187329, 0.99378223865113, 0.993420928305354, 
    0.993085104390459, 0.992697509128682, 0.992270706174623, 
    0.99187402453009, 0.991424538079873, 0.990954205331991, 
    0.990514817796623, 0.989959493100547, 0.989457656717914, 
    0.988919604304662, 0.988362506673778, 0.987729751204878, 
    0.987073077348737, 0.986409359400163, 0.985659484844101, 
    0.984923656531015, 0.984164464947446, 0.983311322997954, 
    0.982386965210602, 0.981429146324529, 0.980429673063104, 
    0.979315060302326, 0.978307143636551, 0.976979267058347, 
    0.975706410621633, 0.974231237140827, 0.972807708403987, 
    0.971250397290052, 0.969642732624233, 0.967775764119967, 
    0.965707478812549, 0.963655480680001, 0.96125034816021, 
    0.959010986172654, 0.956179034224054, 0.953128428807808, 
    0.949834944848519, 0.946298642095474, 0.942651013133725, 
    0.938126596452606, 0.933734990633991, 0.928493337454235, 
    0.922978499736295, 0.916854175207745, 0.909959451981046, 
    0.901864718587472, 0.893266253422424, 0.883262403326096, 
    0.872226325395702, 0.859481613376593, 0.845462939152995, 
    0.828936518574683, 0.809880493857175, 0.787373508479711, 
    0.763220621589403, 0.733131559707855, 0.69911573396521, 
    0.658305132079001, 0.611115592934823, 0.557081956032996, 
    0.492923505948242, 0.423907097290025, 0.342893386162406, 
    0.259355563621793, 0.174409755164743, 0.0975230346023464, 
    0.0370576532636183, 0.00450893376990664, 0.00416666108012863, 
    0.0375031650975481, 0.0984327405406282, 0.175415541801107, 
    0.260791853161579, 0.343053588981871, 0.424237389238896, 0.4959008319981, 
    0.556687823331406, 0.611844480763556, 0.658183923026222, 0.6973589525719, 
    0.732929210653798, 0.762945493513499, 0.787998503908358, 
    0.809314628428321, 0.827952128346517, 0.844989426660308, 
    0.859911544377987, 0.87191159083133, 0.883288554457088, 
    0.893143971040107, 0.902247345121208, 0.909630023027058, 
    0.91688024257478, 0.923344284358436, 0.928812782809041, 
    0.933832943261082, 0.938504200754929, 0.942771703027929, 
    0.94641131069028, 0.949829008557168, 0.953017588543892, 0.95604471551337, 
    0.958737138221061, 0.961271000532393, 0.963662793788692, 
    0.965747851158024, 0.967652425986488, 0.969582186030229, 
    0.971302089900928, 0.97282131782801, 0.974276452779105, 
    0.975677695866958, 0.976988774115399, 0.978235098409709, 
    0.979364215710188, 0.980374544826585, 0.981436025567572, 
    0.982303483248427, 0.983276784821804, 0.984126300076019, 
    0.984900985974629, 0.985710396821089, 0.986419560071577, 
    0.987073616943287, 0.987751639158232, 0.988294905967315, 
    0.988949893420496, 0.989469926145555, 0.989967076337263, 
    0.990479640346769, 0.990972094833251, 0.991445658743706, 
    0.99187042350867, 0.992288368785034, 0.992659014487975, 0.99305237080162, 
    0.993451256833602, 0.993778723714249, 0.994142413830203, 
    0.994456845585039, 0.994734893851788, 0.995067636471225, 
    0.995336690012203, 0.995612174410944, 0.995877830871706, 
    0.996123611538906, 0.996374027147813, 0.996600073504635, 
    0.996836956060745, 0.997049595390141, 0.997255019279059, 
    0.997466158248257, 0.997669265628439, 0.997852823806044, 
    0.998040188614639, 0.998210881965178, 0.998390163083803, 
    0.998549903972194, 0.99870576996272, 0.998859831755826, 
    0.999016681042024, 0.999156969686377, 0.999294979477328, 
    0.999429033846619, 0.999561712931844, 0.999689805810549, 
    0.999812918916885, 0.99993261732152,
  0.999938673374332, 0.999832291255377, 0.999720664352052, 0.99960788243848, 
    0.999489189066317, 0.999367846725875, 0.999239413792313, 
    0.999111820947107, 0.99897862795165, 0.998838465278745, 
    0.998698941956356, 0.998551416231679, 0.998394348406557, 
    0.998240066568218, 0.998081262272252, 0.997898171899182, 
    0.99772809576215, 0.997542827716562, 0.997354091939801, 
    0.997161220649268, 0.996958279278196, 0.996736112607482, 
    0.996526539684181, 0.996302012321272, 0.996080809263393, 
    0.99581995214706, 0.995565529431939, 0.995294200340048, 
    0.995022304702304, 0.994721258756587, 0.994424387204306, 
    0.994121971905232, 0.993796423258305, 0.993451439660071, 
    0.99308513505987, 0.992726682655158, 0.992330024347368, 
    0.991960703094096, 0.99147369782492, 0.991011219662621, 
    0.990541056643573, 0.990073092430383, 0.989529536099449, 
    0.988955877978219, 0.988411921131268, 0.987832321368808, 
    0.987148428500614, 0.986507057359111, 0.985729698475302, 
    0.984962563537624, 0.9841924751011, 0.983316892678111, 0.982382303774026, 
    0.981391322107835, 0.980404433045169, 0.979349855958204, 
    0.978157719108435, 0.976902352018785, 0.975599765655789, 
    0.974143157336028, 0.972548809481869, 0.970832776594778, 
    0.969159973293235, 0.967222952634284, 0.965074374555847, 
    0.962803994538792, 0.960437968649617, 0.957852030121001, 
    0.954860574868822, 0.951614215058679, 0.948145098627005, 
    0.944468687306931, 0.940449686476327, 0.935696651182917, 
    0.930426645539724, 0.924646701285872, 0.918428166665553, 
    0.911365743320174, 0.903002839222887, 0.894302290779745, 
    0.884349431197637, 0.872093361291636, 0.858909106688183, 
    0.843716158923712, 0.826541289458933, 0.805754389168752, 
    0.781828261272268, 0.753579135899943, 0.720006912588451, 
    0.682605205650679, 0.636867576840888, 0.584345574313452, 
    0.521573505929661, 0.44894817187191, 0.369541907400989, 
    0.281386206257767, 0.192891368468498, 0.107517575988351, 
    0.0423913874583109, 0.00435216208319102, 0.00465622246516804, 
    0.0419191996081212, 0.107562522410078, 0.18976685648975, 
    0.281983871550649, 0.370688850569895, 0.447475047015141, 
    0.520994495912842, 0.582842537120928, 0.63550951389976, 
    0.683086271380052, 0.721009436076517, 0.753284213496748, 
    0.781328102962829, 0.804784106225869, 0.82603813191827, 
    0.843553106158793, 0.858473979108107, 0.872463050176977, 
    0.88352858610526, 0.893717168031997, 0.903248370096831, 
    0.911478596004191, 0.918167236813372, 0.924732979914604, 
    0.930655181714711, 0.935632783772179, 0.940048453582914, 
    0.944488580041475, 0.948382448939627, 0.951712047324319, 
    0.954877898084248, 0.957825187086207, 0.960432796335685, 
    0.96298117841406, 0.965252734448414, 0.967170973062534, 
    0.969196111338425, 0.97092129961887, 0.972569197427792, 
    0.974138616612298, 0.975528884521258, 0.976950606146501, 
    0.978152921886884, 0.979342574573687, 0.980333163675756, 
    0.981466493829538, 0.982371293966865, 0.983330104050038, 
    0.984114914064689, 0.984988743434441, 0.985680140160133, 
    0.986474101592803, 0.987173788723212, 0.987758466746238, 
    0.988450274167048, 0.988976293540246, 0.989491290631308, 
    0.990038742765026, 0.990559627829571, 0.99101260590413, 0.99148216660968, 
    0.991929857662958, 0.992358040313027, 0.992728225461746, 
    0.993096409441104, 0.993436560293166, 0.993771702805189, 
    0.994125066198893, 0.994408153313856, 0.994749707706564, 
    0.995011877874693, 0.995299006238261, 0.995571320326937, 
    0.995814493792093, 0.996066881554771, 0.99629169435511, 
    0.996528255843729, 0.996753556675134, 0.996955292730014, 
    0.997160802494115, 0.997358466170612, 0.997540520437821, 
    0.997724601454748, 0.997901384112185, 0.998070921052053, 
    0.998239153433628, 0.998395397841002, 0.99854828397523, 0.99869946958136, 
    0.998840125855344, 0.998980418029648, 0.99911540595384, 
    0.999238274462222, 0.99936906645222, 0.999490324018326, 
    0.999608463610899, 0.999721210324556, 0.999831911852014, 0.999938845135033 ;

 ens_sizes = 5, 6, 7, 8, 9, 10, 12, 14, 15, 16, 18, 20, 22, 24, 28, 30, 32, 
    36, 40, 44, 48, 49, 50, 52, 56, 60, 64, 70, 72, 80, 84, 88, 90, 96, 100, 
    120, 140, 160, 180, 200 ;
}
