netcdf filter_ics.0012 {
dimensions:
	domain_size = 40 ;
variables:
	double state(domain_size) ;
		state:units = "none" ;
	int dart_days ;
		dart_days:long_name = "days" ;
		dart_days:calendar = "no calendar" ;
		dart_days:units = "days since 0000-00-00 00:00:00" ;
	int dart_seconds ;
		dart_seconds:long_name = "seconds" ;
		dart_seconds:calendar = "no calendar" ;
		dart_seconds:units = "seconds since midnight" ;

// global attributes:
		:DART_file_information = "dart output member 12" ;
		:DART_creation_date = "YYYY MM DD HH MM SS = 2016 11 22 09 26 08" ;
		:DART_source = "$URL: https://svn-dares-dart.cgd.ucar.edu/DART/branches/rma_trunk/io/direct_netcdf_mod.f90 $" ;
		:DART_revision = "$Revision: 10669 $" ;
		:DART_revdate = "$Date: 2016-08-29 11:16:35 -0600 (Mon, 29 Aug 2016) $" ;
data:

 state = -3.09036060587693, 2.81639812796183, 5.34211924078629, 
    5.23007480614553, -1.21508873154863, 1.91781539737189, 5.76225453832611, 
    5.48882930669238, -4.90825973729457, 4.94497079278637, 4.86678367613598, 
    3.1090291436312, 6.3055614876701, 4.20027619178106, 1.31667672547683, 
    3.86618711690635, 2.90727714151562, -2.05343786903775, 2.00625312394755, 
    2.47659560157469, 8.25043273780088, -1.75575943161926, -1.40581862798915, 
    1.8077663634748, 3.10567864062924, 3.73182111645618, 6.07156946325131, 
    -3.32964775514527, -0.587074386417673, -2.35282845210724, 
    8.60614408523951, 1.7450800512675, 0.958885278940814, 1.56295965695102, 
    3.53002720318004, 7.81638926728432, 0.827060410710333, 2.73378026516193, 
    6.31445660515181, 5.81340549669425 ;

 dart_days = 41 ;

 dart_seconds = 57600 ;
}
