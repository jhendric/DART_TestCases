netcdf atmos_coupled.res {
dimensions:
	xaxis_1 = 1 ;
	xaxis_2 = 144 ;
	yaxis_1 = 1 ;
	yaxis_2 = 90 ;
	zaxis_1 = 1 ;
	Time = UNLIMITED ; // (1 currently)
variables:
	float xaxis_1(xaxis_1) ;
		xaxis_1:long_name = "xaxis_1" ;
		xaxis_1:units = "none" ;
		xaxis_1:cartesian_axis = "X" ;
	float xaxis_2(xaxis_2) ;
		xaxis_2:long_name = "xaxis_2" ;
		xaxis_2:units = "none" ;
		xaxis_2:cartesian_axis = "X" ;
	float yaxis_1(yaxis_1) ;
		yaxis_1:long_name = "yaxis_1" ;
		yaxis_1:units = "none" ;
		yaxis_1:cartesian_axis = "Y" ;
	float yaxis_2(yaxis_2) ;
		yaxis_2:long_name = "yaxis_2" ;
		yaxis_2:units = "none" ;
		yaxis_2:cartesian_axis = "Y" ;
	float zaxis_1(zaxis_1) ;
		zaxis_1:long_name = "zaxis_1" ;
		zaxis_1:units = "none" ;
		zaxis_1:cartesian_axis = "Z" ;
	double Time(Time) ;
		Time:long_name = "Time" ;
		Time:units = "time level" ;
		Time:cartesian_axis = "T" ;
	double glon_bnd(Time, zaxis_1, yaxis_1, xaxis_1) ;
		glon_bnd:long_name = "glon_bnd" ;
		glon_bnd:units = "none" ;
	double glat_bnd(Time, zaxis_1, yaxis_1, xaxis_1) ;
		glat_bnd:long_name = "glat_bnd" ;
		glat_bnd:units = "none" ;
	double dt(Time, zaxis_1, yaxis_1, xaxis_1) ;
		dt:long_name = "dt" ;
		dt:units = "none" ;
	double lprec(Time, zaxis_1, yaxis_2, xaxis_2) ;
		lprec:long_name = "lprec" ;
		lprec:units = "none" ;
	double fprec(Time, zaxis_1, yaxis_2, xaxis_2) ;
		fprec:long_name = "fprec" ;
		fprec:units = "none" ;
	double gust(Time, zaxis_1, yaxis_2, xaxis_2) ;
		gust:long_name = "gust" ;
		gust:units = "none" ;

// global attributes:
		:filename = "RESTART/atmos_coupled.res.nc" ;
data:

 xaxis_1 = 1 ;

 xaxis_2 = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 107, 
    108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 121, 
    122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 
    136, 137, 138, 139, 140, 141, 142, 143, 144 ;

 yaxis_1 = 1 ;

 yaxis_2 = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90 ;

 zaxis_1 = 1 ;

 Time = 1 ;

 glon_bnd =
  144 ;

 glat_bnd =
  90 ;

 dt =
  1800 ;

 lprec =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2.06907663231558e-11, 2.24267529545436e-10, 0, 
    5.09373001176089e-11, 1.82714001063787e-10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 1.35183041349667e-10, 2.13715890391799e-10, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1.14048837141679e-09, 0, 0, 0, 0, 0, 0, 9.3644065557776e-14, 0, 0, 
    0, 0, 0, 0, 0, 0, 9.00751317420348e-12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9.71508722186967e-12, 5.28973694382363e-11, 1.35745132298535e-10, 0, 
    1.80435705219136e-10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 7.87254746073077e-12, 2.23741556061264e-10, 
    3.42823524054816e-10, 1.11046277413218e-10, 1.14633964722494e-10, 
    2.3183439036176e-11, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8.10610420441251e-11, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.35053153237877e-11, 
    3.96308409941191e-10, 3.11895472593008e-11, 0, 0, 0, 0, 0, 0, 
    5.25002471502178e-13, 6.21280325183436e-12, 1.07923796905985e-12, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5.77433228044009e-11, 6.19626573775271e-12, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.80719896230297e-11, 0, 0, 0, 
    0, 0, 0, 0, 0, 2.31035253520411e-13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.45441853276904e-11, 
    1.15151239120455e-10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6.94756948035979e-12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.19103850199747e-12, 
    0, 0, 0, 0, 0, 0, 0, 2.26941126151096e-11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1.58235420710376e-14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.66149700949812e-11, 3.1553572385361e-11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1.16590680784222e-10, 2.39582008778893e-09, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 5.42013048693896e-13, 1.16655776270519e-11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.10280569315881e-11, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.3543068775463e-12, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  5.25912348706847e-11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.11671190242632e-12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.67712185870478e-11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4.29064615108784e-11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 4.24441575604564e-10, 0, 9.26793634802552e-12, 
    1.53440821171302e-10, 6.61786389427519e-11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4.03870584397031e-12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6.00029255467927e-13, 0, 9.66847498529989e-10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5.28346048173684e-11, 0, 4.40435469972205e-10, 0, 
    4.88958925769064e-13, 0, 0, 0, 0, 0, 8.53177287499202e-07, 0, 0, 0, 0, 0, 
    0, 0, 1.06036124699771e-10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8.92252341102227e-18, 0,
  0, 0, 0, 0, 0, 0, 2.09616619371837e-11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.99028762623319e-11, 0, 
    8.78919962495082e-09, 0, 0, 0, 0, 0, 2.28906575513641e-10, 
    4.14868443709706e-12, 0, 0, 0, 0, 0, 0, 1.5363333395391e-05, 
    6.15144283034124e-05, 4.65504547300504e-05, 4.53051601047829e-05, 
    5.87798132220544e-05, 3.95286349238915e-05, 0, 0, 0, 0, 0, 
    1.6145347982649e-10, 0, 0, 0, 9.84634920362747e-12, 1.81400550838003e-10, 
    0, 0, 0, 1.96903210661987e-10, 4.38798120588402e-13, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.97151927929077e-14, 0,
  1.08476012364341e-12, 0, 0, 7.67259068768038e-09, 3.48360579369781e-10, 0, 
    1.35465035207019e-10, 4.61450541259174e-10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.58668407390639e-10, 
    2.01902914121186e-09, 1.79199642530073e-10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4.0993739370224e-05, 0.000168129929474686, 8.89843257832692e-05, 
    4.30237903443464e-05, 1.20679416006866e-05, 4.78511436569992e-06, 
    5.49386115183584e-06, 5.98646707698567e-06, 1.10561651293749e-05, 
    5.36562182880928e-05, 0, 0, 0, 0, 9.1707417711658e-09, 
    1.99617545868669e-11, 0, 0, 9.13749947889105e-12, 0, 
    4.77077628195039e-12, 0, 1.15969838472846e-11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5.71749600935497e-11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.27203962689813e-11,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.80383996911873e-08, 
    1.63842716797804e-10, 0, 0, 0, 0, 0, 0, 0, 1.28531875655556e-11, 0, 
    5.48645175811233e-07, 0, 0, 0, 0, 0, 0, 9.59714262087129e-10, 
    9.79887591501396e-13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.49533351653071e-12, 
    0, 0, 0, 0, 0, 0, 4.67770201341882e-11, 1.10563116450363e-11, 0, 0, 0, 0, 
    4.65159392650534e-11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.93375367927634e-05, 
    0.000223639795867035, 0.000242107981750432, 9.66396464002553e-05, 
    9.75697141764301e-06, 6.83354219098608e-06, 2.83327202770739e-06, 
    1.88504893335288e-06, 1.40270770841271e-06, 3.07577587160911e-06, 
    4.23445470227598e-06, 5.66937480369549e-06, 1.47935262610494e-05, 
    2.08662933706146e-05, 1.70091035860203e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2.41357153670958e-10, 0, 4.99603585044455e-16, 0, 0, 0, 0, 0, 
    6.65645737659607e-08, 3.23367506409288e-08, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.87560689213391e-08, 
    1.53988314534903e-08, 5.47442256444165e-08, 9.09085913742043e-08, 
    9.4992589993378e-08, 1.45467684066275e-08, 7.5722412339438e-08, 
    1.84343977513211e-08, 1.81656758163755e-09, 1.04284081734123e-11, 0, 0, 
    1.09471967581925e-09, 1.08235240185591e-11, 0, 5.2912514421001e-09, 
    3.3869709736012e-09, 5.10869039662557e-07, 2.67058609824909e-06, 0, 0, 0, 
    0, 1.49735350858827e-10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.87495494513641e-10, 
    9.76211067557866e-10, 1.15993082004033e-08, 1.25877089238184e-09, 
    8.04251933210847e-10, 5.68853310115284e-08, 2.60862823774542e-07, 
    1.3913481761613e-06, 1.3874324053812e-05, 8.32542165564415e-05, 0, 0, 0, 
    0, 0, 0, 0, 1.58666312162198e-10, 0, 0, 9.55001513327058e-09, 
    1.90971694301913e-09, 0, 0, 0.000439158978792203, 0.000448350558955531, 
    0.000304214807917334, 6.28997560314322e-05, 6.73096477918321e-06, 
    5.40686152605084e-06, 6.05702188876507e-07, 4.36627373507556e-07, 
    3.57360606794045e-07, 5.05827325392536e-07, 9.91414433441069e-07, 
    3.33732066862582e-06, 1.68178199864494e-06, 2.47683665373984e-06, 
    6.78607355093915e-06, 2.27922818856677e-05, 1.61691689149526e-05, 0, 
    1.04195855827378e-08, 0, 6.46550909319045e-09, 0, 0, 0, 0, 0, 0, 
    7.35647790016666e-10, 1.94638728463828e-10, 0, 0, 0, 0, 0, 0, 0, 
    2.61879225877336e-07, 3.07476295384276e-08, 0, 1.07070357705862e-09, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 3.86028155200704e-11, 9.7398706764341e-09, 6.06755242410953e-08, 0, 
    6.53617728164721e-09, 2.86155859227203e-10, 0, 0, 0, 0, 0, 0, 0, 0, 
    9.43544864450404e-09, 3.27447197821976e-08, 9.75815889818379e-08, 
    2.94640997147087e-08, 1.04632463226346e-07, 1.74495944374756e-07, 
    1.42369380436471e-07, 5.36346168462154e-08, 1.12357510188997e-08, 0, 0, 
    3.3226628330325e-11, 1.52752081347619e-10, 1.58749735743845e-07, 
    1.87082825789761e-08, 2.50065232021183e-10, 2.41309884686015e-08, 
    6.325046477455e-08, 2.52613119286945e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1.20131392559543e-08, 6.52277575368069e-08, 
    2.48878941592534e-11, 9.04479618035819e-12, 0, 7.02445597413296e-08, 
    1.22240777942819e-06, 2.86640264942254e-06, 5.33252045426324e-06, 
    6.03213878812144e-05, 0.000208083732964519, 0, 0, 2.01423593826237e-08, 
    1.02148697775327e-08, 8.18923415792706e-09, 5.54831851452319e-08, 0, 
    5.20796418190535e-08, 9.78455731263012e-09, 5.73518113325291e-11, 0, 
    0.000394773657585881, 0.000426791438925945, 0.000267090320115656, 
    2.53908030921098e-05, 4.34541239636867e-06, 8.97012949662622e-07, 
    3.2344547427118e-07, 2.19772724165425e-08, 6.9103926522883e-09, 
    1.03363511395999e-10, 8.32339726050135e-09, 1.17377282404408e-11, 
    4.32999729818411e-08, 1.20028364383903e-07, 2.88384510530232e-07, 
    1.38955052740522e-06, 3.6017174735058e-06, 3.85986360997483e-06, 
    6.31996019730426e-06, 1.77439292689836e-06, 1.43797166421883e-07, 
    9.39574201318599e-08, 4.70210954158105e-08, 0, 0, 0, 0, 0, 0, 0, 
    2.22716206676426e-12, 0, 0, 0, 8.77344807005297e-09, 0, 
    4.31874913478588e-09, 0, 0, 0, 2.79870376303762e-12, 0, 0, 0, 0, 0, 
    2.24484868604436e-08, 0, 0, 0, 1.4819909447463e-10,
  0, 0, 0, 0, 1.29028621050491e-10, 4.70188643604061e-10, 0, 
    5.82494864059392e-09, 1.23542339285533e-08, 1.80722129415544e-08, 0, 0, 
    1.54683767456841e-08, 3.94183495818657e-08, 4.53465414834852e-08, 
    5.59934519377333e-09, 4.19107565971255e-11, 1.36579131366855e-09, 
    1.34317745320299e-07, 1.20612777170144e-07, 2.04272626896118e-07, 
    1.62351926026526e-07, 6.10539277866066e-09, 0, 0, 5.12681970396275e-10, 
    5.43152617047126e-09, 1.76407599602304e-07, 0, 0, 0, 0, 0, 
    1.58481090780216e-06, 2.74637309685046e-05, 0, 0, 5.66947569605571e-08, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.5585008912637e-11, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1.56913774340674e-09, 0, 0, 0, 0, 0, 
    1.6240205950683e-05, 3.32675464015229e-06, 4.49187073397403e-08, 
    4.27638085127061e-10, 1.18576718404656e-09, 4.46786817659467e-10, 
    2.94205673015882e-08, 1.10714459988361e-06, 2.40949769915062e-05, 
    2.40806666646451e-05, 3.93987633456488e-05, 0.000145897443836786, 
    5.8730337580458e-05, 0, 1.47016249351692e-08, 1.49917727172271e-08, 
    5.18791046735897e-09, 1.27591025887151e-09, 1.52719721445127e-08, 
    2.24559910536202e-09, 2.18342952024687e-09, 0, 0.00018939019125924, 
    0.000321880598165878, 0.000239230611185298, 3.60986600690697e-05, 
    1.18431948706147e-05, 8.33605853557561e-07, 3.24734067411157e-07, 
    4.58985920650865e-09, 1.08802503113211e-08, 2.21883084874211e-08, 
    2.91037031153911e-08, 8.15258931446439e-07, 5.55729734864961e-07, 
    5.21247816398412e-07, 4.62778982326058e-07, 3.55174054139069e-07, 
    1.60512155550368e-07, 4.33402121030575e-07, 7.42330655338669e-07, 
    2.91099006064907e-06, 5.92425509379985e-06, 2.66359551541342e-06, 
    5.39702055354525e-07, 2.18214637239912e-08, 1.15344225899143e-07, 
    5.27160250030278e-08, 0, 0, 0, 0, 4.00116351961736e-09, 
    3.97594285281753e-10, 0, 1.35558046979226e-07, 0, 0, 0, 0, 
    4.63787366758903e-07, 1.49162217837119e-06, 6.07221537658004e-07, 0, 0, 
    3.59880028199254e-10, 0, 0, 9.62728260383343e-10, 1.17173024413657e-11, 
    0, 1.67705296293815e-11, 0, 0,
  0, 5.50572137932266e-10, 1.09661163487358e-10, 5.67035035389533e-12, 0, 0, 
    0, 6.03612391088968e-09, 2.51183632301234e-08, 6.28879055912998e-08, 
    7.78815865003006e-08, 1.79017571511963e-08, 6.01605789408733e-09, 
    1.44567051211826e-08, 1.10879640604497e-07, 1.33358597250607e-07, 
    1.36092116388316e-07, 3.61110460217633e-08, 2.75512060024367e-07, 
    7.10125526975248e-08, 2.57300278029382e-08, 1.96591295223065e-10, 0, 0, 
    5.23397728810591e-11, 5.33801019156555e-08, 4.2970739043569e-07, 
    2.45506923080486e-06, 1.40448017129784e-05, 5.66518423556529e-05, 
    7.40416858356478e-05, 7.21789311323064e-05, 3.3178905395598e-05, 
    1.71185480219898e-05, 3.82388191625099e-05, 0, 0, 0, 
    1.26444573489109e-07, 0, 0, 0, 0, 8.74047679060611e-09, 
    6.49708088528188e-08, 1.93547711712705e-08, 3.3434885144059e-08, 
    8.33020707213881e-11, 2.51739081239095e-08, 2.01651764360221e-09, 0, 
    5.74186749612584e-07, 2.69110445077826e-08, 1.61223185198611e-09, 
    2.63186711566802e-09, 6.35045989711777e-10, 1.67428005626003e-07, 
    3.77953890811415e-07, 1.85065533177932e-05, 8.70721458102262e-05, 
    0.000101340976011518, 8.21988677907366e-05, 4.08719237883474e-05, 
    9.16229276772229e-06, 3.88543089317702e-07, 1.5166034742443e-07, 
    5.0877212947577e-07, 1.55081244884612e-06, 5.82332158236125e-06, 
    6.12705995146464e-06, 9.46591437483011e-07, 3.54308635748534e-08, 
    6.95239065624295e-11, 5.84724078589752e-10, 1.41371440960829e-09, 
    2.10492560514326e-05, 1.06014170356422e-05, 6.22354269530146e-05, 
    5.26341952026621e-05, 1.10990746915003e-05, 7.8784613459708e-06, 
    4.39767984324243e-05, 0.000158459203705415, 0, 3.56879204253284e-09, 
    1.99833962150203e-08, 6.8531834859746e-08, 1.17624589031407e-07, 
    4.62589451128859e-08, 1.34249939805499e-09, 0, 0, 0.000138143933397376, 
    0.000241869970151557, 0.000140450624438039, 1.89983629724474e-05, 
    8.57925275627602e-06, 4.97534164535367e-06, 6.09685264827104e-08, 
    3.04493297678273e-11, 1.09530929852934e-08, 1.92673000229344e-07, 
    4.18803196366197e-06, 7.08134330369732e-06, 6.58775648199584e-06, 
    1.79011545058698e-06, 6.97470127505348e-07, 1.14919496276452e-06, 
    2.14742336189888e-06, 4.6571099021754e-07, 4.20834357235214e-07, 
    3.54401728486855e-06, 5.96526955472082e-06, 5.58034573127085e-06, 
    7.99207702051612e-07, 2.33925942353496e-06, 3.38884835399364e-06, 
    6.69416273042504e-10, 1.42766519664204e-09, 0, 1.76404569576701e-09, 
    3.67815149997611e-08, 2.65239366771329e-06, 0, 3.79608647635867e-06, 0, 
    0, 8.140997683072e-06, 6.11952575117916e-05, 5.72947480571392e-05, 
    7.94672721139266e-05, 2.03520383528732e-05, 0, 1.10423589281633e-06, 
    4.57421775998165e-09, 0, 4.40394542773725e-06, 4.10402995935443e-06, 
    3.39893158941657e-08, 2.99512252284755e-10, 0, 0, 0, 0,
  0, 0, 0, 2.58371944383306e-10, 0, 0, 0, 0, 5.96515440280353e-09, 
    1.68035525722654e-08, 3.45853196156887e-08, 3.69257712911077e-08, 
    1.36191585770501e-07, 1.44374399987894e-07, 6.99682691076123e-08, 
    1.49958572157504e-08, 1.32254278901151e-08, 3.18647559521186e-08, 
    3.58344672614043e-07, 1.30615855270903e-07, 2.68409364434e-08, 0, 0, 0, 
    4.69365474116538e-09, 1.52310325786258e-06, 6.85844479556107e-06, 
    9.01149471963995e-05, 0.000107987761968477, 9.75387793710201e-05, 
    7.07043191828684e-05, 6.5681093788712e-05, 4.86454617077841e-05, 
    3.07815682304602e-05, 3.77874539024684e-05, 0.000122146732778241, 0, 0, 
    5.84140576414755e-08, 3.0673272067917e-08, 8.36997048749378e-09, 
    3.0148381213405e-10, 6.42469920995172e-09, 3.16048066886809e-09, 
    1.11613401541711e-09, 2.88362214994268e-07, 1.69764541373037e-08, 
    3.2538475953222e-08, 1.99095589559906e-07, 6.49473639134431e-07, 
    2.87401573242137e-07, 7.79371488259829e-08, 2.36693776671164e-09, 
    7.76560278019778e-11, 7.71169057465458e-08, 7.58510475859709e-07, 
    5.53697933840881e-05, 8.71625721835163e-05, 7.98221342733911e-05, 
    5.64821277981737e-05, 4.25741034788569e-05, 4.7074535075023e-05, 
    3.30318017396293e-05, 9.80135831278275e-06, 4.86406132485439e-06, 
    6.28153311792715e-07, 4.88561950369327e-07, 1.79498889321826e-07, 
    1.30922042961047e-11, 6.96374335250916e-09, 3.74675370718646e-05, 
    1.81807148161476e-05, 1.94897141665637e-05, 2.80822145837837e-05, 
    5.18659356162777e-05, 3.1442958565117e-05, 2.84895987956542e-05, 
    2.08683446144297e-05, 1.702618002454e-05, 6.30570458134706e-06, 
    1.67735408794215e-06, 1.63783625828901e-05, 9.6744503044273e-05, 
    5.0073320468207e-05, 0, 3.19833817176858e-07, 4.3661218624783e-08, 
    1.29113983881585e-07, 1.09703165491099e-09, 8.86254236321722e-08, 
    1.08177994971334e-09, 8.11376802987534e-06, 0.000101299618327091, 
    0.000221093357652258, 0.000101982803088115, 1.56031776547801e-05, 
    1.64638057720981e-05, 5.23357629254639e-06, 1.20522994744856e-08, 
    2.52164604347804e-09, 1.25230085123887e-06, 6.89062306343184e-06, 
    1.00476942926954e-05, 9.11782673923028e-06, 5.6776803328531e-06, 
    4.9320108324279e-06, 4.63445169960764e-07, 5.28365753436931e-08, 
    1.79623399677729e-07, 3.11109715265339e-10, 3.86904294270465e-06, 
    1.06519077773751e-05, 9.8867324895224e-06, 1.71031672496478e-05, 
    6.40841917030776e-06, 1.95086649585902e-06, 1.75320483003273e-06, 
    6.22392345602095e-07, 1.21992336005953e-06, 1.12887213366758e-06, 
    7.55633875997372e-07, 2.65244085251977e-06, 4.36170333270217e-06, 
    2.93608867837943e-06, 4.6799742566447e-06, 5.30409609044286e-05, 
    6.91674280073131e-05, 3.65740759479912e-05, 4.15738231512689e-05, 
    0.000155830437129726, 0.000341775773070088, 0.000360063557071754, 
    0.000228574120172713, 3.43689820825814e-05, 1.48620043385892e-05, 
    4.67962933149364e-06, 1.9564378293846e-06, 1.48048571233918e-06, 
    9.3685594616987e-08, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 2.87718857643059e-07, 1.14797960314848e-06, 
    5.07040936431974e-07, 9.05439716325955e-08, 6.44254309449484e-08, 
    6.99008713450461e-08, 3.73705587263625e-08, 1.61764652776263e-08, 
    8.67181040607781e-08, 1.47255436928162e-07, 2.08844010024173e-08, 
    1.27561292894046e-09, 5.78442021776837e-08, 1.37287126815979e-07, 
    3.20431587323953e-07, 2.90417371239236e-07, 4.35775186722495e-08, 
    4.26398097291772e-10, 1.94857865114872e-08, 0, 9.79655880939558e-07, 
    0.000119866144233608, 0.000147680121589864, 0.000120400994445657, 
    5.69111432713204e-05, 3.08223844394482e-05, 1.32238962612251e-05, 
    1.33327681296124e-05, 1.14676268804287e-05, 1.12832266787678e-05, 
    2.05573068585093e-05, 7.32208073769251e-05, 0.000168195860501032, 0, 
    1.57423197748469e-08, 9.70608400185525e-09, 4.667607932091e-09, 
    8.41567786411557e-10, 4.28980522312423e-10, 0, 0, 2.65127174032584e-07, 
    1.61223983748355e-08, 4.78374748385946e-09, 4.19436872383687e-10, 0, 0, 
    5.4362745945393e-11, 3.9245676816423e-08, 6.14394888803774e-06, 
    7.84416402086098e-05, 0.000134205287131067, 0.000120809003078295, 
    5.31370321568039e-05, 1.4770766233322e-05, 5.89232664372691e-06, 
    6.90435756062868e-06, 7.99330520441493e-06, 6.19470474477156e-06, 
    1.0535540884098e-05, 8.40430477027935e-06, 2.76678677710453e-05, 
    3.42163182987134e-05, 5.01302382381637e-05, 2.31172817024839e-05, 
    9.33148186719161e-06, 2.44522317601837e-06, 8.04591526706548e-06, 
    3.55297936695169e-05, 5.12825841053501e-05, 5.8535637399672e-05, 
    4.04000489151241e-05, 1.27690719860201e-05, 3.1091442392281e-06, 
    3.07426238549437e-06, 8.21543406807743e-06, 6.39523547892346e-06, 
    1.21147315758924e-05, 2.80825224512479e-05, 2.8818479849214e-05, 
    1.34449219608265e-08, 2.78276939287974e-07, 4.48158161119271e-08, 
    1.3438762563881e-09, 0, 1.03236210991459e-07, 1.22837718355156e-07, 
    4.43687162776679e-06, 5.63717995802395e-05, 0.000230276694875205, 
    8.33744825346435e-05, 1.62695902343076e-05, 2.32474022110685e-05, 
    3.1584057227237e-06, 2.92312012843224e-08, 3.3035610216599e-09, 
    4.59043399281252e-06, 1.16412189789558e-05, 1.04124982704591e-05, 
    7.86083354558577e-06, 6.78521825292312e-06, 4.48677162925359e-06, 
    2.64508579910843e-06, 1.52762780354266e-08, 1.86701364063093e-07, 
    8.9527057339783e-07, 7.7004732478878e-06, 7.35607494828292e-06, 
    1.30438305015276e-05, 3.8317774825634e-05, 1.41443061279837e-05, 
    8.57515809872358e-06, 4.86060263758682e-06, 1.54642392498909e-06, 
    5.17300179427643e-08, 1.05092283797431e-07, 2.27573226818658e-06, 
    1.18817585866754e-06, 3.02520120287898e-06, 4.30927234029495e-06, 
    4.22502511000195e-05, 3.58512888644562e-05, 1.56700434709951e-05, 
    8.9016867411265e-06, 1.57939271132103e-06, 3.91149446572923e-06, 
    0.000107494801076681, 0.000444962325833569, 0.000415016357368427, 
    0.000196916754558142, 1.4306336889673e-06, 2.50630130265107e-06, 
    6.58805937269168e-08, 1.60840936731982e-07, 6.01768521726561e-08, 0, 0, 
    0, 0, 0,
  3.50589159877895e-05, 9.84989815904277e-05, 8.7055058936261e-05, 
    2.87293735586281e-05, 3.10633761136106e-05, 2.66584093318462e-07, 
    3.89449760638503e-07, 5.49546059000163e-08, 6.18422481435468e-09, 
    9.96777004313256e-08, 1.65732908986118e-08, 5.95032169824661e-09, 
    3.87092761734829e-09, 1.01143037121666e-07, 2.57706434958391e-08, 
    5.34712010536805e-08, 1.08922437148903e-07, 1.06652821112942e-07, 
    1.01766255327398e-07, 6.51436233715207e-15, 2.37081703585629e-08, 
    1.91000748726336e-12, 4.51842064098306e-07, 0.000139439657211102, 
    0.000242938975922837, 0.000219448609066078, 9.6748963735693e-05, 
    2.87090580683277e-05, 4.185505225064e-06, 7.48808670902762e-06, 
    5.56309819442839e-06, 2.59734039114579e-06, 5.3756445680354e-06, 
    6.6049769136762e-06, 9.53964086778037e-06, 2.81664739093256e-05, 
    0.00013847559654808, 0.000154233034965604, 0, 3.05139129611216e-07, 
    8.33728606335762e-09, 0, 0, 0, 0, 9.14869569439153e-08, 
    6.29651418877686e-08, 5.30636163409644e-09, 2.08306083829751e-08, 
    4.37454751704096e-09, 2.58978767878888e-13, 1.10602574060168e-05, 
    0.000125312733365147, 0.000161624792208333, 8.48616545302964e-05, 
    1.55666065878981e-05, 3.77251000695185e-06, 1.57141560833919e-06, 
    4.38090082971765e-06, 6.2251925430014e-06, 4.12836740305671e-06, 
    2.83704423123454e-06, 2.8254982816149e-06, 6.71506056370824e-07, 
    7.52507997250372e-06, 1.02007325210836e-05, 7.44413577118449e-06, 
    2.76507920688685e-06, 3.22076276737332e-07, 1.24464895904489e-06, 
    3.23808092104885e-06, 1.53754735687425e-05, 3.95078265566099e-05, 
    3.2967137002074e-05, 1.23450344362698e-05, 6.06723265615455e-06, 
    2.22263401885492e-07, 5.23398488489663e-07, 6.69401763474072e-06, 
    1.03424302937502e-05, 4.19916228358455e-06, 2.02930600904227e-05, 
    1.2214039292974e-05, 1.11715620329787e-05, 1.43305230023396e-06, 
    2.56888756053208e-07, 2.92589768569896e-08, 7.08486066698623e-13, 
    4.22521427149713e-08, 2.41920804221237e-08, 5.94197323191174e-07, 
    3.02034581370493e-06, 3.09436397888116e-05, 0.000256034109994141, 
    4.30269529620438e-05, 2.11086588474133e-05, 2.2462586332113e-05, 
    7.2914009473582e-06, 1.09677508796339e-06, 3.17768935636783e-08, 
    1.45535187616753e-06, 1.25970751718247e-05, 1.25743930648863e-05, 
    5.40590823801125e-06, 7.2610710229932e-07, 2.634603023734e-06, 
    3.86706539378805e-06, 2.06484549976172e-06, 6.22842856545689e-07, 
    3.03096085406358e-07, 2.02141789240901e-05, 1.21835289437329e-05, 
    1.65091393681863e-05, 3.17832137641149e-05, 6.0642292029656e-05, 
    3.49047143909473e-05, 4.84776476810268e-06, 7.12030366702814e-07, 
    3.40856745372435e-07, 5.58143776480286e-08, 2.95606401475644e-06, 
    6.47292961410419e-07, 2.59402979062377e-06, 2.28012665221754e-05, 
    7.93943584549196e-06, 1.00166762518409e-05, 1.06772388591078e-05, 
    7.09879208858139e-05, 9.50547251155599e-06, 2.43385799834762e-07, 
    4.03094261948557e-07, 0.00023650865163028, 0.000532174711010306, 
    0.000339904039742793, 1.12710088072198e-05, 7.14011128051052e-08, 
    3.6227035122505e-07, 4.6514672687019e-07, 2.50537878946266e-07, 
    1.10313222091351e-06, 8.71969209473674e-07, 0, 5.14544113430323e-06, 
    2.29284682412325e-05,
  5.06092483725684e-06, 8.09595363873112e-06, 5.98416844670382e-05, 
    0.000378574682122784, 0.000182427481067779, 1.09198466865628e-05, 
    2.10149293767374e-07, 1.1475368196322e-06, 6.35175555647276e-07, 
    4.18740972458376e-08, 2.37948490797677e-07, 2.09613584192309e-07, 
    2.53289369454557e-07, 1.66899777979516e-08, 1.09463106012251e-09, 
    8.24648674056245e-11, 1.7354713807464e-11, 5.29177209508614e-11, 
    3.6098345621244e-17, 0, 0, 1.15839163879973e-05, 0.000277068294640821, 
    0.000331883289822418, 0.000174083175980997, 5.14536154738672e-05, 
    6.38174601149508e-06, 3.30880785046123e-07, 1.75147157015507e-07, 
    3.79558648044332e-07, 7.89477127593033e-06, 5.81811630661583e-06, 
    4.10107720692063e-06, 5.25604282865055e-06, 6.7102959973679e-06, 
    1.85480476000078e-05, 8.52469810168283e-05, 0.000168325927431996, 
    4.67925381201745e-05, 1.67666378452505e-07, 3.68414770106882e-08, 0, 0, 
    2.24604071234268e-07, 5.23520667146504e-07, 1.30196922341609e-06, 
    2.83283900133861e-07, 1.34983924463178e-09, 2.00811507858116e-10, 
    6.82021338381792e-08, 7.0437844098324e-05, 0.000203076151675388, 
    0.000126550275295137, 2.78428725334914e-05, 3.00685024390737e-06, 
    1.25497738278692e-08, 2.65789750219767e-10, 5.67454296796961e-11, 
    8.82825653346804e-12, 1.63820433263455e-06, 1.96031676997987e-07, 
    3.67934504212804e-06, 1.84603959962105e-23, 1.67922616819029e-06, 
    1.46900528161161e-06, 1.19824996505145e-07, 4.92317767903489e-20, 
    6.23018223199817e-06, 3.54015256938405e-06, 4.84864399627313e-05, 
    5.83806877878133e-05, 4.08809260149828e-05, 2.06284385396022e-06, 
    1.88577152104275e-07, 5.28164976345483e-06, 1.4045727116258e-05, 
    4.40606772393712e-06, 7.88466824702456e-06, 5.75746532602368e-06, 
    6.38447295425628e-06, 9.23599626726623e-06, 1.32978658793975e-05, 
    2.34013019233798e-05, 4.26792761309792e-06, 1.78766132083541e-06, 
    3.30014663747359e-08, 2.32856290854085e-09, 8.22376080788914e-08, 
    8.79121159879229e-13, 1.06906258050578e-07, 1.23652047231549e-06, 
    3.04888074887386e-06, 2.40688656888483e-05, 0.000282401656113566, 
    2.86405660705855e-05, 2.29426393519842e-05, 1.76942685836463e-05, 
    1.24654655145329e-05, 8.55069039928425e-06, 1.10786338552348e-06, 
    2.62248473636121e-11, 9.91000595855035e-06, 1.17880081250453e-05, 
    9.75611441523329e-06, 1.6848580405995e-06, 1.35279438371539e-06, 
    1.31467933517177e-06, 3.75995774644589e-06, 2.40842538295301e-08, 
    2.76377195911742e-06, 5.16105622922989e-06, 7.45663462008722e-06, 
    2.39266059433535e-05, 8.81008970444709e-06, 0, 0, 2.5623716356217e-07, 
    8.38618358526252e-07, 3.49186216921349e-07, 1.93617488365406e-06, 
    4.9463301696769e-06, 3.79816700406661e-07, 3.84967429379951e-06, 
    2.20111609217062e-05, 2.7682692190827e-05, 1.61433600877735e-05, 
    0.000101577628840996, 0.00010632918769197, 9.37376901885913e-05, 
    2.04083594089995e-07, 8.5706841352064e-09, 4.29617401844258e-05, 
    0.000451047010218628, 0.000434000503116494, 6.09489056804044e-05, 
    8.20278004734079e-08, 9.08106882149336e-07, 6.28685305512378e-07, 
    7.87262644729037e-07, 1.22791069381623e-06, 7.21163533133376e-07, 
    3.0153882313393e-06, 3.45000464614887e-06, 9.04541753256467e-06,
  7.48252179625589e-05, 1.13306327585968e-05, 4.70845882317158e-05, 
    8.92232052134324e-05, 0.000484157685802455, 0.000332090964201719, 
    7.46223083711558e-07, 1.54086899026179e-06, 1.42403154955137e-06, 
    6.45828857979896e-07, 1.18416612813351e-07, 2.84451742815523e-08, 
    3.95217218369591e-07, 2.30615010308807e-08, 5.17183769312662e-13, 
    7.83023481289793e-15, 0, 7.03975602308816e-18, 4.43549377641092e-13, 0, 
    0.000188172343133607, 0.000475201074215314, 0.000383398233274688, 
    9.96154658833094e-05, 2.22030384957402e-06, 7.89567804656237e-08, 
    9.63474564263292e-09, 9.39222549948962e-08, 1.02413911734779e-06, 
    3.71497086116362e-06, 2.88465805374369e-06, 1.4162183470236e-06, 
    7.32874238647677e-07, 1.1676258276246e-06, 1.74901074593406e-06, 
    3.63026256729484e-06, 2.71585675527038e-05, 9.08418392622876e-05, 
    4.45097779291931e-05, 3.34928717815089e-06, 1.23978394212849e-07, 
    6.49001598082669e-09, 1.23043488432561e-13, 4.92677800208764e-08, 
    6.98422926571751e-07, 7.69197997084349e-07, 3.05948686487655e-08, 
    3.19249192721553e-09, 7.41504346346513e-08, 0.000105554054532265, 
    0.000147104505876627, 9.99202558506577e-05, 1.99614011140431e-05, 
    2.02090077839416e-05, 1.20460919189874e-05, 2.58056500130957e-06, 
    7.31448952950232e-06, 4.49086372485851e-06, 2.92471482260125e-06, 
    3.54419385089336e-06, 2.60583691245674e-06, 2.84036429449477e-06, 
    4.17015461731957e-07, 0, 1.17624251525356e-12, 2.96773251841617e-06, 
    3.44719927753909e-05, 5.43465916648355e-05, 3.64552491210799e-05, 
    3.31531911171902e-05, 3.57008738044691e-20, 6.46477110252892e-09, 
    1.44150879841428e-09, 9.64557979111081e-06, 3.59532880981202e-06, 
    8.3351123730153e-06, 7.11399506480285e-07, 4.35132832034381e-06, 
    3.94764433296163e-06, 3.47992923944117e-06, 5.03309278946211e-06, 
    2.10247070720093e-05, 1.7768521406046e-05, 2.48215694648841e-06, 
    1.59995527314629e-07, 1.30950371952846e-08, 5.76375025520011e-12, 
    8.30338309756296e-13, 9.60927647875064e-08, 5.003270382966e-07, 
    5.41798424542355e-06, 9.77531438660044e-07, 1.40445839763588e-05, 
    0.00030280917672924, 3.32261957180547e-05, 4.72048231646585e-06, 
    1.04832215995878e-05, 1.01429612710867e-05, 1.77406228880187e-05, 
    1.78564986477243e-05, 1.56589744342524e-05, 1.17518847714278e-06, 
    4.0196823482466e-06, 2.02721176971021e-06, 6.15613820818883e-06, 
    4.3452445579625e-06, 8.81366759456134e-07, 1.2306213547852e-06, 
    4.31215103017584e-06, 1.64878846505826e-06, 6.58575593642427e-06, 
    1.83662273498046e-05, 2.5935449206562e-05, 2.15779233299884e-05, 
    5.84400744956898e-09, 0, 4.60376459694224e-10, 8.799700205258e-12, 
    1.13227615016893e-07, 2.13901536021402e-06, 3.80639009365751e-06, 
    4.51463346485923e-07, 6.18607400340235e-06, 6.29868385740353e-05, 
    6.21196830046205e-05, 5.22218388762385e-05, 6.46031182351605e-05, 
    0.000123583531122279, 1.70037657825672e-05, 1.32170382672742e-08, 
    1.59790235583851e-07, 6.2977095233072e-05, 0.000393258148665622, 
    0.000334033699125706, 3.75325428681369e-05, 8.97021254811675e-08, 
    4.40053612699152e-07, 4.78226502443588e-07, 1.74025876602636e-07, 
    4.81151406255747e-07, 6.72915909545171e-07, 3.53204258352453e-06, 
    1.15492930015573e-05, 3.25525722913112e-05,
  7.41686069397842e-05, 4.14011840428105e-05, 1.43290545664993e-05, 
    5.41171879362845e-05, 0.000523210393335701, 0.000469077636057649, 
    4.05370956028074e-06, 6.04742465047376e-07, 5.2127595122642e-07, 
    1.49371018083473e-08, 2.6236449665936e-11, 4.38258214757509e-07, 
    1.14762969506629e-07, 7.36919925808582e-10, 9.22217565093801e-14, 
    3.65939146132167e-07, 6.04729144638801e-09, 0, 1.40449496420654e-12, 
    0.00032758074210512, 0.000596405287814319, 0.000384656778965471, 
    1.7426596153277e-05, 4.25486736949989e-07, 5.84895713270236e-09, 
    6.89355601394931e-09, 8.77424508451557e-08, 1.68087864381738e-07, 
    3.64351193976562e-06, 2.31570717255002e-06, 3.24967508167343e-06, 
    4.14255922299255e-06, 4.81193041857195e-06, 1.15505080798264e-05, 
    9.42866377718381e-06, 7.16869061297513e-06, 1.00771702017134e-05, 
    2.85755185625688e-05, 7.1177285423021e-06, 7.87595476200252e-06, 
    1.3653530567602e-07, 2.12160099343463e-08, 1.20008151394263e-12, 
    8.65913179423231e-07, 9.48409297534931e-07, 1.53104995259354e-07, 
    1.07979243807349e-10, 1.05460543321556e-08, 0.000104496194459424, 
    0.000148754996551015, 7.26431593614288e-05, 2.71145180100539e-05, 
    1.43659459181114e-05, 6.38518978147582e-06, 4.1520664589931e-06, 
    4.180687470497e-06, 4.21389596197353e-06, 4.33737185647093e-06, 
    3.62118144385526e-06, 2.55095574734203e-06, 2.08708874696157e-06, 
    5.16040216612254e-09, 3.04600163404075e-10, 2.1744244405906e-07, 
    5.05485369212762e-05, 0.000163688831479452, 0.000187153719072851, 
    3.40321798081064e-05, 1.09343179667082e-09, 9.48316635785223e-11, 0, 
    5.8055923302892e-08, 3.30877347734748e-06, 5.36493680482851e-06, 
    3.12841202622065e-06, 3.87657260120362e-06, 6.23285034183362e-06, 
    1.31794065571503e-07, 2.03815940024752e-06, 1.70242404872707e-05, 
    9.5369690559573e-06, 3.1441289395095e-05, 2.22911687233249e-05, 
    2.160184301052e-06, 1.2867252730291e-08, 1.01940950704677e-09, 
    4.5668658757718e-12, 2.42567682078437e-08, 2.15226582471637e-05, 
    4.54126505734033e-05, 9.73830444251214e-06, 3.57519193824274e-06, 
    2.05488789251221e-05, 0.000327712986447208, 0.000115614459558799, 
    1.41040986072328e-06, 9.32326964231564e-06, 6.24249927616827e-06, 
    1.58539877897097e-05, 5.82923091117515e-05, 0.000140848098265799, 
    3.28552676449908e-05, 2.06079834366425e-05, 7.78493389405279e-06, 
    3.21297744563792e-06, 2.55296792744568e-06, 1.22734959398648e-06, 
    1.70616225048544e-06, 6.27919888458814e-06, 6.85992610758504e-06, 
    6.74470394701882e-06, 2.32842630765315e-05, 2.02144676090413e-05, 
    1.87709304501526e-05, 0, 0, 0, 9.17668358951855e-07, 
    5.73588424993847e-07, 9.26179214096516e-07, 4.86796258500714e-07, 
    3.39078073632244e-07, 8.08437245924448e-05, 8.86438480286058e-05, 
    7.9697941377746e-05, 8.3609372418384e-05, 0.000112013041315036, 
    4.66707580806638e-05, 9.16949584850243e-09, 1.17392629559148e-09, 
    5.76040506356702e-05, 0.000289200397729989, 0.000300656914583468, 
    6.42537929207243e-05, 3.26791066443038e-06, 1.98201804824372e-07, 
    1.12895173611193e-06, 8.53179018194817e-07, 1.56802749247093e-06, 
    4.98628190378729e-07, 9.09719591369501e-07, 3.6497200673518e-06, 
    1.12487300636654e-05, 3.11784823345497e-05,
  8.78681018027317e-05, 5.31597861659724e-05, 4.6637831399928e-05, 
    5.88362570248365e-05, 0.000670271259023456, 0.000585162692343292, 
    2.1184808884595e-05, 7.79755869437058e-07, 8.33242703443012e-07, 
    8.94272629331828e-07, 1.70447278220105e-08, 1.13920524243833e-08, 
    7.92454878912894e-10, 2.91044312886594e-09, 4.08384544602981e-07, 0, 
    2.60519420906231e-13, 9.2618884284178e-11, 0.000375738291444582, 
    0.000616634536403905, 0.000318357936757126, 1.772486442079e-06, 
    2.897488998589e-08, 3.19208974174341e-09, 2.5776685264924e-08, 
    2.5693441975819e-08, 6.75055948674429e-09, 4.97179178069589e-06, 
    8.63130968905983e-06, 1.23873735971025e-05, 8.87690766690422e-06, 
    1.04453086272453e-05, 4.43621791504184e-06, 1.64782062449271e-05, 
    1.44096660913274e-05, 6.80007514390954e-06, 1.62741104566568e-05, 
    1.30255497462995e-05, 1.62740222300412e-05, 7.66426423034588e-07, 
    2.99083272217355e-08, 6.90299571218184e-08, 4.2688102328736e-07, 
    8.33037068041988e-05, 1.27706593659004e-06, 9.94553701761129e-09, 
    1.52904508751774e-09, 7.61660763563585e-05, 0.000150491617473485, 
    9.62057659376693e-05, 1.73495600082164e-05, 1.94719738552138e-05, 
    8.59835684272731e-06, 9.58358691405778e-06, 3.27895999094106e-06, 
    1.09967871365361e-06, 3.35233384376065e-06, 2.68827798462139e-06, 
    2.1295614671141e-10, 3.47944512364442e-06, 2.49883450268597e-06, 
    7.66740115406709e-07, 3.5767081267396e-05, 0.000152180865061176, 
    0.000196220518016791, 8.91281168578589e-05, 5.93918711397672e-05, 
    1.61180573992173e-05, 1.33459996141215e-05, 8.96772572094686e-09, 
    5.87614562916009e-11, 4.04681509051496e-06, 1.06717088492256e-05, 
    7.80420274373359e-06, 8.11088118866218e-06, 5.23094445455081e-06, 
    2.97285739854222e-07, 1.78731570024298e-06, 2.63222527495773e-06, 
    2.36079996646003e-06, 2.33981701333752e-06, 1.41699326263625e-05, 
    2.04989608592719e-05, 2.30789828327126e-05, 3.76994160566341e-05, 
    5.56980518644937e-05, 3.49670820515351e-05, 3.73544007457726e-05, 
    3.44637587070181e-05, 4.5564532456836e-05, 6.05992136965876e-06, 
    3.59433185588688e-06, 1.39778907732946e-05, 0.000345098528307462, 
    0.000227838226589509, 2.97743233397835e-08, 2.83271315654095e-06, 
    8.39297468594091e-07, 8.1526819719375e-06, 5.30806939755724e-05, 
    0.000237737763946124, 0.000176911853442758, 4.09024580902429e-06, 
    1.05663477990809e-05, 4.36161029751247e-06, 5.15604697673661e-06, 
    1.70954093118608e-06, 4.8326619777038e-06, 6.64142099162454e-06, 
    7.11530096950002e-06, 1.20778384931973e-05, 1.21531792581696e-05, 
    2.02434148543218e-05, 2.50544540014294e-05, 5.73036330790522e-06, 0, 0, 
    0, 1.35595926063523e-06, 4.56370982510247e-05, 1.7014249594542e-05, 
    1.46171257927135e-05, 5.67721341263304e-05, 6.06394947989746e-05, 
    9.44357057975978e-05, 6.16825185563152e-05, 1.76064469162504e-06, 0, 
    2.06297302492615e-07, 9.89145114664574e-05, 0.000436035255946275, 
    0.000334486145331308, 3.59855907405768e-05, 6.94852900758756e-06, 
    9.78722038364201e-07, 1.88352023501505e-08, 6.2322362957505e-07, 
    1.23865753840829e-06, 7.32911150083086e-07, 3.68590935912371e-07, 
    6.60779248309047e-06, 2.26018398290432e-05, 4.45217276277542e-05, 
    6.17570258365871e-05,
  4.06959867803237e-05, 1.46533473558277e-05, 7.0079236565348e-05, 
    0.000226895061601964, 0.000565351199379927, 0.000283790836331806, 
    9.03090412150791e-06, 3.63335163038373e-07, 3.1288182946797e-07, 
    6.38569594902626e-09, 1.9842579866383e-11, 4.01430547853371e-13, 
    1.05678511174277e-11, 1.79423021355399e-13, 2.15310716983403e-05, 
    4.38118736702423e-10, 1.02047358481021e-06, 0.000365788210708065, 
    0.000602111108867916, 0.000277837399075249, 9.53493190826339e-08, 
    4.36400696099519e-09, 4.879529200376e-09, 3.58384045293296e-08, 
    9.22944244513051e-06, 1.0193905941425e-07, 6.90451965302482e-06, 
    6.67280280407774e-06, 5.11649118301415e-06, 7.40538226218485e-06, 
    6.87034194536589e-06, 1.185664531266e-05, 1.03650715165419e-05, 
    1.20899800822046e-05, 1.73169994744473e-05, 6.19590245331035e-06, 
    1.19032038163755e-05, 1.68820507661432e-05, 2.49635247564625e-05, 
    2.51429667476544e-05, 2.03777667852048e-05, 7.50164827850468e-05, 
    0.00013191149085863, 7.76207905327567e-05, 3.42859217780087e-07, 
    4.69452456943387e-08, 7.17089747428878e-05, 0.000153217936826297, 
    0.000131053823606189, 5.32857975335282e-05, 1.74318585024146e-05, 
    1.46795925009442e-05, 9.98852939422847e-06, 1.30076015811211e-05, 
    6.9490110694965e-06, 4.80494323657686e-06, 2.31586823212344e-06, 
    1.56818907179969e-06, 3.88798459794778e-23, 9.15607087330044e-06, 
    7.90244873618252e-06, 0.000212264214551409, 0.000166867414519186, 
    5.7597765214734e-05, 2.84117346149623e-05, 1.44833309907241e-07, 
    1.44447787647025e-05, 1.15449652435071e-05, 2.98502497403269e-05, 
    1.37271971880804e-05, 7.12872893324229e-09, 1.29909152624339e-23, 
    4.41087614904683e-06, 3.60577075305791e-06, 7.25912569463736e-07, 
    2.65975089911112e-06, 3.8654083489342e-06, 2.10892227858953e-06, 
    5.34471755350611e-06, 3.72198324294292e-06, 5.24088984110611e-06, 
    9.95868858893103e-06, 1.87003506513587e-05, 3.83370163977829e-05, 
    4.40975671405318e-05, 4.93392412046766e-05, 4.07188407328491e-05, 
    4.10803044181923e-05, 3.110694245565e-05, 3.70690533394373e-05, 
    2.28726629786368e-05, 3.65639868261883e-06, 1.79573925640252e-05, 
    0.000355053151141614, 0.000338159804646995, 4.7247332660262e-08, 
    7.96131209164522e-07, 3.47039487839247e-08, 2.41046827326501e-06, 
    1.93119014395607e-05, 0.000211108046477024, 0.000293702234820837, 
    2.82689263301067e-06, 1.08555863895245e-05, 6.56362841495415e-06, 
    5.36252923315399e-06, 4.37716249788056e-06, 4.29613063232143e-06, 
    5.25552878138989e-06, 6.52050173921233e-06, 8.66359064855804e-06, 
    1.0808908229686e-05, 2.2571860831437e-05, 3.39503975740793e-05, 
    5.35463322545835e-06, 0, 0, 0, 8.0813562508642e-07, 0.000118776413617933, 
    4.26680265685092e-05, 2.47417759276991e-05, 4.37546815182261e-05, 
    0.00014854703690464, 7.9330325928382e-05, 2.04751593854193e-09, 
    3.36998206703994e-09, 3.56514173432769e-07, 0.000139068854752497, 
    0.000728165233198789, 0.000506369504153289, 5.12779124958212e-05, 
    1.00907253801326e-05, 7.66225915840929e-06, 9.3826547417899e-07, 
    2.71626756253329e-07, 1.35834283235736e-07, 1.56284809016943e-06, 
    2.18036597515116e-06, 3.85736679110696e-06, 5.19235477190438e-06, 
    1.23771659001896e-05, 2.17838447350881e-05, 5.47450000260703e-05,
  3.3792093381008e-06, 2.16511457408006e-05, 0.000150036636642686, 
    0.000274657606886673, 0.000151069143290934, 9.08897918686335e-06, 
    5.46432767906745e-06, 4.36781147240459e-06, 2.15477923085222e-06, 
    4.4700610902874e-06, 9.79233489759282e-06, 1.59551829031999e-05, 
    4.59073920923162e-05, 4.61754891556357e-05, 2.48582886239507e-05, 
    2.94239903258045e-07, 0.000222030766371139, 0.000489542907156765, 
    0.000408310892994111, 5.29245431624056e-05, 3.16623715144904e-09, 
    3.66859862549213e-06, 4.94122245724157e-06, 5.95636075530337e-06, 
    9.34142625099246e-06, 1.30468672763097e-06, 5.61823297828383e-06, 
    4.76530982887886e-06, 3.29313018434933e-06, 3.60687276148512e-06, 
    1.72064535481801e-06, 4.27927963303471e-06, 1.41566956922809e-05, 
    9.50832471997987e-06, 1.24079090136068e-05, 1.77729703221207e-05, 
    1.64232026591988e-05, 1.93912612367643e-05, 2.76895589104049e-05, 
    2.35833711187324e-05, 5.15451423508368e-05, 6.62776080442488e-05, 
    4.95585204706172e-05, 1.30223661376998e-05, 2.09882309711622e-05, 
    5.85023061710057e-05, 0.000134081090722189, 0.000100898412520687, 
    4.23261936545913e-05, 3.65244071343484e-05, 4.1636676096391e-05, 
    2.23020505603368e-05, 2.44199597930922e-05, 1.31361885901906e-05, 
    1.0459894104724e-05, 4.50259430626862e-06, 2.78040195922263e-06, 
    1.22493112882296e-06, 2.89223239103647e-06, 5.59898093928233e-05, 
    0.000280368338196602, 0.000308406532178446, 1.06284457925079e-05, 
    4.15653799205924e-06, 3.2505440634132e-19, 1.22305202838796e-06, 
    5.92719889741976e-06, 2.6481042115604e-06, 1.22449670914928e-05, 
    2.2382458717849e-05, 8.43632141442767e-06, 6.92250751269619e-06, 
    3.71801696138161e-06, 2.80031924428249e-06, 1.38832302020396e-06, 
    2.61117105080304e-06, 2.81737322235322e-06, 2.70826136199217e-06, 
    2.32134625778893e-06, 5.05076683465504e-06, 9.53355020427553e-06, 
    1.32737803375266e-05, 2.13452667844347e-05, 4.14233269550225e-05, 
    6.82403193683368e-05, 4.32246763330691e-05, 4.27920411180265e-05, 
    7.9480931236628e-05, 5.44582614164454e-05, 2.86404712822033e-05, 
    7.62442704874368e-06, 1.58447094771297e-06, 1.18920878510487e-05, 
    0.000305302992024585, 0.000372411580428192, 8.54608443852702e-10, 
    3.75220673931209e-07, 2.2493681453978e-06, 4.16847219688898e-09, 
    4.02416042686722e-06, 5.08182289628739e-05, 0.000485977204714, 
    0.000119063077360108, 3.5311526077004e-06, 7.17272154440781e-06, 
    4.96412046069591e-06, 5.5699499504406e-06, 3.99891009536565e-06, 
    4.06131385697368e-06, 6.3101367792744e-06, 9.72177774053791e-06, 
    1.37083239241581e-05, 1.68232650648026e-05, 2.00997798895357e-05, 
    2.34459285842377e-07, 0, 0, 0, 1.41895868379889e-08, 
    9.49580779889508e-06, 1.52164085916498e-05, 1.4054385634782e-05, 
    2.39041887812322e-05, 2.40043458293462e-05, 2.24101562981833e-08, 
    9.36409184635739e-08, 4.85809195338223e-08, 0.000199078029353121, 
    0.00083630898602907, 0.000700923215076046, 0.000143615254374126, 
    1.87026631031677e-05, 1.28809110003848e-05, 9.37008033859826e-06, 
    1.79972191300702e-06, 1.00142987553871e-09, 1.40756771630427e-11, 
    8.02586600134925e-10, 8.38977788835099e-09, 1.23350189885245e-08, 
    2.76184849063306e-08, 1.29785485119846e-07, 5.92375944192066e-06, 
    1.44520144359083e-05,
  3.46248322346875e-09, 9.14796215752025e-05, 0.00012417830751615, 
    7.44342015507594e-05, 6.17557498507574e-06, 1.50523770928525e-06, 
    2.54668662074588e-06, 2.46485201230146e-06, 4.14942571920292e-06, 
    1.68176343835773e-05, 2.07541711653279e-05, 2.64989621201696e-05, 
    6.32543004975128e-05, 5.25954715417002e-05, 1.16686068918118e-05, 
    7.57623632763946e-05, 0.000328326417204979, 0.000237031880045493, 
    9.7145482569495e-05, 2.56777208971261e-05, 7.81871276450631e-06, 
    1.11030992484167e-05, 8.21414375226967e-06, 3.60244081213613e-06, 
    2.0461344855908e-06, 5.70799118808622e-06, 5.10523035366271e-06, 
    2.98417179714083e-06, 6.47838190573986e-06, 2.55444547102671e-06, 
    3.06473040261041e-06, 1.2295150640476e-05, 9.34381271536799e-06, 
    1.36216256800382e-05, 8.76504585648718e-06, 1.48019998562585e-05, 
    2.29133444170459e-05, 2.42275650674687e-05, 2.59315101951801e-05, 
    3.5002967741984e-05, 4.79259235852291e-05, 2.77664249294371e-05, 
    9.30095633639272e-06, 1.74566238599779e-05, 7.21160678745258e-05, 
    0.000120663904146855, 0.000108273176138875, 7.70061125890745e-05, 
    4.7958327360298e-05, 3.92167321863442e-05, 3.52796615146405e-05, 
    1.16036396627212e-05, 6.00978246693145e-06, 3.46842382564412e-05, 
    1.42769672036978e-05, 8.29337767787855e-06, 6.40952268456598e-20, 
    1.11488772928215e-20, 1.11368489604115e-10, 0.000117181724891402, 
    0.000200993961009333, 0.000117478818018998, 0.000154248265085605, 
    4.3639915142214e-05, 2.77816960344154e-06, 5.86662991008111e-06, 
    6.76967807093063e-06, 9.50331730591463e-06, 1.18668462268634e-05, 
    8.96964391571348e-06, 4.55594596424105e-06, 1.36727623689818e-05, 
    6.07727524943098e-06, 6.4383756535129e-06, 7.78290775306532e-06, 
    3.07298883399694e-06, 9.765067831574e-07, 2.68304647275282e-06, 
    2.97466323218384e-06, 5.13360099417979e-06, 8.75009269622774e-06, 
    7.44220566762921e-06, 2.28998542139922e-05, 4.34786230562972e-05, 
    5.5998960522503e-05, 4.79968951146774e-05, 3.56225072876575e-05, 
    7.6050519378493e-05, 6.96182083669096e-05, 4.02347395923705e-05, 
    1.41523122401356e-05, 5.74898817905182e-07, 0.000104726525506368, 
    0.000305440204057858, 0.000345110707647423, 3.58946278632052e-07, 
    1.96721049054141e-06, 2.2397069657032e-09, 3.34994625014353e-20, 
    6.07695600252867e-12, 1.26907638204446e-05, 0.000274321459155385, 
    0.000497119159012857, 0.000183914919963001, 1.32729622512601e-06, 
    2.36386642135986e-06, 5.84881480588002e-06, 6.56107318387878e-06, 
    3.66814067991288e-06, 3.81797223740037e-06, 6.3518527845402e-06, 
    7.10331520442167e-06, 8.60959770735683e-06, 1.12747553511588e-06, 
    1.26555743243966e-10, 3.79907619993059e-08, 9.69184493387794e-08, 
    1.13667249802912e-08, 6.25801442183423e-09, 5.85633349670989e-09, 
    8.00466867809161e-10, 1.01610346508543e-09, 1.84307437700414e-11, 
    7.60108782825233e-10, 5.28803895258732e-08, 1.99569916047149e-05, 
    0.000365914991936169, 0.000583368003607838, 0.000525671929447766, 
    0.000198466878459849, 8.18922280062968e-06, 8.97644509060546e-06, 
    6.99746626999331e-06, 1.58553676587265e-07, 2.55320848603499e-10, 
    4.11543638410797e-10, 3.30906420832503e-11, 0, 0, 0, 
    2.35817030119581e-11, 0, 3.89818172052294e-08, 5.52480324899918e-07,
  8.75710147093307e-05, 6.2388640042594e-05, 5.38295562363192e-06, 
    2.50140719607222e-06, 1.53185500572515e-06, 4.68645252507753e-08, 
    4.25335552327293e-07, 4.27764529567091e-11, 2.2203214885812e-06, 
    1.87750537274022e-05, 5.38901768812485e-05, 0.000132961745772862, 
    0.000109116912779554, 3.13870356108596e-05, 3.81673838186978e-05, 
    0.000370907383750114, 0.000202110228755206, 0.000105585562608006, 
    5.5435959485227e-05, 2.88392423462385e-05, 2.80693488119131e-05, 
    1.27747023077187e-05, 8.5597422855868e-06, 1.77617526111118e-06, 
    1.05676991558343e-11, 1.15930821723033e-06, 1.08545591903989e-05, 
    1.37584361288238e-05, 8.42457815927018e-06, 6.95008046960981e-06, 
    6.08170299593708e-06, 1.05869089905953e-05, 9.7417934648851e-06, 
    1.44364870824802e-05, 1.06404751359948e-05, 1.77482723115587e-05, 
    1.9387924310598e-05, 2.24902022891212e-05, 1.69053438573053e-05, 
    1.19881005914473e-05, 9.85124847948022e-06, 8.3832246577617e-06, 
    1.0828739010877e-05, 4.77690380447304e-05, 7.033077663102e-05, 
    7.03474023030103e-05, 7.57131028713274e-05, 4.0198541419863e-05, 
    1.90697784364852e-05, 2.17912596091788e-05, 3.02753439485645e-05, 
    5.8454544151011e-05, 4.45847863841257e-05, 3.81816885492343e-05, 
    8.70082592786422e-06, 4.9693129788928e-09, 3.07815479665444e-18, 
    3.01176251328833e-20, 4.54285895181215e-16, 1.50501902406639e-05, 
    5.20189790318895e-06, 0.000230536175502618, 0.000297476293316662, 
    0.000158257207193071, 7.05388430471908e-05, 1.11632667296234e-05, 
    9.71404956001609e-06, 1.92891956005774e-05, 1.47245622583696e-05, 
    1.21038957343679e-05, 1.43078854176661e-08, 7.66818185194143e-06, 
    3.96765134139777e-09, 1.04739475391276e-05, 1.06184823721041e-05, 
    8.81010514918057e-06, 1.36409091620053e-06, 2.3321257591626e-06, 
    3.11806698882118e-06, 2.54803291076961e-06, 4.38789557438083e-06, 
    5.12989545097202e-06, 4.9529947306662e-06, 1.64060463111552e-05, 
    2.47492309544575e-05, 6.49807214192895e-05, 5.4076389509288e-05, 
    3.17492872007249e-05, 3.30138184997735e-05, 1.7810875313018e-05, 
    2.08858144972094e-05, 1.72269531362694e-06, 0.000153058745281886, 
    0.000292242023693225, 0.000279975000581565, 5.67722076354614e-11, 
    3.88306509389414e-07, 6.18937237748448e-07, 7.69080169158278e-10, 0, 
    1.01096115631675e-12, 4.82660091312441e-05, 0.00045121144188894, 
    0.000625646300513235, 0.000172010946961419, 1.1820582390232e-06, 
    3.53715496591217e-06, 1.62200855198375e-06, 1.80290660549451e-06, 
    4.10733556160189e-06, 4.62321710222038e-06, 4.25716070902391e-06, 
    7.43681700533556e-06, 3.16162869144493e-06, 7.35409579802043e-06, 
    1.76469310250602e-07, 7.14479474052943e-09, 1.975116305704e-07, 
    1.57219531620891e-06, 2.8993004873703e-11, 3.85986234081069e-14, 0, 
    8.20609074945075e-10, 0, 0.000221022521841611, 0.00031272502801145, 
    0.000245116026686202, 0.000151725004791689, 4.23070804791171e-05, 
    2.7980224282789e-08, 1.66072908144727e-06, 2.53989139453864e-07, 
    4.97410245179515e-09, 1.86919681054527e-08, 7.38445103126579e-09, 
    4.81068112836044e-09, 0, 0, 0, 0, 0, 0, 1.13743075116884e-06, 
    9.76219907020607e-06,
  1.98855045508515e-05, 1.77862700618442e-06, 2.52645202172668e-06, 
    2.55288699117756e-07, 3.93785758455555e-07, 6.95053600666923e-07, 
    1.93268554543798e-08, 0, 0, 1.19864867689485e-10, 3.67283216974899e-05, 
    0.000106550931833563, 8.00351152581455e-05, 7.58908981124645e-05, 
    0.000148145186340136, 0.000280237133946329, 0.000190201690464006, 
    0.000121440172039996, 2.47741114804991e-05, 1.50014718801754e-05, 
    7.66116719846693e-06, 5.57204959081756e-06, 4.70536905450688e-06, 
    1.75035836844935e-06, 4.77982486322653e-09, 8.21813254425509e-06, 
    1.32834269390092e-05, 2.60087300338487e-05, 2.11038371245267e-05, 
    1.34536851075377e-05, 8.99788351877585e-06, 9.6352356933615e-06, 
    1.41116466580586e-05, 1.20103784298187e-05, 1.88694307209634e-05, 
    1.53193919312778e-05, 1.3487004277054e-05, 9.45466007073957e-06, 
    7.70881533652687e-06, 8.60045905870846e-06, 7.04709935646192e-06, 
    1.43874168737593e-05, 5.43027917592766e-05, 9.78368044342525e-05, 
    6.5595134654773e-05, 6.91780935998045e-05, 5.96776353299838e-05, 
    4.26791884939839e-11, 6.41747533918991e-09, 1.07735171888535e-12, 
    2.61499795201091e-17, 3.99049917361388e-06, 1.35509548255122e-09, 
    2.42789652097699e-05, 2.06770377060531e-24, 2.07025764291831e-13, 
    2.24174676138023e-10, 1.55079901043392e-21, 5.4365915291416e-21, 
    4.25815747066239e-08, 0.000178020938895918, 0.000269382153752124, 
    0.000361976067646448, 0.000402583287397459, 0.000171050434422788, 
    2.54472631961648e-05, 1.30392298467567e-05, 1.13795352190119e-05, 
    3.01083491293071e-06, 1.11386290659408e-05, 6.53537723377392e-06, 
    1.09276145776339e-05, 1.35652930859982e-05, 2.30218133843474e-05, 
    1.86997877839172e-05, 1.84941525929114e-05, 1.38537595856291e-05, 
    2.16489976504704e-06, 2.44206768291803e-06, 2.47720186728668e-06, 
    2.31808746509207e-06, 9.18160227182935e-07, 2.63846533928284e-06, 
    1.01624161575378e-05, 3.38935987860449e-05, 3.83634598917708e-05, 
    2.59558999973082e-05, 2.6167892527596e-05, 3.35388679897964e-05, 
    2.00588763543575e-05, 2.00023056152857e-05, 6.14171353868504e-08, 
    0.000201014091473518, 0.000378382870381527, 0.000191707573627018, 
    1.90461227200974e-07, 8.40379407228027e-08, 1.37378658553819e-06, 
    1.60108978560868e-06, 1.65819287791171e-08, 1.30893043240603e-05, 
    2.46522261595002e-05, 0.000252797239574354, 0.000688298887607072, 
    0.000504413989538109, 3.89012107238319e-06, 1.23119930142476e-06, 
    2.03324966135788e-06, 1.95272035571524e-06, 4.46600372704163e-06, 
    2.83607610918533e-06, 2.31544294639336e-06, 2.18187540496248e-06, 
    6.01983337724141e-06, 2.88595661710429e-05, 1.94865657267275e-07, 
    4.19964651191471e-07, 2.30454400388954e-09, 3.35569457576983e-13, 0, 0, 
    5.88546374452334e-24, 8.50446145183591e-05, 0.000391088509591594, 
    0.000276992919483926, 1.1021301794724e-05, 3.7394219449073e-09, 
    1.23618192209693e-10, 3.39764923080455e-10, 2.80644483906292e-11, 
    2.99326496515039e-09, 1.11320529013836e-09, 1.2613492027135e-11, 
    6.87979589101667e-22, 2.59194162717559e-11, 2.52336158002935e-05, 
    1.76139531768433e-06, 8.75515395109444e-06, 6.4154554025949e-19, 
    7.09812918929081e-12, 7.83415922087954e-18, 6.32099731078657e-17, 
    1.64834418838713e-05, 3.63844999326448e-05,
  3.39457412435205e-07, 1.76114399769082e-09, 6.3698238496978e-18, 
    1.40519104790231e-08, 1.22967533636429e-06, 1.13641876384791e-06, 0, 
    2.90745054791178e-11, 5.54447828506394e-11, 0, 1.07408590034815e-09, 
    3.09615904393653e-05, 4.68550828470202e-05, 0.000132254839655579, 
    0.000168000025611731, 0.000233962637371717, 6.23659350257629e-05, 
    3.21380529348827e-05, 2.05151788706888e-05, 3.52027404803707e-06, 
    5.8800235496265e-06, 4.05933252575503e-06, 3.03276504151433e-06, 
    2.04915002801982e-06, 2.64554976106092e-06, 7.24430397682402e-06, 
    1.52124625968983e-05, 2.36114765359681e-05, 2.19001451523838e-05, 
    2.47433800293307e-05, 3.07895110434611e-05, 1.32113953200524e-05, 
    1.42485956076191e-05, 1.30979750382056e-05, 1.15306461729331e-05, 
    1.07653891775591e-05, 1.06275128957502e-05, 8.79619918665187e-06, 
    6.34048783648934e-06, 5.34789973317024e-06, 2.07720130860984e-05, 
    8.42006308298468e-05, 5.59128273501489e-05, 4.34897934755418e-05, 
    2.94275721922256e-05, 5.38596246839478e-05, 6.11846107418667e-05, 
    8.62233061011097e-14, 1.50752467919043e-20, 2.18515638506922e-19, 
    1.51138720425852e-12, 1.20647248277485e-18, 0, 0, 4.13941459021236e-17, 
    2.45103246889397e-11, 1.15097270043585e-10, 5.86868781969004e-15, 
    6.0776804862964e-09, 5.06004004899343e-07, 6.3667930377295e-07, 
    2.24197044175778e-06, 0.000432776941956483, 0.000500958868669915, 
    0.000276758522367342, 9.81185903079476e-05, 1.01373830896867e-05, 
    3.82765141122988e-06, 1.13836563633084e-05, 1.25408946281426e-05, 
    1.53249479146326e-05, 1.73948823810654e-05, 1.03706795417403e-05, 
    4.50934138852248e-06, 6.88084643118557e-06, 3.386157770914e-09, 
    3.53026817214363e-06, 8.84138290523346e-06, 4.66400833025466e-06, 
    2.06138170395988e-06, 1.85711051140189e-06, 4.84881996705888e-07, 
    1.46783045629821e-07, 9.78945424490664e-06, 1.57170091061905e-05, 
    1.5684161188111e-05, 1.3920495496091e-05, 2.81407762726588e-05, 
    1.38545847718992e-08, 1.20488408818049e-09, 2.92528153955946e-10, 
    4.76220211266645e-05, 0.000245818207833103, 0.000327579919274162, 
    1.44926880065669e-05, 3.99660596231334e-07, 1.55400435344526e-10, 
    9.74762735383355e-10, 1.79630304543858e-09, 5.14913014723045e-12, 
    1.58864527898414e-05, 1.41570349629822e-05, 0.000105577492863132, 
    0.000595875178992867, 0.000548656270187994, 0.00013089732908463, 
    1.53180040419787e-06, 1.53251419543066e-06, 1.06709691026545e-06, 
    2.95698876799939e-06, 2.15227701963736e-06, 2.22137582799644e-06, 
    2.174638505219e-06, 2.15815846309241e-06, 3.71345215318061e-06, 
    7.32499142391086e-06, 1.35560522313581e-07, 2.36602729057264e-10, 
    1.16320959702235e-10, 7.7354261859113e-26, 2.6913474144209e-10, 
    2.93070830819704e-05, 0.000244592362946151, 4.3212446819254e-05, 
    3.14094756741119e-07, 1.89788660684381e-11, 1.12354960153081e-20, 
    1.67010917806179e-10, 5.785871151505e-11, 5.44251611013035e-09, 
    5.35874187506144e-08, 2.37990703830278e-09, 0, 2.76783337652701e-08, 
    3.96268111837073e-20, 8.73892672741166e-06, 3.91077548455915e-06, 
    7.12028689385028e-06, 9.44576795242392e-06, 9.42135066086965e-06, 
    1.21805388454514e-05, 1.53573958662011e-05, 1.68803274243439e-05, 
    1.85934536760725e-06,
  2.0219262113937e-09, 5.58303733672226e-07, 4.28224759844069e-07, 
    1.56275662725713e-07, 1.10124865868583e-06, 1.26518172983378e-11, 0, 0, 
    1.00020407294337e-09, 1.01675911665675e-08, 9.74763381985949e-12, 0, 
    1.95065028553581e-05, 0.000234656052592388, 0.0001632462427889, 
    8.8220183397606e-05, 2.31931243161197e-05, 2.53022900121385e-05, 
    4.18629102188843e-05, 3.73346652861009e-05, 4.37938568992273e-06, 
    4.60113174761568e-06, 1.76222152282192e-06, 8.47947452688774e-07, 
    3.91421131746136e-06, 3.82586959189084e-06, 1.03145445514954e-05, 
    2.40747221661307e-05, 2.32689252718005e-05, 2.77926791165147e-05, 
    2.30841264257201e-05, 2.45869330472961e-05, 2.51370701969593e-05, 
    1.48291623364468e-05, 1.37082024893045e-05, 1.38098503781485e-05, 
    1.27452112730148e-05, 8.91871482560642e-06, 1.5222716467771e-05, 
    2.38436508574973e-05, 6.99426609957151e-05, 8.32651263409235e-05, 
    5.67432750885434e-05, 3.19230454783665e-05, 1.20605830861051e-05, 
    6.57767165788364e-05, 1.43571453855066e-06, 2.37486885717879e-09, 0, 
    5.43998983612678e-12, 1.2470573716925e-10, 7.15980363533371e-12, 
    1.02136747206013e-09, 7.92349057544336e-11, 9.65337872915142e-12, 0, 0, 
    0, 2.32948881665645e-18, 7.01482025483475e-05, 3.8896806767903e-06, 
    0.000105281826188319, 0.000106379463871861, 0.000203818031879214, 
    0.000180569198880046, 7.89715006961596e-05, 1.61012354787013e-05, 
    4.91288335721815e-06, 6.97846602563433e-06, 1.21500541159246e-05, 
    1.8108509099423e-05, 2.21071298630711e-05, 2.4068171716989e-05, 
    2.89795977937418e-05, 2.59410414238556e-05, 2.49214805951626e-05, 
    1.74221271103779e-05, 9.3398363739518e-06, 5.70498688215869e-06, 
    3.55404217537245e-06, 1.19675324566915e-06, 2.49262876828682e-06, 
    1.90618721503288e-06, 2.10323318304449e-06, 3.4713606441457e-06, 
    2.37051272958996e-06, 1.37476510665269e-07, 2.56199116089072e-11, 
    3.26645320092027e-11, 1.46198420657532e-10, 2.30916026548516e-06, 
    0.0001180314571661, 0.000166194933575435, 7.69332895741661e-05, 
    1.96045011320649e-06, 1.3609601996757e-08, 7.57616880087065e-10, 
    2.8717422699703e-07, 8.78456658858817e-07, 0, 4.96597481040262e-06, 
    3.51823307831828e-05, 0.000130334053925119, 0.00047565450487996, 
    0.000299453730781193, 7.25270000904592e-05, 3.60494216773533e-06, 
    3.4630631425226e-06, 1.82512377485932e-06, 1.62572754865439e-06, 
    2.45532420250198e-06, 5.03941096297664e-10, 6.33331486714462e-07, 
    5.16029349115125e-10, 4.54567871351045e-09, 2.76507001603994e-09, 0, 
    5.17286409394172e-07, 2.7907452148017e-11, 1.18765559582968e-22, 
    1.96861985893357e-11, 2.93351709737801e-08, 3.94188799594854e-07, 
    2.5563640917127e-11, 0, 0, 3.29677642617444e-22, 1.02442360720528e-09, 
    3.13423618716219e-09, 3.01956239500555e-08, 2.7546677453633e-06, 
    4.22379092541533e-09, 1.51009020011691e-11, 5.85198395783597e-07, 
    3.88280229773352e-06, 7.16885145477878e-06, 4.39369040880312e-06, 
    4.96776713064442e-06, 2.36686993024879e-06, 4.41840380681932e-06, 
    3.48688876136273e-06, 1.86959444339285e-06, 7.44047508349566e-10, 
    2.42640741158839e-10,
  2.16311316979969e-06, 7.14538364786984e-07, 1.00472233040765e-06, 
    3.22430440256043e-07, 1.75540524707583e-08, 0, 0, 0, 0, 
    1.62868016119284e-10, 1.69921761850462e-08, 1.03976982512229e-09, 
    9.33790886411086e-11, 1.47577899101105e-11, 8.40620367984616e-05, 
    3.11687324878763e-05, 1.79265489346216e-05, 4.82751383955226e-05, 
    4.22623643649911e-05, 2.92144791404169e-05, 1.60288944657845e-05, 
    3.03904522712744e-06, 1.81311694233131e-06, 2.50447721717008e-06, 
    7.78032938060195e-07, 4.78287342503477e-06, 1.01061728353127e-05, 
    3.37589346060564e-08, 5.39490766665113e-06, 9.41683111278773e-06, 
    1.55668644172205e-05, 2.12861198772982e-05, 1.8558259730567e-05, 
    1.76888345507791e-05, 1.72705444241685e-05, 2.06938443751556e-05, 
    7.51504170110258e-06, 2.79196157040967e-05, 4.0340081899408e-05, 
    4.97327976057681e-05, 4.10939322522647e-05, 2.93245733633568e-06, 
    9.18681820198225e-06, 2.10364185144056e-05, 2.47930161804096e-05, 
    3.67930963691047e-05, 0, 3.09926617833947e-16, 2.52337900862722e-11, 
    4.54140152421049e-12, 9.64133919876734e-19, 4.45346011113785e-12, 0, 0, 
    0, 0, 0, 7.769166813716e-07, 2.91118317753722e-09, 0.000146714747924882, 
    5.72032042822051e-05, 6.46838081717435e-05, 9.56376228630153e-05, 
    0.000209492115412263, 9.86817892352843e-05, 8.32492352983392e-05, 
    3.86179207975493e-05, 1.6659653252381e-05, 6.96496259652472e-06, 
    1.42943002675465e-05, 2.31192369608613e-05, 2.26795894434295e-05, 
    1.71952290982709e-05, 1.30939115690188e-05, 1.35652558098325e-05, 
    9.19067073688619e-06, 3.22284754734644e-06, 5.12322286636679e-06, 
    7.36621065430312e-07, 7.90702802762831e-06, 1.15262796742102e-05, 
    1.26487434008622e-05, 1.29096612239616e-05, 4.24312008937825e-06, 
    2.11372382725698e-06, 1.26573545605734e-09, 1.78625762300205e-10, 
    1.03140058002833e-08, 7.33745032983743e-07, 7.7625417776009e-06, 
    8.45352590666143e-05, 0.000234515719480347, 0.000157567421275621, 
    1.50516071131511e-06, 4.83921381096798e-06, 1.48609755027008e-08, 
    4.81241299962801e-11, 6.13976044097423e-08, 5.36430383872358e-06, 
    2.7286989813652e-06, 1.45380086579955e-07, 6.57131257876873e-05, 
    0.000206826402095301, 0.000302514349839471, 0.000137476913714373, 
    6.38785915658509e-05, 1.59601579418737e-05, 1.88243569988576e-06, 
    1.29873166918085e-06, 5.46753809297841e-06, 1.35116785505978e-06, 
    8.31303656164302e-07, 3.09166795466013e-06, 4.06840695443807e-10, 
    2.74342552458638e-09, 3.03181846699472e-09, 1.32872333534437e-10, 
    3.18462678384002e-10, 1.42673200151746e-17, 0, 5.18322190823545e-24, 
    4.57929845063297e-20, 2.67577790209491e-08, 2.37193869436002e-14, 
    4.8209524682998e-18, 0, 0, 3.05252965214459e-10, 1.05915204204785e-11, 
    3.61489656024272e-06, 2.07583509539553e-06, 1.26835560658137e-06, 
    7.58383959385503e-06, 5.50618896194796e-06, 1.25472141444779e-05, 
    1.14204026062373e-05, 2.19617890080416e-07, 5.96242170879526e-06, 
    3.50811276518225e-06, 3.28091541406908e-06, 4.28341784677157e-06, 
    2.7596915387662e-06, 6.74515145178889e-07, 1.28535504505076e-06,
  6.57242176840735e-06, 9.27737700227656e-06, 6.89581255730618e-06, 
    2.39806843443521e-06, 0, 0, 0, 0, 0, 0, 0, 1.18340975811368e-18, 
    6.58649626836138e-12, 7.90607075527657e-18, 1.15714366430433e-05, 
    4.07251744095277e-07, 4.56242804488375e-06, 2.69355531712169e-05, 
    3.54386828496888e-05, 5.54941781938384e-05, 4.5212588583275e-05, 
    2.02777911470003e-05, 2.87666457477882e-05, 5.66672121105407e-06, 
    6.81606532989856e-06, 1.03976577153991e-05, 4.54820724452064e-06, 
    8.53887432954897e-06, 2.21716406081065e-05, 2.8917895036434e-05, 
    2.73815286268812e-05, 1.76086169472363e-05, 2.33020369035883e-05, 
    1.44290675871728e-05, 1.47386261232723e-05, 1.38736693788047e-05, 
    1.15237202177428e-05, 2.67945324034698e-05, 2.74894303657312e-05, 
    2.78873226456284e-05, 1.53868204108068e-06, 6.18401236865477e-06, 
    5.64745102823498e-06, 4.25752993111633e-06, 1.29382971259608e-05, 
    1.51883774180763e-10, 1.03201780661704e-24, 0, 2.36419526534499e-13, 
    7.17086396070987e-11, 8.04442840389436e-11, 3.80892760032954e-10, 
    5.85050143932564e-08, 7.93025016414408e-08, 0, 7.24634608740868e-09, 
    2.91600957420373e-09, 7.52045087135399e-08, 1.20851099927142e-08, 
    4.92335747339064e-05, 1.43918855417485e-05, 4.2305280741235e-05, 
    4.20469881446781e-05, 7.60451952527216e-05, 0.000129716840752481, 
    0.000106574658679689, 4.35772174005438e-05, 1.19374825796563e-05, 
    1.44284220393755e-05, 2.07303892551051e-05, 2.84261064928818e-05, 
    6.59772076216615e-06, 5.11315547925109e-06, 6.78051699004077e-06, 
    2.91137487805203e-05, 2.85249076751824e-05, 2.28568744668833e-05, 
    6.05967966261383e-06, 6.14410264972662e-06, 5.31372701598405e-06, 
    9.40258294281795e-07, 1.79322846275132e-07, 4.03097426079301e-08, 
    1.54415198434502e-08, 6.73991939533667e-14, 1.39908929357729e-14, 
    7.10679420097465e-06, 3.35408799898583e-05, 7.40569289962409e-05, 
    9.07977750275991e-05, 0.000118172900958879, 0.000151539331758934, 
    7.95958631412271e-05, 6.63681536770517e-07, 1.55010434430522e-05, 
    2.69226798513531e-06, 4.07411333173416e-08, 0, 1.91813910689762e-09, 
    4.07522735443177e-06, 1.24624253641952e-05, 5.41713660831358e-05, 
    0.000116401043009608, 0.000114630476239234, 5.91630732063105e-05, 
    6.69036944620318e-05, 2.79322319842444e-05, 9.93140914955135e-06, 
    1.33967790312232e-05, 8.4169593963889e-06, 5.14381831320801e-06, 
    3.56839431307095e-06, 1.61998414725036e-07, 0, 2.69310653629999e-10, 
    2.01522184697653e-08, 4.27248106845956e-11, 0, 3.23331799717409e-25, 0, 
    0, 4.2260965562052e-19, 0, 0, 0, 0, 0, 2.59263459590683e-09, 
    3.84662961930076e-06, 4.69481746763958e-06, 2.05268988109819e-06, 
    7.67924581607241e-07, 3.88924298065049e-06, 1.18839102584674e-05, 
    1.14517243064376e-05, 1.43443795247738e-05, 1.21446150994576e-05, 
    5.26566000531688e-06, 9.67496007380018e-06, 8.79449285052137e-06, 
    3.65964345438806e-06, 4.13162205901156e-06, 3.388298925251e-06, 
    5.14360938177082e-06,
  2.76146554622666e-06, 2.07265070570921e-06, 7.68863297563916e-06, 
    1.85258491796887e-08, 0, 0, 0, 0, 0, 0, 0, 4.96666152613617e-20, 
    7.74115856439014e-21, 2.92158200573564e-19, 1.31445158948906e-18, 
    5.43165306748775e-19, 9.22724255847558e-23, 3.95698943410121e-25, 
    5.3821019603374e-07, 0.000106782727079164, 0.000101814363080707, 
    6.34750271845617e-05, 6.03869827019624e-05, 4.17776036533932e-05, 
    1.24567686630961e-05, 2.01411179075922e-05, 1.09438792246006e-05, 
    8.47267325857033e-06, 1.73044920181365e-05, 1.74182440258512e-05, 
    2.10462078749236e-05, 2.81318566626714e-05, 3.70515160310966e-05, 
    4.07345694024871e-05, 2.67559892257925e-05, 1.98109242207948e-05, 
    3.78349963503415e-08, 1.8612098554127e-05, 1.27484887547654e-05, 
    9.33364718763026e-06, 3.60864715884761e-06, 6.99535652844313e-06, 
    4.29918840557521e-06, 1.11278513287641e-05, 7.36324690309732e-06, 
    1.40670478989673e-19, 0, 0, 0, 1.77801536749118e-17, 0, 
    2.37644851845595e-15, 5.33282377536037e-09, 9.762148255884e-10, 
    7.8500978098749e-09, 1.43923767001376e-09, 2.46390849075474e-11, 
    1.94075380881028e-09, 4.4505053631761e-11, 1.89838486201128e-05, 
    8.87742102922994e-07, 2.33353728820667e-05, 5.1972511274716e-06, 
    2.2046620431976e-05, 5.62460379696374e-05, 9.11930774328309e-05, 
    5.25623050764058e-05, 3.20332917809789e-05, 3.54463617324767e-05, 
    3.94194357424344e-05, 2.44823679257117e-05, 8.12705965161012e-06, 
    1.51513073021199e-05, 5.35870277283868e-05, 0.000174930852373565, 
    0.000262733515680473, 0.000204486330287768, 0.000107720574967383, 
    5.35602445016012e-05, 2.11504990155989e-05, 1.65220408348901e-05, 
    9.17522002031397e-05, 0.000439182573520304, 0.000878861643758351, 
    0.000971618266584194, 0.000845203056225714, 0.000601395233324841, 
    0.000366563807073699, 0.000218745074051903, 0.000156410457082319, 
    8.30160290801492e-05, 0.000119185486900329, 2.07450473953831e-05, 
    1.17604242230718e-08, 3.71070485246841e-06, 2.77020664729094e-06, 
    6.47789830639781e-07, 3.71275488436631e-07, 5.85624085533494e-07, 
    8.69120834944511e-06, 4.27209101983662e-05, 1.57316035521811e-05, 
    8.13032093930546e-05, 4.07562403706388e-05, 3.68014483372428e-05, 
    4.60817155736737e-05, 1.67783634287084e-05, 1.28912450381545e-05, 
    1.69339254776561e-05, 1.31343341127171e-05, 5.80441044417061e-06, 
    1.2664352256433e-06, 1.89051832834883e-06, 0, 3.61727755719569e-19, 
    2.03631521204913e-17, 5.41619221208813e-09, 3.06142462774789e-11, 
    9.85987977772481e-16, 7.42166361227755e-18, 4.04314637289158e-17, 
    3.17725320193652e-20, 0, 0, 0, 3.85861208663202e-15, 
    1.32469417947184e-10, 2.0408185042084e-08, 3.10374112538924e-06, 
    3.81904059584438e-06, 7.11190589147297e-06, 3.7824217630109e-06, 
    3.43720747587956e-06, 1.25291297953205e-05, 1.55687281992424e-05, 
    1.3484932485271e-05, 1.57990331057518e-05, 1.60046087882314e-05, 
    1.93012020541236e-05, 9.67967708390119e-06, 8.78943581856247e-06, 
    8.30141387741251e-06, 5.0775878973468e-06, 5.62461032652382e-06,
  3.67885656372126e-06, 9.97522893107002e-07, 1.44463756313244e-06, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2.67619799872879e-24, 1.38061002782746e-19, 
    3.01300351600362e-20, 3.04239423995166e-19, 5.68104993096079e-13, 
    0.000107040150479994, 8.70013986966273e-05, 8.00269997704939e-05, 
    9.25931156262619e-05, 4.28309595801945e-05, 1.62125628214874e-05, 
    2.9348733550003e-05, 1.5959739185305e-05, 9.07344476654142e-06, 
    1.18851987811945e-05, 2.19221937912668e-05, 2.21826266240666e-05, 
    2.02615688359971e-05, 2.05734082885017e-05, 2.36507841943565e-05, 
    2.60034364835989e-05, 2.12857711497095e-05, 1.88907373024399e-05, 
    1.21899948872048e-05, 6.56075533988595e-06, 6.26849784634363e-07, 
    8.53857171346689e-06, 1.09083060232893e-05, 1.09417512259143e-05, 
    8.07854112470088e-06, 2.6846466833111e-06, 3.39207946762478e-10, 0, 
    1.56412451714649e-19, 0, 0, 7.01603021267128e-17, 4.00382632171667e-18, 
    0, 2.39102499983548e-20, 1.34156553788378e-17, 0, 0, 0, 
    7.37234424097866e-12, 1.43875593511114e-05, 1.23098853875093e-05, 
    3.09811446579741e-11, 9.20508910780473e-07, 1.0514664951119e-06, 
    1.35814582340619e-10, 8.55740367779433e-06, 4.2011804917122e-05, 
    2.96291626462177e-05, 2.74913566149175e-05, 2.94194832588821e-05, 
    5.08597415619657e-05, 6.89685542891934e-05, 9.75654177521823e-05, 
    0.000142605695615105, 0.00016196406204168, 0.000186475144963281, 
    0.000143372224578747, 8.20582374058832e-05, 5.64305979326586e-05, 
    5.19717680810184e-05, 0.000220548304315423, 0.000921955938971106, 
    0.00137127156055316, 0.00134300505019925, 0.00112108158361279, 
    0.00068500551139495, 0.000388726024780807, 0.000157858244774235, 
    1.09847343861658e-05, 3.01429454254939e-05, 3.3135821247756e-05, 
    2.47123222543745e-05, 4.45939580138267e-22, 6.56710444134216e-06, 
    8.04182409067589e-06, 7.41712925367547e-06, 5.66017276876031e-06, 
    3.79858078656231e-06, 1.20113305420551e-06, 1.18462006147659e-05, 
    3.10854288712426e-05, 2.0603742811743e-05, 1.40590348676607e-05, 
    2.2288000479888e-05, 2.84515565181455e-05, 2.19493937844869e-05, 
    2.56462760512627e-05, 1.57216425920989e-05, 1.03079550133873e-05, 
    1.06117190752387e-05, 1.04101488669907e-05, 6.51324291451861e-06, 
    2.01127340899977e-06, 2.04835996177536e-06, 8.79775243093617e-08, 
    1.98006350025593e-22, 1.69322463294609e-07, 5.75413876866509e-08, 
    1.97233390037979e-20, 0, 0, 0, 0, 0, 0, 5.73525432726552e-13, 
    2.04530627113898e-08, 1.12507675932073e-05, 4.4111806270553e-06, 
    4.43605763687992e-06, 4.55133364965957e-06, 4.09843640921598e-06, 
    6.53261621030502e-06, 2.47251832010383e-05, 2.52031927877123e-05, 
    2.38986146276723e-05, 1.89194642439676e-05, 2.45416921204158e-05, 
    2.71628460226024e-05, 1.36046659132417e-05, 1.52788601648371e-05, 
    1.35606002080996e-05, 1.33891572033261e-05, 1.06125614972615e-05,
  2.56522936188245e-06, 2.7953974943186e-06, 2.51765317724774e-06, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1.94583109751942e-06, 1.71054833219721e-12, 
    4.3137186206032e-24, 0, 1.32514629993282e-21, 4.25698415098519e-05, 
    4.08675770417558e-05, 9.85146458083425e-05, 0.000101466202586644, 
    9.88956972042222e-05, 6.35015364016444e-05, 4.35739707401984e-05, 
    2.42521351563816e-05, 2.29382238069394e-05, 1.84783255566875e-05, 
    2.0480678857317e-05, 3.43260226028321e-05, 3.79084109991804e-05, 
    3.96050941230078e-05, 4.01378946426848e-05, 3.61829548732696e-05, 
    3.3186176438506e-05, 2.30937807152465e-05, 1.74013842391945e-05, 
    1.87047496969448e-05, 2.16304487027847e-05, 2.29292967149968e-05, 
    1.84841398164416e-05, 1.20105176959644e-05, 4.6609986574764e-06, 
    7.00179271024933e-08, 1.75530232528133e-10, 1.23528826034126e-11, 0, 
    5.81031232230979e-19, 3.79475553550863e-19, 1.11988220928994e-18, 
    4.86818699078263e-18, 1.00087802345772e-18, 0, 0, 0, 0, 0, 
    1.31649194444263e-07, 0, 7.77903616610734e-06, 3.93169556136301e-06, 
    5.36844484432231e-06, 1.12229293186707e-07, 2.35492868257799e-07, 
    3.33476726437744e-06, 1.07355106865642e-05, 3.44821605066271e-05, 
    3.10330991920361e-05, 1.83994245884646e-05, 4.51216599066062e-05, 
    4.24278137355617e-05, 5.52104544535331e-05, 5.5559683338876e-05, 
    2.90742586149534e-05, 2.50135200212182e-05, 2.14648492340784e-05, 
    2.61407073049234e-05, 6.89907515705431e-05, 0.000185399710374923, 
    0.000820791891444948, 0.00114499674107047, 0.000830946666350442, 
    0.000439909577964473, 0.000336106493963289, 0.000214814752679285, 
    0.000105960545321523, 2.62294197081288e-05, 3.25316036059539e-05, 
    1.6911648333449e-05, 2.61608939714633e-05, 4.89428795757644e-05, 
    3.18567176013324e-05, 7.26788611476988e-06, 8.64919585287568e-06, 
    6.66913057559937e-06, 6.54048209295433e-06, 6.19675347583651e-06, 
    1.28877029368374e-06, 1.41031915825724e-05, 9.99221293184392e-06, 
    8.50453717317243e-06, 8.55874284418783e-06, 1.23202518876397e-05, 
    1.26227084825905e-05, 1.93912210699006e-05, 1.53989899842502e-05, 
    1.64498638785016e-05, 9.69442884164826e-06, 1.02817335481103e-05, 
    1.21023786043639e-05, 4.17117120332636e-06, 1.93471137997137e-06, 
    3.28137650766632e-06, 1.6415121067093e-05, 2.73756225113076e-07, 
    6.9108568614146e-07, 1.49874188483459e-07, 7.81816524347847e-10, 
    7.15839642474508e-15, 0, 0, 0, 8.63323561407218e-19, 
    3.57047691595391e-16, 6.72780330844204e-11, 5.14771146849466e-07, 
    4.53720087106269e-08, 3.65641351530046e-06, 8.03873782870298e-06, 
    4.0699756183087e-06, 1.40398033238321e-05, 2.30844092785041e-05, 
    3.13277949222869e-05, 2.61547884464092e-05, 2.62507018823958e-05, 
    2.08353163130841e-05, 2.237536888619e-05, 1.36322213267796e-05, 
    1.59198938662065e-05, 1.1954375911786e-05, 2.18171621655014e-05, 
    1.55107272543323e-05, 5.91081154769803e-06,
  2.12744063172515e-06, 3.00094139160577e-06, 1.65963085009417e-07, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4.62753077088116e-09, 4.72413682538079e-07, 
    1.38311997598822e-06, 2.23593792242378e-06, 8.64483044684385e-13, 0, 
    1.18418068957434e-11, 1.80012886642864e-05, 4.64630432962784e-05, 
    8.16865324373439e-05, 0.000117891103996158, 0.000101994844241054, 
    8.51077497761623e-05, 6.76301392349893e-05, 2.99291943404919e-05, 
    2.32091684421704e-05, 2.20522243654398e-05, 3.29807953632745e-05, 
    3.42604565558951e-05, 3.40199416053573e-05, 3.96015250381912e-05, 
    4.30660037366121e-05, 3.33615535375503e-05, 2.29155396091402e-05, 
    1.81877684686739e-05, 1.9968002657916e-05, 1.92088378223782e-05, 
    5.56928463544136e-06, 5.79890026029309e-06, 3.13990500784992e-05, 
    2.12892807965954e-05, 1.22966165418191e-05, 1.23981053109045e-05, 
    9.17648193599583e-06, 7.93294948150912e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 8.93933784365242e-24, 1.44781407725266e-06, 6.20538459923769e-06, 
    1.6735167320155e-06, 9.61652139140964e-07, 9.38203141011456e-07, 
    5.87906429556482e-07, 3.91849915329953e-06, 5.85978541944145e-07, 
    2.93500678333731e-07, 9.58945315264e-09, 1.13167540820321e-06, 
    2.606515045101e-06, 2.57125326434957e-06, 2.14640302834321e-08, 
    2.19733179204804e-11, 1.81484375213793e-08, 5.25396571379922e-06, 
    0.000155873144984108, 0.000331705922279507, 0.000288869050834031, 
    0.000379790767627002, 0.000438771488455087, 0.000250361266117484, 
    0.000194707120000357, 0.000129545649396707, 8.24031799175301e-06, 
    6.44008422300153e-05, 9.24918684168429e-06, 1.88083747775728e-06, 
    2.10823968774269e-06, 6.25458110837412e-06, 5.60775978779501e-05, 
    2.94029501207131e-05, 2.78394820809613e-05, 5.01409024401503e-06, 
    6.76168526808848e-06, 5.15618677832221e-06, 6.30955268313733e-06, 
    3.62681186393938e-06, 2.34356854429062e-05, 7.56796248812463e-06, 
    6.52116417458994e-06, 6.44275923348477e-06, 5.24148083105465e-06, 
    1.03797712713571e-06, 1.93553242550715e-06, 2.33156326150291e-06, 
    2.20613485003091e-06, 2.05722177108797e-06, 3.52223012108061e-06, 
    5.63593642614599e-06, 6.21044034254926e-06, 4.44848140886294e-06, 
    1.12601214934056e-06, 1.43621209908629e-06, 1.15473212210486e-05, 
    4.45156034528784e-06, 1.55424758484147e-05, 2.22476127084012e-07, 
    4.01228296379201e-12, 0, 0, 0, 0, 1.28986573467212e-18, 
    6.99148682434357e-12, 9.2981737499212e-11, 1.53191718426412e-08, 
    3.69902614910062e-08, 1.64441151337868e-07, 5.12807257662295e-06, 
    7.7987369034014e-06, 1.74824516891309e-05, 1.56150184961117e-05, 
    2.45696852527308e-05, 3.26811037125869e-05, 1.83531904455219e-05, 
    2.39486141185084e-05, 3.25840563903342e-05, 2.64736665122644e-05, 
    2.83368891702907e-05, 2.23878792206986e-05, 1.3375226102274e-05, 
    1.41217476281233e-05, 8.71310279402785e-06,
  1.45199169822762e-06, 3.06398563948061e-06, 8.51981720760065e-07, 0, 0, 0, 
    0, 0, 0, 0, 0, 8.38998453900403e-12, 3.87298146079667e-09, 
    3.28336406069313e-08, 5.59176004897224e-07, 2.02505599720391e-11, 
    6.29718618728797e-07, 5.72851596690063e-13, 1.13001109095253e-11, 
    7.27258301293901e-06, 5.92938318594409e-05, 4.6276521191024e-05, 
    7.26653193326604e-05, 5.81263752400118e-05, 7.25810688339422e-05, 
    5.08692305774134e-05, 2.03380676350665e-05, 2.06176763020262e-05, 
    2.50468896407863e-05, 2.49886102713407e-05, 2.49992491350235e-05, 
    2.81213587777788e-05, 2.72287251914262e-05, 2.67978988778716e-05, 
    2.34492913600474e-05, 3.19969823709028e-05, 5.13077456541912e-05, 
    5.62733090383851e-05, 5.2432431965898e-05, 4.27296052608458e-05, 
    4.30391039215679e-05, 4.34201383038053e-05, 4.71068585704318e-05, 
    3.70566310200184e-05, 3.18895734969493e-05, 2.20127894680697e-05, 
    8.66608595324795e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3.08385408472787e-13, 1.47941126347937e-06, 1.28932791508523e-06, 
    1.28084440308239e-06, 2.20837278286637e-07, 0, 2.61507673486924e-06, 
    1.71669438268098e-06, 0, 0, 2.84879417365996e-12, 7.69748565993175e-07, 
    2.21063228247562e-07, 1.64479290488388e-06, 3.53164627274567e-06, 
    4.97729450195967e-06, 9.58562962523987e-05, 0.000244647778016472, 
    0.000308464214699749, 0.000306332831467006, 0.000289924305691247, 
    8.54199704590652e-05, 4.9502327120775e-05, 3.58252656561839e-05, 
    2.08897429860066e-05, 6.51999874908852e-06, 2.04206504135932e-06, 
    3.71928817767817e-06, 2.79574945848632e-18, 1.64809689514353e-07, 
    1.10564880242683e-05, 2.40013394129843e-05, 2.90169379663656e-05, 
    1.86850189799368e-05, 1.19473517836248e-05, 2.44045816929102e-06, 
    9.65381407848544e-12, 1.59280835814158e-06, 2.64159961661903e-06, 
    1.1717009843571e-05, 8.86500184745842e-06, 9.09007534571237e-06, 
    6.15533131082223e-06, 1.82668620506096e-06, 3.11555902647078e-06, 
    2.8633768597797e-06, 3.39405439189993e-06, 1.67592216668296e-06, 
    1.27815975849461e-07, 6.28129607433615e-07, 1.3237846719861e-06, 
    3.23375419627118e-06, 6.05592203036109e-07, 1.17981715967349e-06, 
    5.94353805207561e-06, 1.03865358156908e-07, 1.48091602894005e-06, 
    2.17841220249498e-05, 1.72001442011186e-05, 2.12051854649854e-07, 
    2.91615336785689e-08, 2.21686445962839e-17, 0, 0, 0, 
    4.68644091140654e-17, 1.40681613561299e-16, 1.13045643629502e-10, 
    4.25614726976194e-10, 2.60153040653402e-06, 3.67229737907933e-06, 
    1.00168535847734e-05, 9.44859302769826e-06, 1.87674060479115e-05, 
    2.55821570288807e-05, 2.92566978554254e-05, 3.24023346004835e-05, 
    2.95893651922704e-05, 1.6846315187502e-05, 3.52383373946886e-05, 
    4.33468398293021e-05, 3.75672396134256e-05, 2.26523328276809e-05, 
    1.11568760282008e-05, 1.05771287524223e-05, 2.33585582557241e-06,
  7.61291796014036e-06, 3.44988917800497e-06, 4.7137429262737e-08, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3.67842118477887e-10, 3.4878930506369e-09, 
    3.65408337041749e-09, 4.4329333191506e-12, 6.29475067599499e-06, 
    1.18209248736148e-05, 1.38135582130139e-06, 5.60904066732317e-05, 
    7.27985337073599e-05, 6.95054895908757e-05, 5.35102113254796e-05, 
    4.81324023520561e-05, 4.43485436395616e-05, 5.38578419811139e-05, 
    4.53647950362213e-05, 2.81977842308624e-05, 1.64162112776232e-05, 
    2.38006981088665e-05, 2.46307801251278e-05, 2.28359892203321e-05, 
    2.44322518072477e-05, 2.98199600462695e-05, 4.76454793268459e-05, 
    5.38279550237857e-05, 8.38179465106277e-05, 7.39686254340695e-05, 
    9.89737660854651e-05, 0.000100910271072883, 9.4733054157424e-05, 
    4.46781466327058e-05, 5.12300123713392e-05, 3.44187295638352e-05, 
    4.26447689517763e-06, 1.0981265551222e-06, 1.05459675812845e-06, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.55566280495789e-07, 8.940076284467e-07, 
    1.34022080949312e-06, 6.30826769735924e-07, 1.93859989326495e-06, 
    5.4167328725099e-06, 1.05687091149436e-09, 0, 3.82116002699553e-21, 
    3.16852899262983e-10, 1.80385228333844e-06, 1.39028544555466e-06, 
    1.96346914878224e-05, 0.00016358163687756, 0.000323745938140712, 
    0.000223169195486419, 0.000196063163167985, 0.000132688814891567, 
    0.00012412842270463, 9.02668769644322e-05, 4.17112167745436e-05, 
    1.11381994038246e-05, 2.70047665557407e-06, 3.47016028377962e-06, 
    1.17830956204377e-06, 2.63563222534597e-06, 1.38058253697314e-06, 
    2.64502509354856e-06, 3.06276644182427e-05, 4.28725650085458e-05, 
    2.41118818034999e-05, 1.0390951929272e-05, 3.59805565076905e-06, 
    2.97924576715198e-06, 8.39699235510922e-09, 7.91496324799123e-06, 
    7.63992550903381e-06, 7.57806205598241e-06, 7.31628200940704e-06, 
    8.52879349129309e-06, 2.06134168681114e-06, 2.17324441776941e-06, 
    1.83467515748194e-06, 1.84894446966084e-06, 1.77289748495484e-06, 
    1.25548135277412e-06, 1.49638684077327e-07, 1.45055317480931e-06, 
    5.63464924972697e-07, 5.60203468139898e-07, 9.64039388545844e-07, 
    1.90729198505553e-06, 7.53182808653815e-06, 1.35199811755385e-07, 
    4.4390745763966e-06, 2.74899816925148e-05, 9.7415151596296e-13, 
    1.80533493540126e-18, 5.26766707356806e-09, 0, 0, 0, 0, 
    4.32665118426619e-18, 3.45030615255855e-16, 7.96784152260996e-16, 
    6.50191332936646e-08, 4.98764184163018e-06, 1.43395041705947e-05, 
    2.93199494424817e-05, 2.50317262377462e-05, 3.17801306579777e-05, 
    2.65328818773359e-05, 2.61213148693021e-05, 2.6674583264278e-05, 
    1.91921040348872e-05, 1.77378452976728e-05, 2.61754006300154e-05, 
    2.28007646430674e-05, 1.96539272293709e-05, 1.73882051347703e-05, 
    5.47579865619301e-06, 8.62303756884605e-06, 4.14167394205517e-07,
  3.17426654525235e-08, 4.75010061483753e-08, 6.3401534145661e-10, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 6.26354040335907e-12, 7.42877557054996e-10, 
    1.34372834215115e-09, 2.98452080094311e-12, 7.38407816792614e-06, 
    1.2577263974857e-05, 3.90921567477748e-05, 5.90852612633591e-05, 
    8.14105048518321e-05, 5.80642292025e-05, 6.4525314094827e-05, 
    3.45219986401621e-05, 2.62542876748698e-05, 2.89785019409876e-05, 
    2.85789772524662e-05, 2.32858472832081e-05, 1.74900942222858e-05, 
    2.68764813008352e-05, 2.52265717757802e-05, 2.01278770469158e-05, 
    3.12663376386255e-05, 3.90914711323785e-05, 4.52762314420216e-05, 
    5.20353737228769e-05, 5.8616398416373e-05, 5.79841690154266e-05, 
    3.93717026357738e-05, 5.00420132433744e-05, 3.69721935186462e-05, 
    4.65504212210591e-05, 2.45499564229722e-05, 9.64507208985547e-06, 
    8.88762145847876e-06, 4.60656954353657e-06, 3.388162360957e-06, 0, 0, 0, 
    0, 8.25263958501514e-12, 2.34794723920713e-08, 6.68672195930645e-09, 
    8.44244401407335e-08, 2.91681276450737e-21, 6.5411797109785e-13, 
    2.03136126674365e-08, 2.86796900447704e-06, 3.86004079800318e-06, 
    2.38809466624894e-06, 4.00801157766167e-07, 3.2940439795726e-06, 
    8.08239846422944e-06, 7.5932300311253e-06, 6.88703799086293e-06, 
    2.42585341564042e-06, 2.13932405562644e-06, 1.79625753690481e-06, 
    3.46835042208045e-07, 9.6459095371446e-07, 5.1005796497629e-05, 
    0.000210721278297761, 0.000287061135556496, 0.000164719650006202, 
    8.81872283694418e-05, 6.74312120108731e-05, 7.93854776674407e-05, 
    4.8999051038849e-05, 2.3673803541317e-05, 6.44921795815281e-06, 
    2.36279375249367e-06, 1.73615861069367e-06, 1.99422332799146e-06, 
    2.76183021438384e-06, 1.21108271463974e-06, 1.48234247521651e-05, 
    2.09379004761312e-05, 1.75502656064361e-05, 1.98111894411419e-05, 
    1.00021320490076e-05, 5.49496939744751e-06, 5.05567053448217e-08, 
    2.61575685825365e-09, 7.76171975133091e-06, 1.37293920343866e-05, 
    6.9422528612516e-06, 3.11454784164295e-06, 4.40625587515074e-06, 
    4.37283476931152e-06, 4.19561388955796e-06, 4.16271349295096e-06, 
    2.2650825323812e-06, 1.76510658267875e-06, 1.58846869821604e-06, 
    1.04106318763404e-06, 3.50285250474829e-08, 8.77414047301432e-07, 
    1.09343228351933e-06, 5.06935754933304e-07, 3.1739156221576e-10, 
    2.0047594150082e-08, 4.4367047123002e-07, 2.82856691226896e-06, 
    1.20623659040673e-05, 3.41985144277224e-06, 0, 8.58280664876919e-28, 0, 
    2.42777493978545e-24, 1.07497165623042e-17, 0, 0, 0, 
    8.54961487291986e-17, 5.15857083135984e-16, 6.00367078839439e-20, 
    9.01536816991124e-07, 2.15321794105488e-05, 4.37346334772669e-05, 
    3.3363175872157e-05, 4.01276311450321e-05, 4.13322896714278e-05, 
    4.22458059659857e-05, 3.45731473160137e-05, 1.73725605588173e-05, 
    2.32843515927218e-05, 2.79657970513937e-05, 2.70217314084865e-05, 
    1.97174964841218e-05, 1.37898492834239e-05, 6.04141730712237e-06, 
    5.5913448260263e-06, 3.46376229424175e-07,
  1.00248052660443e-06, 1.45666466742441e-19, 1.21809616293638e-19, 0, 0, 
    1.85811946105547e-14, 0, 0, 9.63037150401149e-17, 0, 0, 0, 
    5.31639608564481e-12, 1.87298304900325e-11, 3.37427950546321e-10, 
    5.26712117823028e-06, 3.2281481406411e-05, 3.15249087961631e-05, 
    3.23952822654301e-05, 6.25407168498915e-05, 4.52461820031296e-05, 
    4.25621727994078e-05, 5.80654597513208e-05, 6.32918891932798e-05, 
    2.83542795120873e-05, 1.30804453373857e-05, 1.00076048453445e-05, 
    1.40555317295574e-05, 1.28469125518865e-05, 1.69023244035657e-05, 
    1.72134857044885e-05, 2.68279885267618e-05, 3.15145800016247e-05, 
    3.27724113566013e-05, 3.90480374503822e-05, 2.20837995577505e-05, 
    2.5236743635434e-05, 1.36596035561082e-05, 1.21399426914927e-05, 
    2.77115918963743e-05, 9.8855887727489e-06, 1.69097966816829e-05, 
    1.23582392485213e-05, 1.69414172841891e-05, 2.04547474263696e-05, 
    1.02320195768655e-05, 8.89993473792038e-07, 1.97800383723675e-06, 
    1.35443321479643e-06, 8.31542272111139e-07, 1.75017270409989e-06, 
    2.655568634112e-06, 8.64440770802388e-06, 4.09714092352493e-06, 
    2.95355628100048e-06, 3.26761094296037e-06, 4.99116003151848e-08, 
    3.30862756929059e-06, 2.94881485181916e-06, 2.80694334814056e-06, 
    6.58367216595445e-07, 7.38671767766176e-06, 1.67301663723591e-05, 
    4.84180443947768e-05, 5.6304717774326e-05, 3.28199585224744e-05, 
    1.18313802734423e-05, 2.31179520772821e-05, 3.2778043520241e-05, 
    8.83210354636122e-05, 0.000198901739438036, 0.000303978623726939, 
    0.000149294036593485, 0.000101779761140473, 5.64233478666587e-05, 
    1.6597119141026e-05, 1.89432416072351e-05, 2.52455672069579e-05, 
    2.42774708749215e-06, 4.31116494299074e-06, 3.82195004207119e-06, 
    2.68045986202723e-06, 3.15425355448587e-06, 2.85968431376106e-06, 
    7.29152454237038e-07, 1.3095435654165e-08, 2.07392276911593e-05, 
    2.27712761575566e-05, 2.08802330780496e-05, 7.94660700054129e-06, 
    7.78251785777295e-06, 9.75304894213475e-06, 6.64497181991669e-06, 
    6.77982718258826e-06, 1.08392818331751e-05, 1.38068462055624e-05, 
    9.52460627048817e-06, 7.64609145443947e-06, 1.13859523261916e-05, 
    1.39714232591753e-05, 3.35634626104109e-06, 3.7376453695575e-06, 
    2.94123206506825e-06, 2.13562100298064e-06, 1.4248389708223e-06, 
    1.30245292749921e-06, 2.153663570416e-06, 1.59011435730827e-06, 
    8.80057217193072e-07, 9.06721338805891e-07, 1.25795964397709e-19, 
    9.54169901227699e-16, 4.65281098971624e-06, 1.81597298678472e-05, 
    3.74379876772325e-08, 8.42645618205878e-22, 5.00970462054035e-304, 
    1.67554225854368e-53, 1.99856809451436e-11, 4.18692896835266e-21, 
    2.18335308700634e-19, 2.77684790039076e-11, 2.67069906562172e-16, 
    4.78048567961385e-19, 1.86265084775089e-11, 0, 5.16018836553487e-09, 
    3.73218632251963e-09, 6.47231404622241e-09, 7.03108214203436e-05, 
    4.63412571619161e-05, 4.74826961012598e-05, 3.47763524591844e-05, 
    2.559028521178e-05, 2.87534226335847e-05, 3.79293233886312e-05, 
    2.1750526083185e-05, 3.15336822373557e-05, 2.85113409660298e-05, 
    1.72767773230793e-05, 4.26211726885812e-06, 5.21225981558285e-06, 
    2.11073360740923e-06, 1.43910854144601e-06,
  8.63785266417267e-08, 4.56274719808249e-07, 2.03577348070126e-06, 
    2.78992792150078e-06, 3.56604374407136e-07, 2.47469416164498e-22, 0, 
    3.32907232476806e-17, 0, 0, 0, 0, 0, 1.02155801305595e-10, 
    2.07037629884219e-08, 2.33229466045308e-05, 1.65161316694194e-05, 
    1.01621464269995e-05, 1.63632895938394e-05, 2.80829542146249e-05, 
    2.47363773244e-05, 2.03548622158553e-05, 1.9937269142406e-05, 
    3.86200139681542e-05, 2.69915372571651e-05, 3.20059222072077e-05, 
    1.10098389460626e-05, 8.6786457523514e-06, 7.26044169874127e-06, 
    9.45814371038683e-06, 1.52618489536523e-05, 2.01706256028998e-05, 
    2.11926643767312e-05, 3.30075601542515e-05, 3.86427163575944e-05, 
    1.58508998909359e-05, 2.0232054674312e-06, 9.28102821791468e-06, 
    9.07890655410843e-06, 1.43022499490418e-05, 2.2959274294277e-05, 
    7.33037571119439e-06, 1.52555014276675e-11, 1.59610215370746e-09, 
    7.84762915701328e-07, 3.83978407863405e-06, 5.69913032143351e-06, 
    2.21942855186047e-06, 3.60177319645189e-06, 2.56054074325221e-06, 
    9.95434455604245e-06, 1.24510568784754e-05, 1.30340004562691e-05, 
    5.93015939207558e-06, 1.25022828018911e-05, 4.15165022402766e-06, 
    1.05300315321568e-08, 4.5844149030022e-09, 2.26424035394425e-09, 
    1.32266166981406e-05, 2.14543302368447e-05, 2.43675936788862e-05, 
    5.78180016445221e-05, 9.03614158857394e-05, 6.48787320432641e-05, 
    6.30749939520168e-05, 6.77917881479212e-05, 0.000138001431567942, 
    0.000215590535814714, 0.000312374219554351, 0.000271632613848399, 
    0.000151187699320886, 5.81504651949987e-05, 2.33686212990801e-05, 
    1.16797872531563e-06, 1.5997012173532e-06, 2.08560320724602e-05, 
    3.26382634201112e-05, 1.74589575154671e-05, 9.68048798107602e-06, 
    3.65674573536462e-09, 1.45540176626732e-06, 6.88580496181203e-06, 
    3.81005294420875e-06, 1.87833752313435e-06, 6.88684790872595e-06, 
    1.5575967443523e-05, 2.06973154116519e-05, 1.01891061952179e-05, 
    8.12190298818903e-06, 1.19232095573165e-05, 1.10500955530681e-05, 
    1.92816731089608e-05, 1.55088879053991e-06, 9.81620341878469e-06, 
    1.61696872861614e-05, 1.66490674790519e-05, 1.95478515085159e-05, 
    2.13687042153726e-05, 1.26136923221637e-05, 8.52941139338963e-06, 
    3.61016146631579e-06, 2.03759720842308e-06, 1.96971691437596e-06, 
    2.27817941407524e-06, 4.76309530349938e-06, 1.01447294700854e-05, 
    4.92867300027445e-06, 2.86117603404721e-06, 1.37323105205116e-06, 
    2.23135614691746e-07, 1.32697951246493e-08, 2.16825251459427e-23, 
    5.85880224580908e-05, 3.47392627353652e-53, 1.37661150291887e-47, 
    8.24489693976444e-21, 1.4310260626472e-11, 2.31716799192106e-15, 
    3.10942365237966e-11, 5.16100920555977e-07, 3.49063852381312e-11, 
    4.85528932290681e-22, 4.88291685470746e-20, 0, 1.74287136426469e-16, 
    9.52974993329292e-56, 2.72599820515959e-30, 8.80923815250824e-10, 
    4.11133553580198e-05, 3.91433745919248e-05, 4.11988162042996e-05, 
    4.8802721441125e-05, 3.2377940896661e-05, 1.95132251875289e-05, 
    2.27230451393219e-05, 2.86412746694538e-05, 5.86633752506794e-06, 
    9.34695083275689e-07, 7.42746502701976e-06, 4.10372387546033e-06, 
    3.72852570906019e-06, 3.82453190211134e-06, 1.66578847390883e-06,
  4.54179630627521e-06, 5.40537171892812e-06, 2.2128533188369e-06, 
    5.90832813487684e-07, 1.626549768054e-06, 2.55925637473446e-07, 
    2.80845442127402e-11, 5.05442162382491e-11, 1.0308287760195e-19, 0, 0, 0, 
    3.9565928775866e-11, 1.4904749533444e-08, 9.58665795746688e-07, 
    2.69998475469955e-05, 1.94781155795256e-05, 1.50749883719973e-05, 
    5.34855386185584e-06, 1.05176471258976e-05, 1.80153349272063e-05, 
    1.71304099153166e-05, 1.34199872517058e-05, 3.21632978217681e-05, 
    1.06350510320189e-05, 9.02417883906197e-06, 1.03403667978081e-05, 
    1.91097597928726e-05, 1.59922833881503e-05, 1.49641355109421e-05, 
    1.73265949756589e-05, 6.35537833490819e-06, 2.66957135604184e-05, 
    4.29788823825868e-05, 3.50145342579874e-05, 1.56399978358269e-05, 
    1.52685064080831e-06, 5.41289572355811e-06, 7.26923317023216e-06, 
    5.53469569171265e-06, 1.74978902423271e-05, 6.27522775251769e-06, 
    5.67403036447464e-10, 8.27475248600739e-06, 6.43486234410222e-06, 
    5.28559222025386e-07, 7.71714298235128e-07, 2.49327465901925e-06, 
    5.6009606437676e-06, 1.59669098502859e-05, 1.56772189266044e-05, 
    1.34761613376326e-05, 1.46640648888422e-05, 1.34039767672894e-06, 
    2.75205575480079e-05, 2.58792725832924e-05, 2.40206166156576e-05, 
    5.0874119677311e-05, 2.3877502806562e-05, 1.03104447803426e-05, 
    4.56215478872377e-05, 3.53454464122332e-05, 1.49722880016046e-05, 
    9.3923096971354e-06, 8.96739852742194e-06, 8.66832941065689e-06, 
    2.58608124433962e-05, 9.09970317462484e-05, 5.83894316999579e-05, 
    9.59702395980781e-05, 5.22096936419002e-05, 1.029568349598e-06, 
    5.09414473883337e-06, 3.10808092502536e-06, 4.48081681353961e-06, 
    2.2202086970418e-05, 4.47012348636839e-05, 2.7301694737997e-05, 
    3.38970355790738e-05, 1.19645395269913e-05, 3.87272222606964e-06, 
    8.09913053811142e-07, 2.4014764152883e-09, 3.19045286362926e-06, 
    6.20760668455815e-06, 6.9061318239586e-06, 9.71126494352083e-06, 
    6.65698991757313e-06, 1.18815391261938e-05, 1.0847054008078e-11, 
    1.19568438491185e-08, 1.07747189424981e-05, 1.14262126311077e-05, 
    1.21155295539771e-05, 1.54557982662866e-05, 6.42584355978536e-06, 
    1.61403139462281e-05, 2.15156149152984e-05, 1.26217418667774e-05, 
    1.47230572736891e-05, 9.94380115940654e-06, 6.10126406319195e-06, 
    3.59711602242536e-06, 3.39087910321091e-06, 6.65932897932108e-06, 
    8.74803310107208e-06, 1.06174982184994e-05, 1.29025442191499e-05, 
    2.13952080157328e-06, 1.31257575321293e-06, 8.24411907196915e-07, 
    1.90958437896005e-08, 2.24126740807573e-09, 3.07349443778037e-07, 
    5.9896967975106e-09, 0, 3.18884447180225e-10, 3.8002127206808e-10, 
    2.04931729347015e-19, 1.57002177972284e-11, 1.69463805335833e-16, 
    1.66347984852453e-11, 1.28703813972958e-19, 5.03822445455993e-06, 
    6.82123429037425e-16, 4.02273207043757e-16, 1.65866712102075e-45, 
    3.30467982333129e-11, 1.71445093065858e-09, 2.23203135429834e-06, 
    3.04775845577219e-05, 2.17649721555126e-05, 2.27143513975715e-05, 
    1.6588526601022e-05, 2.21551015043111e-05, 2.40513215337486e-05, 
    2.17736239587604e-05, 1.39134007224226e-05, 4.77123459073847e-06, 
    3.66254282184939e-06, 9.69034060474591e-06, 8.93610093064244e-06, 
    1.14073039931027e-05, 6.48220582684962e-06,
  7.06545186041171e-06, 1.43177471153758e-05, 2.78519992706833e-06, 
    1.35750340991397e-05, 2.96197523857234e-07, 2.05578475802793e-10, 
    6.53334123732134e-11, 7.99052648880988e-08, 1.92224935451057e-08, 
    1.09712709034878e-06, 6.29453261511789e-07, 1.86893667873329e-11, 
    3.21929404470958e-22, 4.75917150624554e-09, 2.84690986781399e-08, 
    1.6751045283424e-06, 2.08930129672507e-05, 1.82423823909976e-05, 
    1.07027521197411e-05, 9.56924296549594e-06, 2.35641740892674e-06, 
    1.26327338012715e-05, 5.37634294456297e-06, 2.21187446810252e-05, 
    3.35137844137659e-05, 6.58078532313526e-05, 2.24184952246289e-05, 
    5.10881596793853e-06, 1.25563893747261e-05, 5.95411582831388e-05, 
    7.5201566002105e-05, 7.33143856751981e-05, 0.000132124718451183, 
    0.00015947942137345, 0.000177571075039382, 0.000117920116657516, 
    6.71625548613705e-05, 2.58404769556373e-05, 1.45753806223268e-05, 
    1.00936491028925e-05, 1.96624239262682e-06, 5.59462531197097e-07, 
    1.33110117571726e-06, 6.87799150735339e-06, 1.52507966246825e-06, 
    1.32185553423199e-06, 4.71713107412499e-06, 8.06916603959537e-06, 
    4.52514364043269e-06, 1.40268919223813e-05, 2.3456164912506e-06, 
    3.39240767787632e-06, 3.64288172615726e-06, 7.93163376166299e-09, 
    3.66704860585878e-07, 2.62137806426771e-05, 0.000125235343994514, 
    8.52219870769058e-05, 4.88061752571582e-05, 3.48114236960427e-05, 
    1.52437788941013e-05, 7.18305594054687e-06, 0, 5.54480464866587e-07, 
    2.5293455675599e-06, 1.10708378666401e-05, 1.66449812751064e-07, 
    8.70351899496275e-06, 4.75306870413068e-06, 4.51034228973259e-06, 
    9.24952138797538e-06, 8.395939214431e-06, 2.39040419476033e-05, 
    1.69444503275692e-05, 1.13961290998756e-05, 2.19340318508215e-05, 
    1.06463755814205e-05, 1.88198141172122e-05, 2.68239220281707e-05, 
    1.11274566185869e-05, 2.42680077166958e-05, 2.13865244853334e-05, 
    3.20956632043516e-06, 1.06273808382943e-06, 9.9152719568292e-06, 
    5.9343388980461e-06, 5.27271570506547e-06, 5.34458508288506e-06, 
    4.11074834329008e-06, 0, 6.26314875161355e-06, 1.03519243985629e-05, 
    9.80992948459722e-06, 8.33362854021597e-06, 1.26684945919282e-05, 
    9.09762604996172e-06, 1.66982152889978e-05, 1.73959765740945e-05, 
    1.3683001083338e-05, 9.75530213701658e-06, 5.97700097341594e-06, 
    4.01422993975324e-06, 5.8590422514279e-06, 4.46773958305502e-06, 
    8.53082544294114e-06, 1.69763986233002e-05, 1.50319240076429e-05, 
    1.33169193223382e-05, 2.59627785316003e-06, 2.39805135803122e-07, 
    7.33554899959973e-07, 3.22577421386624e-07, 2.09844251926677e-08, 
    6.0132198829683e-06, 3.67990834099947e-09, 0, 1.57299056791295e-08, 
    2.38216812395688e-08, 1.91128014231903e-10, 7.71818581549447e-09, 
    4.43490444730136e-09, 5.56812563473984e-06, 5.51982909627473e-08, 
    1.54462824690296e-17, 0, 2.04860826685783e-16, 1.33795854744649e-17, 
    5.89872656721682e-10, 2.02889277118117e-07, 1.04120884238839e-05, 
    7.97136218162688e-06, 4.19734223490384e-06, 5.03987460636005e-06, 
    1.59743155262578e-05, 2.17263741270617e-05, 2.0873593029922e-05, 
    1.01658751516968e-05, 4.79566305811022e-06, 9.22908912875465e-06, 
    7.21693112797925e-06, 9.62967007715557e-06, 1.00779319257863e-05, 
    1.38704091724155e-05, 9.23331893375358e-06,
  6.88242166655547e-06, 5.41735511043552e-06, 2.27540675312469e-06, 
    1.86104206801783e-07, 1.46373866189134e-06, 5.92539468897272e-09, 
    2.11954995546576e-10, 5.22639682893157e-07, 1.39428050425528e-09, 
    8.11920516333922e-06, 8.56754278156517e-06, 1.58634277732669e-06, 
    1.00499673998503e-08, 5.65180145648536e-10, 2.4571865709916e-09, 
    2.50767896385438e-10, 5.40659143571365e-06, 1.77607930014921e-05, 
    1.10574324835446e-05, 1.71534608124838e-05, 1.37284740410345e-05, 
    1.87082038004303e-05, 2.04870910696734e-05, 2.58338380814207e-05, 
    1.38638095590504e-05, 7.22836437046021e-05, 6.98042313793984e-05, 
    3.40201080657921e-05, 8.55403518386937e-05, 0.000224908046317825, 
    0.000260250366998268, 0.000351162053549534, 0.000354959686943153, 
    0.000239393379261453, 0.000209531835500422, 0.00019048459096611, 
    0.00014364062198499, 2.37998825651942e-05, 7.22117610468792e-05, 
    1.62298929563255e-05, 5.44341459511569e-29, 1.00789571470556e-06, 
    3.0234570779584e-06, 8.14008552499405e-06, 4.71153268033408e-09, 
    7.93161941109753e-11, 3.09772842746974e-05, 4.51823087407575e-06, 
    9.56927302280221e-06, 9.50614652994697e-06, 5.1926128241739e-06, 
    1.88316179466285e-06, 4.81792422853094e-06, 1.52893369335973e-05, 
    5.20572546686443e-05, 8.37679823178943e-05, 6.70677144896446e-05, 
    2.60764426248918e-05, 3.00672553145538e-05, 2.2032986982239e-05, 
    1.02979282691043e-05, 2.82820728733514e-06, 1.53108431143447e-05, 
    4.09907637514425e-06, 4.3284233069454e-06, 3.73268390248863e-06, 
    4.01448954978129e-06, 3.1441909925952e-06, 2.62269854352837e-06, 
    2.27453135673448e-06, 2.94894900763356e-05, 5.46014995683177e-05, 
    5.82704238869852e-05, 1.92472695203784e-05, 5.96902065829472e-06, 
    7.25521603321718e-06, 6.9014437705512e-06, 7.31401255270587e-06, 
    5.47772666984007e-06, 9.2815863809515e-06, 6.91929701558219e-06, 
    6.07828751947534e-06, 1.3380385656369e-05, 1.23895299921547e-05, 
    9.78580305353491e-06, 6.4079139300072e-06, 5.95591966542731e-06, 
    3.21658090134131e-06, 3.23411642978952e-06, 3.66160030473509e-06, 
    8.9987576046439e-06, 8.97061844368773e-06, 8.36882298631523e-06, 
    6.35961380590485e-06, 1.2933443715013e-05, 8.41984460202999e-06, 
    1.14213686832018e-05, 9.19708415034976e-06, 5.58754894637811e-06, 
    6.88676669974393e-06, 4.74480849536385e-06, 2.67590856262879e-06, 
    1.1251806780534e-06, 7.70312755849483e-06, 2.60157833373433e-06, 
    1.54436075747153e-05, 1.58557960825531e-05, 1.04622099817782e-05, 
    2.18642089898279e-06, 2.9845465936464e-10, 1.68694239596074e-06, 
    4.72680206357142e-08, 2.97320340798132e-08, 1.12958187746996e-05, 
    1.33259133319023e-07, 2.96266235461866e-08, 1.6998363568109e-07, 
    1.2569668402388e-06, 4.54609897057318e-10, 1.96595047965097e-07, 
    5.41120276869899e-09, 1.46833827475294e-05, 4.08652542756003e-06, 
    1.55115739611129e-05, 2.63911442839692e-20, 5.31431464144393e-17, 
    1.8971936032092e-07, 3.26942329983197e-06, 2.62077076357266e-07, 
    5.38172393075979e-06, 5.83788083505008e-06, 4.99472538827799e-06, 
    4.58229677132087e-06, 1.60015570915195e-05, 1.55204164715328e-05, 
    9.45756494626273e-06, 1.03649685531497e-05, 7.09295152493346e-06, 
    1.39042218150251e-05, 1.73060566872846e-05, 1.00378484159337e-05, 
    1.0771832709077e-05, 6.01743178146247e-06, 6.55112077228897e-06,
  1.18657440800797e-05, 9.8356178903775e-06, 3.95339798705062e-06, 
    4.77451714495019e-08, 1.26498113141785e-06, 4.46454753710494e-08, 
    4.85425471311894e-11, 5.29531224474787e-07, 2.77739517225788e-11, 
    8.34358030777493e-07, 6.15682106666546e-06, 1.13585951887338e-06, 
    2.00359885320687e-08, 2.37604063154233e-09, 1.31707636925379e-08, 
    7.32048209964524e-11, 6.14719110009615e-06, 2.69178597721751e-05, 
    1.04550482890829e-05, 1.7850112550086e-05, 2.10139462035433e-05, 
    2.30490861332555e-05, 8.65721623085561e-05, 9.70970810587965e-05, 
    6.98532674894883e-05, 0.000115475648626228, 0.00019411516683042, 
    0.00012371807154944, 0.00010569142923572, 0.000191297674790745, 
    0.0003422299023724, 0.000373129705615441, 0.000322973498796137, 
    0.000119844042951509, 8.81070430881454e-05, 0.000113277604428367, 
    1.63306236888549e-06, 2.10224294706395e-05, 0.000123784743903007, 
    5.23026175541091e-05, 8.62901068829807e-18, 7.60567626654076e-06, 
    1.48062727619167e-05, 1.78542249464287e-05, 5.99205056147891e-10, 
    2.02085495578226e-10, 2.74080015523639e-05, 1.3035225995015e-05, 
    9.30556784308414e-06, 1.33956016498277e-06, 2.12545080783796e-06, 
    7.32705891553967e-07, 4.44798018934729e-06, 3.73561845788173e-06, 
    2.06900913640135e-05, 4.02704232628375e-05, 2.66597743177944e-05, 
    3.02378615519533e-05, 4.35320324913101e-05, 3.37570317104766e-05, 
    1.53428370924619e-05, 9.26880793424501e-06, 5.45026258358701e-06, 
    3.43316732378808e-06, 2.27491244527299e-07, 7.1425200953625e-06, 
    9.90929161775585e-06, 5.88960675500509e-06, 7.62415511258103e-06, 
    1.93831489269858e-05, 5.74061247091094e-05, 9.92673093695849e-05, 
    8.24260377416466e-05, 3.32085707433796e-06, 5.43789293286481e-07, 
    9.0568111778062e-06, 5.0061429801992e-06, 2.50715235770527e-06, 
    8.73862026517152e-06, 1.69697327598108e-05, 1.8613066757351e-05, 
    1.45978648942851e-05, 2.06799897398815e-05, 1.77058177559771e-05, 
    2.24405175202253e-05, 1.61763182659327e-05, 1.41435036146613e-05, 
    1.10802247845439e-05, 9.31029523138002e-06, 9.3383644108648e-06, 
    8.32582946487644e-06, 6.86463643128939e-06, 5.79553242507852e-06, 
    5.42540589714211e-06, 5.60911565012738e-06, 3.43905373291537e-06, 
    6.15566557761601e-06, 6.95349062516239e-06, 5.63328537219193e-06, 
    4.28600648518277e-06, 3.37909468491235e-08, 1.53396185461003e-06, 
    1.05323232693854e-06, 1.75861459714848e-08, 6.77725583233065e-06, 
    8.70259856236052e-06, 6.77272676117862e-06, 7.77571083474011e-06, 
    7.84337989249062e-06, 1.41145651023034e-06, 2.04662178139497e-06, 
    1.07057568039095e-05, 3.33220572599618e-08, 1.97896936953198e-05, 
    9.12794884035903e-08, 0, 3.65043820068686e-06, 3.31237857874627e-06, 
    1.39593659276401e-05, 1.79507635601211e-05, 1.6354371470398e-05, 
    2.41191464321822e-05, 2.71225356511599e-05, 1.09290520919425e-05, 
    3.57944065336591e-06, 3.38377861269999e-09, 2.78275985912559e-06, 
    5.02002043542758e-06, 4.64842540400309e-06, 9.76033995737947e-06, 
    1.02507701363591e-05, 1.37273508851649e-05, 1.74375175405145e-05, 
    1.51937846074716e-05, 9.4838667199344e-06, 6.68909138721856e-06, 
    3.2860111741825e-06, 8.44303561328356e-06, 7.37082448004107e-06, 
    7.33668187731759e-06, 8.94156214471158e-06, 1.31225115482159e-05, 
    8.02835617139256e-06, 4.17912800575528e-06,
  4.88879253038466e-06, 7.69561932088741e-06, 9.44570994412009e-06, 
    3.72689410064168e-06, 8.74384548713163e-07, 6.34698089569249e-08, 
    1.57437266910652e-09, 5.77672995998795e-07, 1.13297996067669e-09, 
    7.95272945453015e-10, 1.61878376902759e-08, 3.14579283482422e-07, 
    1.03496004993622e-07, 1.00415024526555e-10, 5.31993988837095e-12, 
    1.88169920167662e-15, 4.27285804180902e-08, 1.27965298214981e-05, 
    2.91681030874674e-05, 3.07807030270218e-05, 2.55733888682067e-05, 
    3.47897333484789e-05, 9.77403060719936e-05, 0.000122877807275879, 
    0.000109343751043528, 0.000112367770648509, 0.000136723897749199, 
    0.000207626403034345, 0.00028569871959655, 0.000269281093854333, 
    0.000366294010852448, 0.000360980483929859, 0.000311451256490292, 
    0.000296441339118854, 0.000184186469737502, 0.000117328450089361, 
    0.000105487859914245, 3.03835557046827e-07, 0.000156638872027493, 
    3.62048040531473e-05, 3.76563236112824e-06, 3.72188512786552e-05, 
    5.33320442868889e-05, 5.13909592737086e-05, 1.75340405100868e-05, 
    2.26750500880586e-05, 3.02774636368164e-05, 3.41444162444292e-05, 
    9.37509721226715e-06, 1.21280837558663e-05, 5.34931617726121e-06, 
    1.29699486556443e-06, 4.35267438190612e-06, 9.56702720403259e-07, 
    1.55680158713502e-06, 6.41738445443066e-06, 1.12155477523133e-05, 
    1.5846394190652e-05, 3.74354512517807e-06, 8.98167633465325e-09, 
    2.48453606979553e-06, 2.70556242712861e-06, 1.1412652979418e-05, 
    1.16175488668341e-05, 1.35630639145142e-05, 2.61483770648917e-05, 
    1.84508815538605e-06, 1.77556400495997e-06, 1.91818665749068e-05, 
    2.20996194359341e-05, 4.62498262310327e-05, 0.000131121860998152, 
    0.000221544655377214, 7.89710335514827e-05, 4.26971577300849e-05, 
    7.2916708315563e-05, 8.55023998844236e-05, 7.82068869017953e-05, 
    7.77344093857799e-05, 6.22062304725847e-05, 5.04194278176196e-05, 
    4.01714443996196e-05, 3.03031424652066e-05, 4.73992945863766e-05, 
    5.23490448313322e-05, 4.09942482487575e-05, 3.07908375628753e-05, 
    2.13494239342607e-05, 1.79447285967093e-05, 2.19466578796793e-05, 
    2.36672733564173e-05, 1.17059645482155e-05, 9.62439023553692e-06, 
    9.20477093937308e-06, 1.06620953608117e-05, 1.08498655824128e-05, 
    7.44962305253191e-06, 6.38589378891904e-06, 3.06632090222814e-06, 
    5.11207569207514e-06, 4.04122868189931e-06, 2.29885558986637e-06, 
    4.60948446402391e-06, 2.06645058714635e-05, 9.34831526083702e-06, 
    9.55057991920209e-06, 1.38999588236692e-05, 1.85731538839792e-05, 
    1.80545991251693e-05, 2.72971786148764e-05, 9.63056933652166e-06, 
    8.44510935141838e-07, 3.86620155171846e-08, 7.51212503126296e-09, 
    5.09602464895096e-06, 1.69407817865485e-05, 3.97274391704466e-05, 
    3.8711318034289e-05, 5.59600395410584e-05, 2.08220066745965e-05, 
    7.37454510768303e-05, 3.84408895879882e-05, 3.04410869755773e-05, 
    5.0465039433536e-05, 1.32252440938713e-05, 3.69050540730661e-11, 
    5.96562907559726e-09, 2.09718292589395e-06, 3.58505539049882e-09, 
    4.7258222325054e-06, 6.93014651559365e-06, 1.9768166684194e-05, 
    3.79227003623723e-05, 2.21698256143686e-05, 1.33244176570741e-05, 
    1.21079927614363e-05, 7.69751971468921e-06, 1.04527151479667e-05, 
    1.23976517902638e-05, 1.49240389691098e-05, 1.74880499309564e-05, 
    1.09756676890438e-05, 1.39668588555715e-05, 7.25595828956479e-06,
  1.53912012683786e-06, 1.04891350056083e-05, 1.25619807576177e-06, 
    1.836710291356e-05, 2.01997549143396e-08, 1.46419336391509e-08, 
    4.434543778677e-08, 1.12536237593324e-10, 8.84691083318653e-10, 
    9.44711368197887e-14, 3.70779161173285e-11, 3.18913508374758e-09, 
    2.09617991033916e-11, 1.54908113818907e-18, 5.23302053456589e-10, 
    5.81628254399363e-09, 3.53713900957629e-09, 4.74101561346321e-08, 
    8.69442193181911e-09, 2.04682904999251e-05, 2.04782871999343e-05, 
    1.45537290759051e-05, 5.16888543142392e-05, 0.000173283114782018, 
    0.000186988532602741, 0.00013414503019916, 0.000222280758413788, 
    0.000219503873674343, 0.000260847755647929, 0.000275333208831862, 
    0.000288726720625402, 0.000326152369360341, 0.000215254766835664, 
    0.000146158511875156, 0.00012440959129009, 9.83845732200308e-05, 
    7.7724018633079e-05, 6.42539304210856e-05, 4.64288027503962e-05, 
    8.78370096993713e-05, 2.06564812918813e-05, 0.00011470572215045, 
    0.000151576228007757, 0.00019362949620517, 0.000146604075051922, 
    9.40052717915204e-05, 5.19158099244635e-05, 1.84488652573642e-05, 
    1.49621592347187e-05, 4.33435405800879e-05, 2.1837689818627e-05, 
    3.8829440169666e-06, 7.65486012003222e-06, 8.59072187728893e-06, 
    9.87734397582584e-07, 1.48336463086866e-06, 7.1973988069979e-10, 
    6.80834604790132e-07, 3.72188680344246e-06, 2.74483944073009e-05, 
    5.04948717258032e-05, 1.27887712041231e-07, 2.39842865535697e-05, 
    9.54794949680345e-06, 2.24519984201667e-05, 3.7962718980891e-05, 
    4.13943246960225e-05, 4.95118345584967e-06, 1.48264110303247e-05, 
    4.34832408656704e-05, 5.11683115681742e-05, 0.000158699582953045, 
    0.000357341516205015, 0.000370514391851671, 0.000260624703528196, 
    0.000289016217514203, 0.000284654760511942, 0.000383267323599169, 
    0.000378903690946826, 0.000259065581881101, 0.000151576924814589, 
    0.000100259249845109, 8.43004386508747e-05, 8.07356770540869e-05, 
    5.89909818671011e-05, 4.79193385831478e-05, 6.57415206570914e-05, 
    6.21037409164686e-05, 3.48541190634112e-05, 3.26948828600643e-05, 
    2.86021555009528e-05, 3.87608870787993e-05, 3.72612880897712e-05, 
    3.23430126752903e-05, 3.27884045459305e-05, 2.91014001120424e-05, 
    2.84846921562076e-05, 2.03722486995946e-05, 2.40323976210401e-05, 
    2.18816991990493e-05, 1.67173522865699e-05, 2.67643375556894e-05, 
    3.43402158320601e-05, 3.5481424705505e-05, 3.09879924812666e-05, 
    3.18779517750339e-05, 3.10884764165468e-05, 3.3725772785242e-05, 
    4.80976703540358e-05, 6.34085426085594e-05, 4.3828495186591e-05, 
    4.5740133668526e-07, 3.19618557566869e-06, 1.39048046237925e-05, 
    3.52024179960881e-05, 9.17671556228787e-05, 0.000115602880457201, 
    0.000117039554756931, 7.83592441588248e-05, 9.16377088128138e-05, 
    0.000120320640023992, 9.19179107387317e-05, 9.5151475905618e-05, 
    0.000155717668178985, 4.85552627734815e-05, 3.1131981577728e-05, 
    8.80561232777369e-06, 3.39952300301695e-06, 4.81211471689406e-06, 
    4.58161859985447e-06, 1.51250641503173e-05, 1.10138656531668e-05, 
    2.24222838428547e-05, 4.17575145014417e-05, 4.83940725910637e-05, 
    1.93913639067385e-05, 4.01136243277062e-05, 2.77026116658925e-05, 
    2.93564458134186e-05, 2.67154304617181e-05, 1.36930835828076e-05, 
    1.11970740192959e-05, 9.73528950398663e-06, 1.79067119324696e-06,
  8.02120394481049e-07, 1.47194158017354e-09, 1.30888283729853e-05, 
    2.83228134070272e-05, 2.30721753572701e-05, 4.42896441362275e-05, 
    2.63756159802965e-05, 2.79019653176873e-05, 0, 0, 0, 0, 0, 
    2.67270471265188e-05, 2.50239855616015e-05, 2.6748141508419e-06, 
    5.17069591956143e-08, 2.21033582418982e-07, 3.9540135404268e-08, 
    1.51068075200046e-07, 1.36588253252441e-18, 2.35718963856259e-18, 
    1.7927302784332e-05, 9.09346660615642e-05, 0.00017223621573694, 
    0.000453905112241186, 0.000409916390013804, 0.000263524460551455, 
    0.000192674662051682, 0.000121653674810348, 0.00012306395259912, 
    4.49298010836764e-05, 4.34533600547678e-05, 0.000107742298194164, 
    6.19219645357101e-05, 0.000151715438601923, 0.000121151120732019, 
    0.000110119554158688, 6.15547859545621e-05, 2.33462342399232e-05, 
    9.98643324054177e-05, 0.000108868230562827, 0.000181444609051996, 
    0.000265873625858564, 0.000282667537549428, 0.000263514113210992, 
    0.000158257595902388, 3.91018465103609e-05, 7.54936370556319e-05, 
    5.55211255032655e-05, 4.4186091090416e-05, 1.79056044261171e-05, 
    9.62453994039335e-06, 1.66411181471446e-05, 1.04683701246089e-05, 
    3.75926480806519e-06, 1.5627323776602e-06, 2.9972832273973e-06, 
    8.72072282174123e-06, 8.26007624292668e-07, 1.67790640413169e-05, 
    4.44244251718579e-05, 5.40696641916652e-05, 1.04599213809345e-05, 
    2.46053415448954e-05, 3.67166845588115e-05, 1.11533426610436e-05, 
    2.1968451687443e-06, 1.21330449414298e-06, 6.04042182160207e-05, 
    8.89714361543361e-05, 0.00026115315744083, 0.000335988955186904, 
    0.000350395830766398, 0.00032436001612272, 0.000299913754378293, 
    0.000293869775115907, 0.000280853920125721, 0.000264809457002654, 
    0.00024801475161829, 0.000226134030452137, 0.000134161193845285, 
    8.72570528796318e-05, 6.87431072307502e-05, 5.28464847696775e-05, 
    4.40961496936156e-05, 6.28432880085068e-05, 6.11471277415102e-05, 
    4.82863822286529e-05, 4.90019297597685e-05, 4.81168158692136e-05, 
    4.80638813348818e-05, 4.70151265749427e-05, 6.21820719098065e-05, 
    4.23132975861107e-05, 4.00554814165856e-05, 6.25899840779202e-05, 
    6.22489199279489e-05, 4.81271339717152e-05, 9.03042811708926e-05, 
    8.09825687659866e-05, 0.000100707964408344, 0.000112963449212618, 
    0.000132257782740134, 0.000158221136827333, 0.000102817992453501, 
    5.15038641690542e-05, 4.28826061996595e-05, 2.71180359918847e-05, 
    6.57614348163213e-05, 8.77435388130801e-05, 4.30805560101453e-05, 
    7.80846176375345e-05, 3.11017477374962e-05, 9.71498224023232e-05, 
    0.000228609367699873, 0.000164172422063783, 7.46790442668615e-05, 
    6.98307076262876e-06, 7.46287168959696e-05, 3.01093549875564e-05, 
    0.000108163911792696, 0.000131117601279633, 0.0001475622711415, 
    0.000110741579487013, 0.00010929424066027, 3.17039995392195e-05, 
    2.08564317415993e-05, 1.81997332408695e-05, 1.94629922164307e-05, 
    1.88155425212787e-05, 2.55768694613712e-05, 2.50098628365645e-05, 
    2.34562081172959e-05, 3.72066811130845e-05, 3.14782291441897e-05, 
    4.8532135354666e-05, 5.54951541492543e-05, 6.29355202653108e-05, 
    5.8086038870059e-05, 1.82402216286009e-05, 1.02907097570485e-05, 
    7.14640354777129e-09, 9.01064332719985e-10,
  2.09875372061088e-09, 4.81706374556641e-06, 3.26146794283351e-05, 
    2.24074828006573e-05, 1.52548333453355e-05, 3.43734638229393e-05, 
    2.56705149312457e-05, 2.68629899760006e-05, 3.65003169469654e-05, 
    3.31281244544855e-05, 1.26904497035799e-05, 0, 1.42003738564572e-05, 
    4.88921533692516e-05, 5.06704940156339e-05, 4.24020861957279e-06, 
    3.0893509216804e-07, 1.22892179740542e-05, 3.74248845034502e-09, 
    3.60649136071058e-16, 8.79677539371151e-19, 2.58187025236633e-05, 
    6.90621558640023e-05, 1.75289336119493e-05, 0.00015722304321977, 
    0.000323546058009588, 0.000356044269813026, 0.000233249384122213, 
    0.000160863841447619, 0.000139283553479472, 9.31234962849529e-05, 
    4.75754621163099e-05, 0.000110912221723203, 0.00012369195079478, 
    0.000143393492674414, 4.70531393081021e-05, 0.000154117881265853, 
    0.000132909402486391, 0.000125401747940721, 3.70839748758121e-05, 
    6.90680914951179e-05, 9.22994032468645e-05, 0.000140403283981629, 
    0.0002112375884491, 0.000487109639700608, 0.000520531326470881, 
    0.000387724153794178, 0.000146237362363591, 0.00012398370426604, 
    3.97146923583271e-05, 4.15263278432936e-05, 1.46163239776322e-05, 
    1.86280546043639e-05, 2.88718933497874e-05, 3.01588733409468e-05, 
    1.7117749159559e-05, 3.01064813250367e-06, 2.11150740201264e-06, 
    3.20301059122082e-09, 6.04204491289887e-06, 1.73485491649948e-05, 
    4.58985903049412e-05, 3.35215618053447e-05, 9.45185707944423e-07, 
    8.1560957702893e-06, 4.41268006429961e-06, 8.14043937617843e-07, 
    4.56291139446371e-07, 9.52725464830028e-07, 1.87393997979361e-05, 
    0.000155879378426529, 0.000272127912837374, 0.00027539735790434, 
    0.000255519196004815, 0.000138046072553509, 0.000118191839396533, 
    8.32106305384969e-05, 4.73299645110725e-05, 5.63652855098366e-05, 
    7.22738483528545e-05, 8.135542035339e-05, 8.21775498764577e-05, 
    7.13707674498779e-05, 6.80515082442388e-05, 3.73919024020872e-05, 
    2.095811725605e-05, 3.79132616331456e-05, 5.61852749389245e-05, 
    6.21504177627912e-05, 7.55282758131444e-05, 5.2549266487479e-05, 
    3.41240421876331e-05, 5.66205735815188e-05, 2.92249029160942e-05, 
    2.09000463875954e-05, 2.07216440654704e-05, 2.84823118358341e-05, 
    2.38097998389296e-05, 5.8855283711393e-05, 3.90837143506119e-05, 
    0.000103829989564216, 0.000132294136946816, 0.000243306697721927, 
    0.000276042657230522, 0.000281010266705433, 0.000126814715928514, 
    5.01430566007874e-05, 3.06299801783067e-05, 1.30188284142481e-05, 
    3.15322081612057e-05, 0.000174837109801311, 0.000229050087824264, 
    0.000234486366745916, 4.14826352769406e-05, 9.56695905922129e-05, 
    0.000143720211387361, 0.000146855503476698, 5.23252176509465e-05, 
    2.89652131850501e-05, 5.74931826347107e-05, 2.07679563758642e-05, 
    1.35433031289669e-05, 2.09964749666521e-05, 0.000131660048455233, 
    0.000149241034099822, 0.000155980527176117, 0.000167410410846564, 
    0.000194191621682524, 8.49991875339316e-06, 0.000173567389983868, 
    7.92135000068658e-05, 4.61767029700943e-07, 1.39188254527741e-05, 
    2.11225511555624e-05, 2.28618447374066e-05, 2.78827621574349e-05, 
    3.05641778938357e-05, 7.71496252521411e-05, 0.000198085272176657, 
    9.56117077423899e-05, 1.61515792807397e-05, 1.31125508639856e-05, 
    1.13888091501957e-06, 3.915121390041e-20,
  1.20123033966404e-09, 4.5112801817706e-17, 3.72099053877157e-06, 
    1.34668631663849e-05, 2.04116495438981e-05, 2.05337627171443e-05, 
    3.0414877751955e-05, 4.21565292871623e-05, 4.45228187285438e-05, 
    3.317400257859e-05, 4.73188707446166e-05, 2.85241996783066e-05, 
    1.17670046944582e-05, 2.92290154208812e-05, 1.47252859551486e-05, 
    9.89882658965017e-10, 1.07724605199774e-09, 1.12440161074399e-09, 
    7.18395149010529e-09, 1.35072199079658e-06, 1.03370586541352e-07, 
    5.76212644410713e-10, 2.74989265747924e-06, 8.01581048795959e-06, 
    0.000158709990394855, 0.000188797248137849, 0.000260740462172492, 
    0.000279472759008052, 0.000296844081931237, 0.00023728035698963, 
    0.000222594323064097, 2.14829125422312e-05, 0.000101663554480213, 
    0.00023105792907735, 0.000192134220426764, 0.000257255972055851, 
    0.000221102879492024, 0.000241633053464335, 0.000170537197266205, 
    3.94042518762176e-05, 0.000113202009523224, 0.000131455807053849, 
    0.000147463410532222, 0.000204395429289673, 0.0003799066273296, 
    0.000437956107228903, 0.000348752181692029, 0.000196434358671009, 
    0.000174181047741713, 0.000168286466580907, 6.12419714051956e-05, 
    3.33355815222939e-05, 3.49455373844281e-05, 4.55753823468237e-05, 
    5.17659098671299e-05, 4.55027119475991e-05, 3.5440801403846e-05, 
    3.2464654875278e-05, 5.54602269083767e-07, 8.98863334640573e-06, 
    6.00647314067209e-05, 0.000113540472337698, 0.000136281790236477, 
    3.0472546518433e-05, 4.5376138295556e-06, 1.06344528992564e-06, 
    2.6964196797949e-07, 1.0592848154798e-06, 1.14867961387473e-05, 
    6.67293084725373e-05, 0.000181144097332677, 0.000165937298531241, 
    0.000111971770991537, 8.13922733980744e-05, 4.07666219633069e-05, 
    2.75031250802233e-05, 3.37014430272915e-05, 3.71352558390773e-05, 
    3.30645449104324e-05, 3.7688194497935e-05, 3.17284082865774e-05, 
    3.02965271029969e-05, 1.7737477329165e-05, 1.72272272587983e-05, 
    4.14106998394074e-05, 3.6940640114751e-05, 3.86224250358337e-05, 
    3.7640676568686e-05, 7.9740789308476e-05, 0.000104808177517484, 
    6.43673803038834e-05, 7.16134379040894e-05, 0.000104223005353082, 
    3.42589348106966e-05, 4.21859191608458e-05, 2.08372874295022e-05, 
    1.90030592174376e-05, 2.40259052039931e-05, 3.30503655444072e-05, 
    2.12495536658894e-05, 8.17222735502863e-05, 0.000129961518737824, 
    0.00017446322214894, 0.000111991807917362, 0.000215740088166112, 
    0.000148963567704056, 0.000113113825928058, 8.66011848346622e-05, 
    7.5483541748108e-05, 0.000119035048677428, 0.000224098188684411, 
    0.000168282144706671, 0.000124045548473527, 3.84230775311378e-05, 
    4.73227944569276e-06, 4.0093538935517e-07, 2.34054341909817e-08, 
    2.11129718368337e-05, 3.24370046861511e-05, 6.13793493617198e-05, 
    0.000144736805816828, 0.000149848030689661, 1.27720447807778e-05, 
    0.000146007203901572, 0.000204393709098037, 0.000206367860537508, 
    1.78689746616036e-05, 2.01517595287957e-05, 0.000206235579939827, 
    9.33882055115585e-06, 0.000137404271345174, 0.0001220352357803, 
    9.65639291594207e-05, 7.93304313326017e-05, 3.65606500472654e-05, 
    4.86855411147485e-05, 0.000188611807798979, 0.000220135142799285, 
    0.000244479224964973, 0.000124188903245433, 0.000214725778612546, 
    0.000160931529976461, 1.09044704966072e-05, 8.64861664340564e-09,
  2.53053028046036e-07, 3.22885408871116e-05, 8.95786801685723e-05, 
    0.000210337544613297, 0.000209848231924786, 3.11107060784295e-05, 
    0.000207809052740722, 0.00017357138689245, 1.30851505002113e-05, 
    0.000115594946325787, 3.93687416522891e-05, 3.54064492442724e-05, 
    1.99962749353174e-05, 1.75049602595526e-05, 2.78874545391142e-09, 
    3.04971076036575e-07, 1.70733498188112e-16, 2.71248156924622e-16, 0, 0, 
    0, 2.18027131350444e-08, 1.22337965567207e-07, 4.38075945759037e-05, 
    9.54055564959509e-05, 0.000138369764724334, 0.000177119155074143, 
    0.00020604140114075, 0.000200640124839666, 0.000229409166156283, 
    0.000218734345155912, 8.40679614621601e-05, 2.35574813454933e-05, 
    0.000327818771712642, 0.000297121933068278, 0.000324560900272522, 
    0.000317232408332432, 0.000308588724166096, 0.000201524970534042, 
    3.64341521957896e-05, 5.1579509837894e-05, 0.000158581421176543, 
    0.000121528609145263, 0.000143770793527214, 7.29423534313766e-05, 
    5.72875116485101e-05, 6.72481109041144e-05, 0.000195027527885448, 
    0.000230919753135652, 0.00016628716236319, 3.27862999455703e-05, 
    5.15116081626955e-05, 6.03050070848376e-05, 7.48032950988022e-05, 
    5.50926315879507e-05, 4.75459728356565e-05, 4.47455818386678e-05, 
    7.15470099991713e-05, 8.44084114808268e-05, 2.27516126126267e-05, 
    0.000100465462830706, 0.0001540191693853, 0.00026936448234142, 
    0.00023564868627479, 2.13075312224391e-05, 8.04774884716507e-07, 
    9.44466897655919e-07, 3.44278915151518e-05, 9.35817263067536e-05, 
    8.60580784034212e-05, 5.53673970690062e-05, 9.66248360990587e-05, 
    1.31416949894309e-05, 8.68343542214446e-06, 1.80053398654841e-05, 
    1.88077844382704e-05, 2.87520658682601e-05, 2.78808598800361e-05, 
    1.46947875309258e-05, 1.87862346483172e-05, 2.06456522558645e-05, 
    1.58776017892843e-05, 1.46666507995176e-05, 1.94874639236862e-05, 
    3.67546040399341e-05, 5.83570455850062e-05, 9.71699254392666e-05, 
    0.000104569342059108, 0.000125147042249084, 0.000140215729170864, 
    0.000161283403982898, 0.000195011131899013, 0.000172321590120124, 
    3.62145323426433e-05, 2.37475724088942e-05, 4.77364669972485e-05, 
    8.076488599425e-05, 0.000102415617108309, 0.000131577558041649, 
    3.40192457667173e-05, 6.29462817950281e-05, 0.000187388285273583, 
    5.37206105711642e-05, 4.80522222320682e-05, 5.73400074198052e-05, 
    4.58528129549312e-05, 6.66391119038089e-06, 5.26257722163429e-06, 
    7.05962866803873e-05, 0.000102519436823915, 8.34211032173832e-05, 
    3.80064663579314e-05, 3.94068312437784e-05, 3.14316273040938e-05, 
    1.66135932888677e-05, 2.50051741309801e-05, 7.94072091953883e-06, 
    6.67747348536361e-06, 3.85793001827126e-05, 4.32707000484373e-05, 
    6.64570011843135e-05, 9.50119250729865e-05, 3.0864979121898e-05, 
    2.83625564579315e-05, 1.96493420894851e-05, 2.01050514846593e-05, 
    1.8060879815883e-05, 1.84401046445813e-05, 1.84889398942742e-05, 
    2.11168915025853e-05, 1.81423899384103e-05, 9.97510667528648e-06, 
    1.31982466168771e-05, 9.69732042755302e-06, 4.79439311686969e-08, 
    2.35616389765484e-05, 0.000154199776281069, 6.28768491219755e-05, 
    5.78401247983525e-05, 0.000101634462623086, 0.000187476287223506, 
    8.86855859640618e-05, 8.58082738372502e-05, 2.11732292405371e-09,
  8.01131587071351e-05, 5.13231834980034e-05, 0.000141468833712639, 
    0.000194331075585472, 0.000154555864742948, 0.000268330053370444, 
    0.000230455046084229, 0.000177809358568029, 1.57405552359066e-05, 
    7.16806221769806e-05, 0, 0, 0, 4.16891137954021e-07, 
    6.51011533661655e-06, 1.10735311505432e-08, 1.32557975713398e-16, 0, 0, 
    0, 0, 1.23579827685888e-08, 4.34564705693565e-06, 1.08445369547997e-05, 
    7.43924179689289e-05, 0.000102350066326332, 9.73742117500366e-05, 
    0.000119623878089288, 0.00015815358824489, 0.00020202666710415, 
    0.000154495082911941, 4.49643420563871e-06, 3.49437364692314e-05, 
    0.000261840194611199, 0.000294000633458626, 0.000300906429965174, 
    0.000226764436796148, 0.000174423786785992, 0.000180916181260192, 
    2.31514649169734e-05, 7.22549290321509e-05, 0.000110764848612343, 
    0.000117824138717793, 0.000109959486240444, 1.45203432273624e-05, 
    2.05801331369516e-11, 4.73297234550559e-06, 5.42283180926596e-05, 
    9.43138115846576e-05, 0.000354299220099786, 0.000156238888437667, 
    4.18430954496126e-05, 3.79388157592895e-05, 5.4846033651071e-05, 
    3.44724387667412e-05, 4.47519380882963e-05, 7.11913508657264e-05, 
    0.000192111847510233, 0.000111627257539278, 0.000122536676611762, 
    0.000164617688491446, 0.000299506679253642, 0.000222894446813503, 
    0.000222644746856015, 0.000156481662324825, 9.11209145932713e-06, 
    2.2470812779739e-05, 0.000162375871914152, 0.000201335548771845, 
    7.58544466728162e-05, 6.82815543450809e-05, 3.23831251377185e-05, 
    9.98607629754067e-06, 8.09895538808965e-06, 6.40703100526928e-06, 
    5.36837833939942e-06, 6.69132750217241e-06, 1.59788183089344e-05, 
    2.60147617924628e-06, 5.74833276351283e-06, 8.67727592380099e-06, 
    1.13120668166741e-05, 1.13867680285856e-05, 7.61831979517613e-06, 
    1.27479498717253e-05, 3.28794389328271e-05, 2.95565031385522e-05, 
    3.36252098549299e-05, 8.75819724823141e-06, 5.84541237022604e-06, 
    1.17903854656721e-05, 1.0724901127054e-05, 1.03995853997244e-05, 
    1.979217547639e-06, 1.43439631527492e-06, 7.11211105659496e-06, 
    5.21830703075359e-06, 6.19268657457218e-06, 4.61101522101032e-06, 
    6.84254840468369e-07, 2.5568329479683e-05, 0.000137140445113795, 
    2.60033787033404e-05, 3.81757349128348e-05, 0.000206217155460039, 
    0.00018413161077858, 0.000107507219606397, 0.000145232326854031, 
    0.000167983973763823, 0.000116623048236012, 2.96898710921182e-05, 
    5.64529318392293e-05, 4.93144628128209e-05, 3.34986394788996e-05, 
    4.10321453921526e-05, 8.81360913952418e-05, 7.84013360643909e-06, 
    1.18717761281857e-05, 1.43693726186778e-05, 1.24861215159532e-05, 
    1.56566551987777e-05, 1.57542943386323e-05, 1.24827401581427e-05, 
    2.08983481516375e-05, 2.17898839208673e-05, 1.71267805987478e-05, 
    7.5258107887823e-06, 1.3892153821934e-05, 1.17680599885141e-05, 
    1.16513393778645e-05, 9.49129997620071e-06, 7.02639867564115e-06, 
    5.92951964040632e-06, 5.98797149268334e-06, 2.70897126441594e-06, 
    1.63535655414057e-06, 1.45544836691742e-06, 2.97214198656233e-10, 
    1.6283028754715e-05, 4.22568272788584e-05, 0.000170163525075184, 
    2.54236147857681e-05, 7.62797715738214e-05, 7.17896454706447e-05,
  2.95549841906432e-05, 6.49525642770465e-06, 4.0018576181508e-05, 
    2.10185538391949e-05, 1.03839166246117e-05, 4.40468665917397e-05, 
    6.34790667337333e-05, 8.87787325809415e-05, 7.39732957198183e-05, 
    2.53532574140231e-18, 0, 0, 0, 0, 5.95349195106316e-13, 
    3.64083517227082e-14, 0, 7.18304137948667e-16, 0, 4.74330451821151e-20, 
    4.90957512730329e-20, 1.31538271457497e-10, 6.00404789013489e-07, 
    1.86005538955416e-05, 4.70426035569721e-05, 0.000105943046358797, 
    0.000116147512275435, 0.000112124070290414, 0.000174618590045405, 
    0.000158091054639449, 9.30200239504452e-05, 9.61954331369594e-06, 
    2.01985841307947e-09, 0.00015242765567965, 0.000182245669997514, 
    0.000187218697580624, 0.000147600412698148, 9.40679274012537e-05, 
    8.81191350568898e-05, 2.36809400984274e-05, 6.65267496123988e-05, 
    0.000113856983829457, 5.90089441662074e-05, 7.97660039072733e-06, 
    7.90505139538367e-06, 5.60123018050206e-11, 8.28765811652158e-06, 
    1.24862965125986e-05, 4.46713202731228e-05, 0.00095425820197036, 
    0.00073086033417592, 0.000224578693931433, 2.94021693310788e-05, 
    3.73063267996905e-05, 4.84580821018747e-05, 7.57400903661231e-05, 
    0.000206436967347634, 0.000270194963921947, 0.000293499256396186, 
    0.000264661643155523, 0.000263513808359944, 0.000230859778190849, 
    0.000119889437392483, 0.000123211282943787, 0.00016047967285756, 
    3.83480255333083e-05, 0.000108658101628606, 0.000183993859627598, 
    0.000188607243193337, 9.60054437489072e-05, 4.4165747175614e-05, 
    2.52729251592504e-05, 2.19618077295365e-05, 1.12967022925732e-05, 
    4.81536431908898e-06, 1.10100686817051e-05, 6.30977331767377e-06, 
    1.03116580831568e-05, 9.2160392048696e-06, 5.08150198035668e-06, 
    5.69020997835171e-06, 7.95461956300217e-06, 9.0121514248352e-06, 
    8.56087279377581e-06, 5.91689136180899e-06, 6.51619281366058e-06, 
    5.97050581985944e-06, 1.67470368978483e-06, 2.20378572163826e-06, 
    1.59427225715681e-06, 1.69739517610065e-07, 5.56566073925949e-07, 
    1.35941589547514e-06, 6.01059061405652e-07, 1.29920025872254e-16, 
    1.65262146732982e-09, 4.8663634759315e-09, 4.6463779304177e-19, 0, 0, 0, 
    9.99927532006579e-05, 0.000267595048799859, 0.000378839663380921, 
    0.000289667192561614, 0.000218066158942188, 0.00020413101928752, 
    0.000191963708859321, 0.000164225937856238, 7.35797577058252e-05, 
    1.29319867591958e-05, 8.50611570774235e-06, 3.12352495338715e-05, 
    9.27279883309428e-05, 7.99456073552901e-05, 1.34606259050946e-05, 
    1.62641755992498e-05, 1.92148387010564e-05, 1.1650561332966e-05, 
    4.62366629014919e-06, 1.16269127920482e-05, 1.15101494019585e-05, 
    1.84688090461477e-05, 1.50190536260123e-05, 1.44230422108536e-05, 
    1.55419809844541e-05, 1.48339038415649e-05, 1.62544063038134e-05, 
    8.65983981967745e-06, 5.28946640756748e-06, 1.09370614820084e-05, 
    6.48583449519396e-06, 1.1770206205633e-05, 2.52729158859504e-06, 
    4.02993105066171e-06, 5.87944128068684e-06, 3.82355291135293e-07, 
    7.14495542544456e-11, 4.12856521517419e-10, 3.36922882939505e-11, 
    5.9625174731877e-06, 2.13437988500446e-16, 3.13165306647102e-23, 
    9.47433053764863e-05,
  1.27905043772616e-07, 0, 2.55163882048501e-07, 0, 7.80229379520163e-07, 
    1.74638410578605e-18, 1.95589183551199e-17, 1.72510103748733e-05, 
    8.34948323995908e-17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.63133028087999e-18, 0, 
    6.27771581855819e-18, 4.1666815041257e-14, 5.20743771870917e-07, 
    3.42382512217338e-06, 2.95043729621904e-05, 3.24417477724744e-05, 
    7.09512478254623e-05, 8.49121727937204e-05, 0.000132371990147246, 
    0.000121390546536581, 4.85309668788913e-05, 8.45965463539506e-05, 
    0.000105204989873059, 9.58506946685214e-05, 0.000140137829403644, 
    0.000136836271765194, 0.000109118383634136, 7.61151018057562e-05, 
    5.04710610230801e-05, 5.42037850707997e-05, 7.97291576472552e-05, 
    4.83607609578352e-05, 1.40143039119245e-06, 1.58929835467198e-05, 
    1.93855319913973e-05, 2.39073326866134e-05, 2.11928701926118e-05, 
    2.37643560158218e-05, 3.08082058255804e-05, 0.000140786780442301, 
    0.000743274289375022, 0.000343645771790625, 7.78944772981233e-05, 
    6.44434288301469e-05, 0.000132745035681298, 0.000168662803025729, 
    0.000282619497853491, 0.000325023636171622, 0.000333170646699752, 
    0.000305823595572329, 0.000213052628482386, 2.54644844101396e-05, 
    6.49191109689884e-06, 7.49711917659255e-05, 0.000156321020317867, 
    9.34849677467911e-05, 0.000149632446827677, 0.000156051853204407, 
    0.000159609012161181, 0.000117463309801052, 9.24302036693217e-05, 
    5.90027957621278e-05, 1.7915078392562e-05, 1.6946913808025e-05, 
    1.39293874879597e-05, 5.2318404098393e-06, 5.364755228961e-06, 
    2.05501909000806e-06, 8.29849159552452e-06, 3.33617214631694e-06, 
    2.74730551432949e-06, 4.89861071869235e-06, 2.82860934671454e-06, 
    6.29161234793229e-07, 1.60837533775517e-06, 2.04303849283921e-06, 
    1.55858244679142e-06, 2.39242652515582e-06, 4.94517838874808e-06, 
    4.08485338791058e-07, 4.32850927684473e-09, 8.30763963976762e-11, 
    2.53446521463615e-11, 1.45266249014478e-13, 0, 0, 0, 0, 0, 0, 
    2.05495164862669e-19, 5.59662274758572e-05, 6.94033570601726e-05, 
    0.000341317775008752, 0.000145203996540816, 0.000198719750590641, 
    7.86436673651251e-05, 4.55930573529605e-05, 1.6483264446616e-05, 
    4.93041748146395e-06, 1.02137657987946e-05, 0, 3.0429947952388e-23, 0, 
    1.76911343414833e-19, 3.20598906173403e-07, 7.66344562108967e-06, 
    5.70666969211064e-06, 5.42219889116184e-06, 6.11027555519382e-06, 
    9.85015480870629e-06, 1.24919217660131e-05, 1.20631888586026e-05, 
    1.04170098087548e-05, 1.29038685731743e-05, 1.02228185410827e-05, 
    1.21316443841143e-05, 9.40796273462988e-06, 9.87108236863351e-06, 
    3.17478312365334e-06, 9.00878494737073e-06, 1.01594903977334e-05, 
    4.47582033586745e-06, 5.57431093665882e-06, 2.6240257763869e-06, 
    3.98513256988498e-06, 3.0420076044807e-07, 0, 4.59844627555815e-12, 
    2.69916508696005e-22, 7.26007903270669e-05, 5.47608579662335e-05, 
    1.29951674319182e-22, 6.75927161980427e-06,
  0, 2.24069970089125e-05, 0, 3.8388526936501e-22, 7.73996001734294e-25, 
    8.19335693018415e-23, 1.66576143362809e-18, 9.48917014926926e-11, 
    1.59852363001935e-17, 0, 0, 0, 0, 0, 9.04983333963993e-19, 0, 0, 0, 0, 0, 
    0, 0, 2.842199899013e-11, 1.95936398335845e-07, 2.87168882498384e-06, 
    2.61133602048514e-05, 3.2608422904817e-05, 5.08299936511459e-05, 
    3.07408169053914e-05, 2.43874738597379e-05, 1.93691707808272e-05, 
    6.64085446708066e-05, 0.000155075770502116, 0.00018675732368063, 
    0.000132202045662551, 5.47306914973032e-05, 8.07514763008281e-05, 
    1.50973133268545e-05, 2.87982490198551e-05, 6.08778896294333e-05, 
    6.8892967220592e-05, 1.19543872205755e-05, 1.26709986281256e-05, 
    2.45024050167081e-06, 2.40573180332692e-06, 4.19880011031165e-06, 
    1.70836341909653e-05, 1.95925669536409e-05, 4.11503546994535e-09, 
    6.72060776081852e-06, 6.06201864750102e-05, 7.92793235318021e-05, 
    0.000127452926772691, 0.00021864539511477, 0.000272050547501842, 
    0.000266150313979403, 0.000245577261134314, 0.00031324704448569, 
    0.00039626775641735, 0.000272437446022782, 0.000229787165961605, 
    9.28044788289031e-05, 8.676842908697e-05, 0.000122353993700348, 
    0.000193756591610452, 0.000200300316470102, 0.000229795276948015, 
    0.000252316466193538, 0.000278295888445373, 0.000271214269504928, 
    0.000161694733530409, 0.000102571611535881, 4.39617610367251e-05, 
    3.71129650327113e-05, 2.31674731365469e-05, 3.66030838116618e-06, 
    1.38569406176611e-09, 4.24477620341798e-07, 3.86411899614703e-06, 0, 
    2.29395986964966e-06, 6.10844472805875e-06, 2.62855404392703e-06, 
    6.07358999230211e-07, 1.53759173671032e-06, 1.61112770363319e-08, 
    7.13777950549999e-07, 2.73869809264178e-06, 2.30049046609418e-06, 
    1.45277785612526e-06, 1.97544140011781e-06, 5.05707413861977e-08, 
    1.51136182919504e-11, 2.86717434475503e-10, 2.96077663747976e-20, 0, 0, 
    0, 0, 1.25158669643235e-21, 3.95848060118655e-18, 1.32409807132327e-09, 
    0.000142182602676737, 0.000100216675063312, 0.000215710906276431, 
    0.000180556744099257, 1.69893185719719e-05, 4.4912118658453e-07, 
    1.85716382438767e-09, 3.15730665899809e-06, 5.07133400202955e-06, 
    7.8562721602251e-61, 3.60303908189531e-18, 0, 5.70920638026858e-06, 
    9.85484054013624e-06, 6.66521113403321e-06, 9.59678541890641e-06, 
    9.57598490882126e-06, 7.47587573858608e-06, 6.26622579042598e-06, 
    7.88003447042891e-06, 1.13388034568153e-05, 1.07480732866269e-05, 
    8.99797596123155e-06, 9.01371738163352e-06, 8.93988433953757e-06, 
    1.36924544322275e-05, 1.26284923472512e-05, 9.98623409335745e-06, 
    1.06014064273522e-05, 5.66243479549325e-06, 4.2213718154079e-06, 
    3.01121641086025e-06, 1.58572037575514e-06, 2.58011609720282e-08, 
    6.25059931997231e-07, 0, 6.57369383233631e-16, 0, 6.83038910890255e-18, 
    8.08510431880813e-05, 1.6966270843347e-18, 3.36570401504066e-19,
  0, 4.19171375116666e-06, 0, 3.28707490271351e-22, 3.15038470654746e-18, 
    9.16007174491219e-20, 4.44788160586765e-08, 1.18325471509848e-17, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.55350949136854e-17, 2.77304201735211e-18, 
    1.36254766738279e-17, 2.1713149897424e-10, 6.53316820854757e-07, 
    9.98719225140015e-06, 1.8637181947948e-05, 8.04240355777446e-06, 
    2.3116597258646e-06, 6.95337204874397e-06, 1.81328835906495e-05, 
    2.50929807024218e-05, 6.6761733048133e-05, 0.000207265467139942, 
    6.00167530486143e-05, 5.50540739656793e-09, 6.84839932158789e-08, 
    3.99065666108814e-05, 2.55644684332389e-05, 7.09473663939956e-05, 
    6.85672830090586e-05, 3.37113090653317e-05, 1.81406556030885e-05, 
    1.22161252352162e-06, 1.29513671910669e-06, 8.42373769087355e-07, 
    6.95330992416767e-25, 4.11080252566967e-08, 6.34460625721182e-10, 
    9.04538179256536e-06, 1.84240301251795e-05, 4.52638009615388e-05, 
    9.68869773011134e-05, 6.22648450642718e-05, 0.000152157566679531, 
    0.000208461023222541, 0.000265491942417667, 0.000266457653149487, 
    0.000316696753717572, 0.000305824480282733, 0.000213942459836084, 
    0.000192649327472145, 0.000183890709787333, 0.000181077838610341, 
    0.000299282489263625, 0.000307994361354778, 0.000374590704919585, 
    0.000355576142499309, 0.000391990646475597, 0.00038382061359734, 
    0.000184729631477416, 7.51357728965668e-05, 0.000125622834176046, 
    0.000151593657666956, 9.69615342558057e-05, 6.5134414240846e-05, 
    5.89094234382945e-05, 3.1668238319179e-05, 4.87891158708208e-05, 
    6.61624613201678e-05, 6.04174625369088e-06, 4.60151892420456e-06, 
    2.85430584442207e-06, 3.00011347539689e-08, 4.71417695081143e-07, 
    7.32532035555696e-07, 1.68253961712921e-06, 1.06682954284835e-06, 
    2.07514423471758e-06, 1.68438715284059e-06, 1.45995004769362e-06, 
    9.70778574668195e-07, 4.44414304207413e-09, 3.91495930858121e-08, 
    1.56369694482685e-09, 0, 1.32230651508894e-08, 0, 0, 3.5603754268507e-20, 
    3.93343864750855e-19, 2.4419443384848e-10, 0.000384694094073909, 
    0.000136620027889565, 0.000174150293400246, 0.000129488389675489, 
    2.73590183616852e-07, 9.4942902493553e-06, 8.75728452273196e-06, 
    1.98769821174949e-08, 1.81187341026282e-10, 0, 4.67042624375091e-11, 
    1.34352388092637e-07, 2.06207811399445e-07, 1.03552819908347e-05, 
    8.57710691804347e-06, 1.02636393049487e-05, 8.4728705412661e-06, 
    5.97926929873473e-06, 4.61162990429822e-06, 4.75200592195134e-06, 
    5.78237970673261e-06, 8.39172042381243e-06, 9.21045405905039e-06, 
    9.48081634480178e-06, 1.03151184323585e-05, 1.15170584458057e-05, 
    1.24103014951624e-05, 1.46582607585574e-05, 1.29421417691039e-05, 
    6.64827437388442e-06, 4.41590922684405e-06, 8.77241401529098e-06, 
    3.53816024125994e-06, 4.28233442741607e-07, 1.2649674205868e-06, 
    2.15039845138658e-07, 0, 2.55809098363952e-17, 0, 0, 
    4.41633944756383e-06, 0,
  3.39485886390867e-05, 0, 1.28775932446842e-23, 2.04870523784926e-23, 
    7.94417364463339e-47, 1.72059144816486e-17, 0, 1.65441514242275e-10, 
    6.88826715344026e-21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.24662316519571e-21, 
    0, 0, 4.5238247248605e-14, 9.58916845912524e-10, 9.46726072616563e-07, 
    6.34885895778665e-06, 4.06524574370355e-06, 2.08046747603421e-06, 
    1.75761583003959e-06, 5.48285303154191e-07, 1.79504388780386e-06, 
    1.23773154524316e-07, 0.000149446517351314, 0.000192876954056706, 
    0.000104965029552338, 1.92404443955657e-05, 1.43224657467338e-07, 
    5.5640799035461e-05, 4.98172205188308e-05, 6.62720416286099e-05, 
    7.93674420119177e-05, 5.15712256835532e-05, 1.83566266440484e-05, 
    1.021737541445e-05, 1.99592769324254e-06, 5.13030912759636e-07, 
    8.78087878402716e-09, 2.51007442128592e-06, 1.65852176895573e-05, 
    1.93038257776917e-05, 3.561582255154e-05, 1.94874474953184e-05, 
    1.66768319155148e-05, 1.55756538528699e-06, 7.67710506106003e-05, 
    0.000263089676026007, 0.000245245604792484, 0.000310740991880011, 
    0.000358358108934927, 0.000162136038274604, 0.000136607005424404, 
    0.000192286642752996, 0.000268192242758683, 0.000429757516932853, 
    0.000463435748149267, 0.000331736156921084, 0.00019857369149133, 
    0.000178147970715704, 0.000230025066639987, 0.000210594855517481, 
    2.06463327252009e-05, 1.12137600046666e-06, 7.98959410929038e-06, 
    5.11611579128381e-05, 4.66500034906596e-05, 1.43128420832087e-05, 
    1.26785843132736e-05, 3.50617808384465e-05, 0.000108913509926949, 
    1.1374528846544e-05, 8.32209599156897e-06, 4.55332593292175e-06, 
    2.24701177418013e-06, 5.233438611302e-10, 5.27272163478947e-07, 
    1.89626422357824e-07, 1.16943824834265e-06, 4.62242568122582e-07, 
    1.04087291218488e-07, 7.49276700422865e-07, 6.65423049636059e-07, 
    1.37164513308032e-06, 1.50024603344538e-06, 3.57704842593739e-07, 
    5.03799435518551e-08, 0, 0, 1.82806604256639e-08, 0, 0, 
    1.50765370640294e-16, 1.67690995661803e-16, 2.18209084693406e-05, 
    0.000154140296450308, 7.35823557672648e-05, 8.98919651239328e-05, 
    5.11602495621017e-06, 0, 0, 5.89049901234382e-06, 1.33230176071846e-06, 
    8.67159205560758e-07, 3.92625599348894e-07, 5.50481394326833e-11, 
    1.19158299812405e-06, 4.61105103021793e-06, 6.70794918690224e-06, 
    6.18926661477498e-06, 5.34804203381652e-06, 3.54041485310003e-06, 
    3.443838035014e-06, 2.89357722175458e-06, 3.32010768803854e-06, 
    3.93838104289832e-06, 4.10758807925202e-06, 5.15975057475697e-06, 
    6.62194886511929e-06, 8.26825821028247e-06, 1.60761508052352e-05, 
    1.59570292439275e-05, 1.48571903183364e-05, 6.47692743367237e-06, 
    8.0938329448747e-07, 3.91237583610421e-06, 1.25223581194319e-06, 
    5.69031904200241e-07, 1.98615795827448e-06, 7.35609806883823e-07, 0, 0, 
    0, 2.60108999484238e-17, 4.21727408845312e-06, 1.65002758756029e-24,
  0, 0, 0, 6.09402470816819e-20, 0, 1.09249656867234e-22, 
    9.01589030488684e-21, 8.86888086809125e-19, 1.50093055167006e-19, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2.03206843724196e-14, 0, 2.69939037314597e-20, 
    4.42597445715406e-11, 8.45514271333577e-08, 8.23563029343733e-08, 
    9.2436210823674e-08, 4.51982938491634e-07, 9.59193671556389e-08, 
    4.95058411173305e-08, 1.97728743882867e-10, 6.44089889271357e-05, 
    8.95032544472006e-05, 0.000459960885690628, 0.000806459608044716, 
    0.000328199436113291, 4.24286224402737e-05, 7.09252509107555e-05, 
    5.0288596942721e-05, 3.33394454527421e-05, 3.89679930344029e-05, 
    4.43228372363929e-05, 2.53517685627511e-05, 1.32811608304961e-05, 
    4.24888964471529e-06, 1.34065454265415e-05, 6.47227940698562e-06, 
    1.57329790644377e-05, 2.02890885397763e-05, 5.16313892745332e-05, 
    8.93374164593336e-05, 4.048595979971e-05, 2.29912328282598e-05, 
    2.41264624217975e-05, 0.000233305914026446, 0.000216967770402956, 
    0.0002472920097786, 0.000170820356231889, 9.85095267404746e-05, 
    0.000150432083049533, 6.82766972465945e-05, 0.000160898882036928, 
    0.000220869792865529, 0.000314985602118068, 0.00016920542097697, 
    0.000128999373707545, 4.0261074654468e-05, 1.84370754638912e-05, 
    4.63253019595204e-06, 3.85137589326503e-05, 9.98919477685196e-06, 
    2.57391575360952e-23, 3.59828502333306e-05, 7.25888992165958e-05, 
    2.03241296311063e-10, 2.49549464755488e-06, 1.02338843302762e-05, 
    2.43055914524422e-05, 0.000104967880038697, 0.000132766036384787, 
    4.91925582246166e-06, 4.46809154521338e-06, 3.79982113045179e-08, 
    5.3696389777838e-07, 1.88958431802623e-07, 1.40203457698593e-07, 
    1.19521219083474e-06, 1.50733965769829e-10, 2.4241781369174e-07, 
    7.70283704947762e-08, 1.01137953033057e-06, 3.97413765291187e-07, 
    5.95457620068795e-07, 1.87873364554155e-06, 9.55990549400882e-07, 
    5.89957448786368e-11, 0, 0, 0, 1.74857686808956e-11, 
    9.29801520976114e-11, 7.01932568665524e-09, 3.0547518480932e-07, 
    1.75486904284583e-06, 2.6541486835135e-05, 5.09015517935266e-05, 
    1.32783153031187e-05, 4.58364459239221e-07, 0, 0, 0, 
    1.47066805998937e-06, 1.18524006144277e-05, 1.46996008602238e-07, 
    1.85702590523891e-06, 2.44106475459202e-06, 3.02880319866385e-06, 
    2.81509203551336e-06, 3.15662151116435e-06, 1.07949873030002e-06, 
    2.63342621784306e-06, 2.26324961945921e-06, 1.37237319805427e-06, 
    1.90099408559008e-06, 1.96092541602132e-06, 1.7494829628543e-06, 
    1.97119484142944e-06, 3.97995197288296e-06, 1.62763240179863e-05, 
    9.51984195801972e-06, 1.07843789390993e-05, 4.9062270328806e-06, 
    5.97512663387769e-06, 3.4283536948118e-06, 2.82208456003225e-06, 
    1.68443995593072e-07, 8.22578132368631e-07, 4.39272017811647e-07, 0, 0, 
    1.20461478079437e-16, 7.34696926012983e-08, 8.52253835658616e-05, 
    7.87327930853012e-06,
  1.61694228349081e-16, 1.44755186393873e-25, 1.24565595505605e-23, 0, 
    2.40322015943668e-11, 1.60357075765584e-17, 2.54933991827617e-21, 
    1.13192957255233e-16, 0, 2.75760450091192e-23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 8.27558927584115e-13, 0, 0, 3.78653234506084e-29, 
    1.96386192754542e-14, 4.93196856184289e-15, 3.3097558061641e-13, 
    1.32679844500898e-08, 6.51380771417536e-09, 4.27583576579255e-11, 
    6.16554621951034e-05, 0.00036865875398512, 0.000332814102217215, 
    0.000414423460412392, 0.000327064478894382, 1.15952159206123e-05, 
    1.6591615362711e-06, 3.36457566860231e-05, 3.2574788984308e-05, 
    4.77286024261011e-05, 6.42165938980796e-05, 3.05045518133851e-05, 
    1.30475527406147e-05, 5.13944754715787e-06, 1.30742505843129e-05, 
    3.87998879636223e-06, 1.20190597817615e-05, 9.16711384682632e-06, 
    5.06596237827254e-06, 0.000760367964280645, 0.0018331844376075, 
    0.00115149195900938, 0.000156840134623697, 0.000146116085255217, 
    0.000176534166762296, 9.83988272030757e-05, 0.000203052810034877, 
    4.68768617284717e-05, 3.52904134612033e-05, 9.91163757230049e-05, 
    0.000139937359524378, 0.000180903776613593, 0.000182820161685992, 
    7.47625513005609e-05, 3.87133673500129e-05, 6.44299260853805e-06, 
    3.88497587866836e-05, 1.7797399014308e-05, 1.62256328644712e-05, 
    5.9292916518858e-05, 4.61297544606232e-05, 0.00013967594399775, 
    7.34633304781573e-05, 4.57754534807354e-06, 1.34485148384186e-05, 
    1.2194442669612e-06, 8.22384393370996e-06, 4.1042285833239e-05, 
    7.32818006785166e-09, 6.77013498885557e-05, 3.79758505733438e-06, 
    6.34917184640908e-07, 5.74880395844885e-07, 2.35725408416111e-06, 
    1.42452267775985e-06, 1.08364367705265e-06, 2.91920991317799e-08, 
    4.93189380117982e-07, 8.88726610492286e-07, 1.02231584960574e-06, 
    9.01213190599141e-07, 1.52818121936879e-06, 5.03990612204486e-06, 
    3.90792292862421e-07, 1.9246310852772e-08, 4.43849822579529e-08, 0, 0, 
    2.93888693518645e-16, 1.40632521716668e-06, 2.06193501378179e-08, 
    7.96208220871047e-09, 8.63338061977949e-20, 1.73894765972268e-09, 
    1.18479839666617e-09, 0, 0, 4.9390138296285e-10, 3.97020881134079e-10, 
    4.58428221515864e-08, 0.00010785812932456, 6.88421678883749e-05, 
    3.45330808530499e-05, 5.16578740034408e-10, 2.57985732817534e-06, 
    3.92784214433047e-06, 2.52370432181738e-06, 3.58613451948651e-06, 
    3.84464515457156e-06, 5.6555693155766e-06, 7.15165777153532e-06, 
    5.54821854959429e-06, 5.08947294387836e-06, 1.92771561744436e-06, 
    8.77864854668396e-07, 2.43346778840241e-06, 2.74651435036285e-07, 
    1.35466092921618e-10, 1.44577382204038e-06, 6.24536902630369e-06, 
    5.6099851036317e-06, 4.70479835211861e-06, 3.25281195262475e-06, 
    2.46960192049194e-06, 2.04218581980116e-06, 7.27837317792775e-07, 
    1.87880995889729e-09, 0, 0, 5.72620955780369e-18, 6.50004741348751e-09, 
    0.000111200362097114, 3.87804890638245e-12,
  2.97996087079745e-06, 5.69978395535013e-07, 7.59645345011318e-18, 
    9.00809715689179e-11, 4.33745393257043e-11, 0, 4.12080859884674e-19, 0, 
    4.90475286111901e-19, 3.2273114035836e-18, 8.20460776039536e-24, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1.61408357233294e-10, 4.38147379526152e-13, 0, 0, 0, 
    0, 0, 1.37997357239641e-18, 8.97272563233676e-11, 0.000107355915311424, 
    7.20089179320338e-08, 2.64195539030124e-10, 1.89252271339156e-07, 
    3.62023328797658e-07, 1.01209645015673e-05, 1.40419168628179e-05, 
    1.1419274593226e-06, 1.12899116573313e-09, 2.54700629991108e-05, 
    4.07909178972735e-05, 8.8100514845181e-05, 7.03922865528926e-06, 
    2.89370222332383e-06, 3.91180100151229e-06, 7.92697412656637e-11, 
    2.04075723769606e-07, 1.74919685129525e-05, 4.174784745049e-06, 
    4.28851623600791e-11, 0.000436703822890965, 0.00182003533023195, 
    0.00162629627684789, 0.000243007873967389, 8.79996087929173e-05, 
    0.000109319915126416, 1.66174696803027e-05, 1.08010818155809e-05, 
    6.08920578984047e-06, 1.62930472201761e-05, 7.5036582572141e-05, 
    3.12023778664207e-05, 7.20226665584101e-05, 9.83275758686165e-05, 
    2.36079339582123e-05, 1.45299348755978e-05, 8.77061818697058e-06, 
    4.8697951349555e-06, 3.39714668641411e-06, 4.18171546865586e-18, 
    4.58313578041889e-05, 2.36705489890654e-05, 5.43515624227666e-10, 
    3.3159931427099e-06, 4.93636423055361e-06, 3.39875468629093e-06, 
    2.7806283881884e-06, 1.18857165431249e-10, 2.27783944580782e-06, 
    3.83583359287869e-06, 4.03881781733694e-06, 3.33534827278632e-08, 
    3.47782975585143e-06, 2.07442357814966e-06, 1.37274102912328e-06, 
    1.77361702770105e-06, 2.0304531324495e-08, 1.71961581820055e-06, 
    1.27484137076165e-06, 2.11780545800519e-06, 1.88834576665478e-06, 
    1.57236996213254e-06, 2.33161665708165e-06, 7.71995974019492e-07, 
    6.10723823131281e-07, 1.73707315907366e-07, 0, 0, 0, 0, 
    6.65198997888524e-10, 1.06356975111643e-05, 1.78768761491517e-10, 
    1.9021551012857e-24, 0, 2.24294666569317e-11, 1.23155711989322e-09, 
    5.59726576227203e-05, 2.88101730562256e-05, 1.18074395584102e-05, 
    1.97741485192316e-05, 0.000189591410380219, 0.000148042812759644, 
    0.000105098425655102, 0.000109112942662821, 7.05266137334514e-05, 
    1.0374962357268e-05, 4.38158343257986e-06, 7.70509468819309e-06, 
    7.60768390346685e-06, 1.32129913551622e-05, 3.98181171166701e-05, 
    4.57734079994361e-05, 2.01921142339587e-05, 9.0970360543416e-06, 
    6.37108451185157e-06, 9.37755991073721e-06, 7.88515280671945e-06, 
    9.1327691620314e-09, 4.523133598927e-10, 2.64415101109219e-06, 
    7.7969135649904e-06, 5.9374006259268e-06, 5.98015125650599e-06, 
    1.28814224713869e-06, 3.613281293655e-06, 2.43930841649397e-06, 
    5.65482095040565e-20, 0, 0, 0, 7.27834087303402e-09, 
    1.49627640477205e-05, 1.64312039134243e-05,
  9.51514870276153e-24, 4.31952796785191e-05, 3.06141924847325e-05, 
    1.69093646023878e-05, 4.19886593096696e-24, 2.40412666507425e-19, 0, 
    2.05162410455546e-19, 3.22403343952888e-17, 7.77969438756235e-23, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8.20520270766513e-21, 0, 0, 0, 0, 0, 0, 
    2.97060215971665e-18, 1.99289847777427e-12, 8.79091577148842e-18, 
    9.26587065637503e-09, 5.86129072075635e-10, 1.20613820732878e-07, 
    5.98892685388535e-09, 1.79110544118726e-07, 1.22997035948537e-08, 
    2.63834072733121e-06, 8.37197269548813e-05, 0.000121958198411081, 
    0.00010404250600897, 0.00015942612642242, 7.75033725390394e-06, 
    2.22848633325708e-09, 1.16878798670527e-09, 6.51928380518885e-11, 
    3.942984898888e-08, 2.32327847706204e-08, 4.09850208708097e-09, 
    4.30925098495424e-12, 3.11076386457865e-10, 2.39676727473497e-07, 
    1.15591769274481e-05, 7.17571720237882e-07, 8.65656885687254e-06, 
    4.12726078783947e-06, 1.83886756756563e-05, 1.97134592911307e-05, 
    8.22812186772522e-08, 1.02056466910411e-05, 1.57203754884812e-05, 
    2.13022059715484e-09, 9.17514195437086e-21, 8.38207194869157e-06, 
    1.64108539618738e-06, 4.2134909143658e-06, 3.85314917532984e-06, 
    2.04166403812976e-06, 2.80834853974081e-06, 3.64330958337498e-06, 
    3.70692660764788e-06, 3.82337321746529e-06, 1.49426727579883e-06, 
    3.65803176137101e-06, 3.13650898379707e-06, 2.28025696231735e-06, 
    8.36066651320971e-07, 4.03934827712251e-08, 6.64523575582103e-09, 
    4.64216501949502e-06, 1.66405648826762e-06, 2.2879464698073e-06, 
    7.95624808649095e-06, 5.28226265079496e-06, 4.50038474223566e-06, 
    2.07150550016734e-06, 7.10202694026119e-07, 6.96794252807388e-07, 
    1.41898356174509e-06, 1.7934070098091e-06, 5.49860642124874e-06, 
    6.48168014557245e-07, 7.60055639954159e-07, 1.19757192571981e-06, 
    7.05996613874357e-08, 3.31963769541845e-09, 0, 0, 0, 0, 
    4.04914099714734e-12, 2.23334957894518e-08, 2.04918591746689e-05, 
    4.32488731918906e-24, 0, 1.01054272172245e-09, 9.22920391337708e-08, 
    0.00010614124468899, 0.000182280253556949, 1.0036520710644e-05, 
    2.41777607372437e-06, 7.26710002800477e-09, 7.79760347333316e-05, 
    3.52836121289621e-05, 2.72032715650072e-05, 1.24752545444042e-05, 
    1.97387034510381e-05, 6.47856990343658e-05, 6.8467378250797e-05, 
    6.4108993104712e-05, 2.79134025990811e-05, 4.11081712756581e-05, 
    8.6130463581989e-05, 3.26821833773758e-05, 1.83069974337125e-06, 
    3.09562693525837e-07, 2.15104041443969e-06, 6.48737888914255e-06, 
    1.17604622203452e-20, 5.02917692946169e-06, 6.60740028009812e-06, 
    6.04520793778955e-06, 6.94154995108796e-06, 2.68992839242729e-06, 
    3.24654366559222e-06, 3.61354861535916e-06, 2.1482430113278e-06, 
    2.55944113401091e-10, 0, 0, 0, 4.86060452303258e-15, 
    8.57625268317347e-12, 5.53497391939874e-09,
  9.47451028327012e-09, 6.76777683130557e-05, 0.000142952884401433, 
    0.000105569084091738, 1.78196242285553e-06, 3.83752547254332e-19, 
    7.03622251240994e-18, 0, 0, 0, 0, 0, 0, 5.10185985763463e-25, 
    5.42191042134367e-23, 0, 0, 0, 0, 0, 0, 7.99768462313441e-19, 
    2.18170954512392e-20, 0, 0, 0, 0, 0, 0, 2.10778365423145e-12, 
    2.83505508377642e-12, 3.47146498215168e-19, 4.32348514099163e-11, 
    1.56825507802677e-10, 2.88342564731577e-10, 0, 6.18223833701406e-09, 
    5.7418091583808e-08, 1.13300143703178e-05, 0.000151449220941512, 
    0.000163894148500167, 0.000172901794891672, 0.000546068141000518, 
    0.000202613689524985, 9.5259865309915e-09, 4.21008596376926e-10, 
    1.06328728771745e-08, 5.2241518198566e-09, 2.17063538297247e-08, 
    7.63261646248202e-10, 7.82142812240365e-09, 9.47154031320813e-08, 
    1.42436782007945e-09, 1.34957359947923e-08, 1.78394481161902e-06, 
    6.38354806944518e-05, 2.87266956019094e-05, 1.48707819812038e-05, 
    7.8695183787606e-10, 1.03714459850807e-07, 4.99878242954237e-06, 
    1.12126864174023e-06, 1.92348229528941e-11, 9.45414262881299e-12, 
    2.02833154803381e-08, 4.89733370475472e-06, 1.31359590658049e-06, 
    1.34783079582954e-09, 1.84741479202023e-08, 2.74347978916107e-06, 
    6.12917219773e-09, 5.5943002632801e-06, 2.7484980091013e-06, 
    2.06155224666966e-06, 2.08918837394389e-06, 4.01378747213325e-07, 
    2.4627660937282e-09, 8.68315025729016e-07, 1.85233064148309e-06, 
    1.75776716538013e-07, 4.73932430553261e-07, 3.59600002328325e-05, 
    3.10798732921194e-07, 9.90586398464563e-06, 6.72615994388597e-06, 
    1.78659944426688e-06, 9.08872192919453e-07, 2.42127045011099e-06, 
    1.8190515679108e-06, 1.49533411172425e-06, 6.49248510995228e-06, 
    2.25809531332437e-06, 3.01031129861596e-06, 1.70706099783807e-06, 0, 0, 
    0, 0, 0, 7.49689039290272e-18, 3.05050625868016e-19, 
    8.76857435036567e-11, 2.46875017680938e-05, 2.01248592408131e-19, 
    1.000046798101e-11, 9.24647428493644e-06, 3.59144066418865e-08, 
    8.42595017616746e-05, 0.000113815075169294, 3.80774902051638e-11, 0, 
    3.53012089468888e-10, 0, 2.68542905092608e-10, 0, 0, 0, 
    4.08672113112159e-07, 6.28264598454855e-05, 6.00171880559447e-05, 
    4.28467344945761e-05, 2.26513131998717e-05, 2.10527021896666e-05, 
    7.43793350748537e-06, 7.37429498458119e-06, 3.49151299015781e-06, 
    2.9629748823548e-06, 4.1940153698626e-06, 1.25944144197441e-06, 
    1.27423340546625e-05, 4.15007654078174e-05, 3.63469888045191e-06, 
    3.96205400755086e-06, 2.0285753242305e-06, 1.51395160546731e-06, 
    2.99927185248771e-06, 1.09274692646157e-06, 9.23590494719016e-08, 0, 0, 
    0, 8.36235785877882e-24, 1.28674370747444e-16, 5.28141546964636e-12,
  4.51095259820253e-17, 1.32058030936694e-19, 8.15341977928283e-05, 
    0.000136889892996526, 3.74317539106112e-05, 1.2190785913445e-11, 
    2.82935292876456e-17, 7.36368024018167e-19, 0, 0, 0, 0, 0, 
    5.63068426483033e-10, 4.11272234950428e-15, 0, 0, 0, 0, 0, 0, 
    8.45985634348976e-19, 0, 1.57432586567363e-18, 0, 0, 0, 0, 0, 
    4.3582941061943e-12, 1.89613668819647e-11, 0, 3.12920534192198e-12, 
    4.46058664581686e-12, 1.02679297358737e-07, 3.13878657446927e-09, 
    1.7459968115544e-10, 4.48018046256736e-08, 4.23970065449604e-07, 
    5.58077297979569e-09, 7.24277177605634e-12, 1.1011221097995e-20, 
    0.000450310475634586, 0.000600424077845748, 5.93622411325357e-06, 
    2.35649358351957e-11, 3.18906939027623e-09, 2.432085359337e-09, 
    1.64512716440366e-07, 2.7728039878033e-08, 1.20467683901546e-06, 
    4.78552443686829e-07, 3.41919224440452e-09, 1.04792756630653e-11, 
    8.71633772505299e-06, 1.11814487462435e-05, 1.85838256344394e-05, 
    2.51538324958565e-07, 1.12124027676496e-06, 7.24193732555567e-08, 
    4.83030056444068e-06, 8.01070241238645e-06, 3.8343853016033e-06, 
    2.75233770125933e-06, 5.9861208059317e-06, 6.64529552529086e-07, 
    1.59893885483033e-06, 2.1695348221179e-06, 0, 3.95334462765719e-06, 
    5.10141694914848e-06, 9.61744355147693e-09, 4.04525516673941e-06, 
    4.23121783205248e-06, 2.66506070645046e-06, 3.05370052239471e-07, 
    2.61411017120009e-06, 9.40915718992265e-10, 3.95529805724937e-06, 
    2.80427496000321e-06, 1.06007912752816e-08, 6.69484934761099e-05, 
    2.93257201895194e-05, 2.90019952755501e-06, 8.65998762214043e-06, 
    2.51666577161153e-06, 2.32527536504382e-06, 2.09912202631016e-06, 
    5.89086454359539e-09, 1.37223786050495e-06, 1.32497145450287e-06, 
    1.52842335901117e-06, 2.26590125844243e-07, 2.58856353627199e-07, 
    4.58816902569605e-08, 0, 0, 0, 0, 0, 0, 1.07502594145789e-09, 
    5.5634357830948e-08, 6.17392025734205e-06, 2.24268356201642e-05, 
    1.44442932890541e-05, 6.74620305192817e-05, 0.000161877190815225, 
    0.000102402628243079, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.50303097346877e-07, 
    1.86935941845912e-05, 5.77110268005499e-05, 4.27028821850334e-05, 
    1.2772623901374e-05, 5.1882985313793e-07, 1.94170042962439e-06, 
    1.28811217134378e-06, 4.42797347456324e-06, 4.70296494709755e-17, 
    5.79801210626823e-21, 3.78164053232414e-07, 8.58069647379929e-05, 
    7.96551914497666e-06, 3.12497426641525e-06, 2.31874603980403e-06, 
    3.56829740345444e-06, 2.28799132919581e-06, 1.89541644156336e-06, 
    8.46261276434173e-07, 2.90462037293854e-09, 0, 1.34500191385235e-13, 0, 
    0, 3.22896679896157e-12,
  2.79048721303451e-06, 4.08187446638325e-06, 7.91270394971859e-06, 
    1.13223544135134e-20, 1.18327560588112e-06, 0, 0, 0, 0, 
    3.12220268242076e-05, 1.99893004678899e-05, 0, 0, 3.68293930538866e-24, 
    6.7241821254936e-11, 0, 4.43561001458312e-11, 5.44189037165997e-08, 
    3.1149630428147e-20, 3.31554114903932e-17, 0, 9.08044890671011e-18, 
    6.22640124274061e-20, 0, 0, 0, 7.62253797521325e-28, 0, 0, 0, 
    3.43804530609344e-18, 3.0338262964316e-17, 1.09529720137045e-09, 
    8.91161462557488e-09, 8.41118687782269e-10, 2.41424521497789e-07, 
    7.23170338821699e-08, 1.6620309448218e-10, 9.93972369305624e-12, 
    3.49694372396112e-08, 2.72610747530142e-21, 2.90926131623476e-09, 
    0.000113754815024615, 0.00063218435978405, 9.16381912017495e-05, 
    4.18920636217971e-08, 3.36900431002564e-07, 6.72273707545158e-06, 
    2.45510677864215e-09, 4.23462291741453e-07, 2.37278304900595e-06, 
    2.1870432327732e-05, 3.0817149803669e-06, 9.45096876932643e-10, 
    1.96570361307742e-07, 4.30133931966294e-07, 1.67787638714242e-05, 
    8.96563808977249e-07, 2.73820925946429e-07, 2.66900877039372e-08, 
    7.46790137995905e-08, 6.39232043160835e-08, 1.27221162232138e-07, 
    5.52228369771394e-07, 2.51744388334758e-07, 2.41611305588745e-07, 
    1.74557380029971e-06, 5.53379095156069e-06, 6.06648300253112e-06, 
    5.67252348025766e-06, 2.91971684603021e-06, 4.29661198284043e-06, 
    4.62644087321963e-06, 4.02450280484989e-06, 4.09811552555509e-06, 
    1.79750790051129e-06, 1.76019810657368e-06, 1.72460618734681e-06, 
    1.6900855798496e-07, 3.90306486498862e-07, 3.00233344169065e-07, 
    0.000127276606687475, 0.000307992248067349, 5.21371918466403e-05, 
    7.27597086153941e-06, 2.36104820925537e-06, 2.40829463919372e-06, 
    1.99919442981553e-06, 1.10619622316032e-06, 6.84434154046346e-06, 
    1.42850263221374e-06, 1.59201275281431e-06, 1.79848520792246e-06, 
    1.07159529543485e-09, 0, 0, 8.74323160986438e-10, 3.70934656919685e-06, 
    3.20029195051026e-06, 2.29630964077736e-06, 1.60801454406485e-07, 
    3.06431519699515e-07, 4.22814914149711e-11, 1.10274418281047e-05, 
    8.24882618750598e-05, 0.000102687647096721, 0.000127355424139061, 
    0.000201005947463613, 7.92705480962984e-06, 2.45585979933172e-20, 
    2.18066499568138e-21, 4.73912943706601e-18, 0, 0, 0, 
    2.62694993862999e-17, 0, 0, 0, 6.02512970137197e-06, 
    2.50386944787054e-05, 8.02994920254572e-05, 5.20538631556688e-05, 
    4.93681934855305e-08, 1.80443070675365e-09, 4.29703054405329e-06, 
    1.10218025034157e-06, 5.51254802681186e-07, 1.89850921062179e-11, 
    5.28733670193798e-20, 7.23259463256793e-05, 5.84990130343708e-05, 
    2.96747148714943e-08, 5.05436917201378e-06, 2.21071191041538e-06, 
    3.30957789948342e-06, 1.08990763609649e-06, 4.7198887982307e-09, 
    1.73420780564057e-07, 2.39421912714175e-10, 0, 2.03797094670554e-09, 
    6.70847530394216e-09, 1.00261004587696e-10,
  1.8283877139303e-07, 1.38433077738542e-07, 5.36651515813813e-05, 
    2.75363822859269e-05, 7.50620197439642e-06, 2.32592917507756e-07, 
    5.45421002946961e-21, 0, 7.05249965971803e-05, 6.74645636849178e-05, 
    1.86889843287522e-18, 1.10136710137773e-22, 4.05994407056072e-18, 
    5.87406139951782e-19, 1.89175295652792e-23, 2.98445919293708e-10, 
    2.84340724764039e-06, 1.35854737642474e-21, 3.70651560065712e-11, 
    2.95931356768844e-19, 7.23796066740436e-18, 0, 5.69638303720058e-19, 
    1.3322026495108e-19, 0, 4.41767860318745e-08, 3.53090303034687e-21, 
    1.40412719848481e-19, 1.35833375570229e-19, 2.35648758164999e-10, 
    1.59759528641517e-16, 7.61700573383564e-18, 8.29622244598558e-08, 
    5.93727359383603e-17, 1.83435950927211e-07, 2.17869098233048e-08, 
    5.05764239929256e-07, 5.59261205406886e-12, 3.54544948942745e-07, 
    2.16279304561977e-08, 9.89902831916182e-09, 1.9809093147617e-05, 
    1.33387259645904e-07, 0.00016154975217575, 0.000141091389225561, 
    1.52772003004488e-05, 1.14630029378175e-05, 1.4519142123805e-05, 
    4.16105870577826e-09, 7.74907221507387e-08, 7.74948905621364e-06, 
    2.67476526802396e-05, 1.40030669181481e-05, 2.84309432547269e-06, 
    3.56665659812137e-07, 3.98315634480902e-07, 2.36155215082296e-07, 
    7.8732945473248e-07, 1.3507520797752e-06, 1.29038695495965e-06, 
    1.18177433174533e-06, 1.27068282063498e-06, 4.58319425913699e-07, 
    5.14820706127812e-07, 8.45245352629184e-07, 7.03799613662908e-07, 
    9.092910055675e-07, 1.64339393157014e-06, 3.74692123114916e-06, 
    1.50234374400615e-06, 1.49898758133898e-06, 7.79309888605873e-07, 
    1.22126869973204e-06, 1.07890412305426e-06, 7.28346947238738e-10, 
    1.10562129402558e-05, 9.44571480841646e-09, 1.22666580017347e-07, 
    1.66584129121764e-06, 2.27611131161001e-07, 1.13541976809276e-05, 
    0.000233889208722765, 0.000342514578122403, 0.000183568548261825, 
    0.000142832747249806, 3.03845075584047e-05, 3.88324454706052e-06, 
    3.23684429476982e-11, 2.38880264878977e-06, 1.67544185866814e-06, 
    1.46855508992249e-06, 1.72260709707241e-06, 1.09217953643468e-06, 
    7.74514523843855e-09, 1.69428855246472e-09, 3.76644708081385e-11, 
    1.32410973863684e-06, 4.4722315972383e-06, 1.12682915851261e-06, 
    1.20743494806932e-05, 2.80181502914617e-07, 1.49762086483606e-07, 
    3.83308029853074e-13, 0, 4.04214098513645e-05, 0.000105213418977064, 
    0.000147352047495301, 3.38311822423716e-05, 3.37849658251594e-08, 
    2.78495417553198e-17, 6.56199412298615e-18, 1.08776491097208e-23, 0, 
    8.73998872615515e-12, 2.09443240131356e-10, 6.4482746704338e-09, 
    4.89211336714339e-12, 6.0759958244887e-10, 1.49715262002346e-09, 
    4.60546575369474e-11, 1.15803594794442e-06, 6.85393812140515e-06, 
    2.97340485618134e-05, 1.03833542306373e-05, 2.49616116197091e-09, 
    9.45160095433981e-07, 8.30681424098461e-07, 1.25755907566641e-09, 
    4.07646960853975e-10, 5.26363725060372e-12, 3.22544792140145e-05, 
    9.46628366697651e-05, 9.08741661972007e-05, 1.21308768333038e-07, 
    4.957129071111e-06, 2.56755451700277e-07, 4.04331666504486e-09, 
    1.44688610556778e-06, 3.50625527524027e-06, 1.01324038956291e-08, 
    2.37940472373342e-07, 4.10699504428741e-08, 1.37090886075136e-05, 
    1.48025557914482e-05,
  6.50204499776534e-11, 6.13527476204779e-09, 7.11372221800362e-05, 
    6.10642572125098e-05, 7.80073024272439e-05, 3.31334146151155e-05, 
    1.15495424760356e-19, 6.59669897976239e-24, 2.84542414435888e-24, 
    4.40775255009658e-22, 2.38357466766323e-20, 9.17462222258862e-20, 
    4.564498895843e-17, 0, 0, 5.58915899675733e-23, 9.54729005948076e-06, 
    1.77049498579348e-07, 2.32385831620081e-10, 2.0626743109577e-26, 0, 
    9.43960672287628e-23, 4.25286194016543e-24, 5.24109349170361e-19, 
    1.87711447692498e-20, 6.69737068700222e-17, 2.08310690379504e-19, 
    5.04870979341447e-29, 4.4374377291015e-16, 1.07904738375363e-05, 
    8.4220545439588e-06, 2.30992556621005e-18, 8.71021407051183e-16, 
    2.77682763792558e-09, 6.44711766735201e-23, 4.98824384897577e-11, 
    3.96386802627744e-20, 7.31893513898797e-10, 2.14354360851442e-12, 
    3.7488298301083e-07, 2.83794266094595e-07, 9.48095936217522e-06, 
    1.35200871089273e-06, 6.51698935398971e-05, 0.000215488208256343, 
    8.62523858444876e-05, 3.64956662929721e-05, 3.23629021191796e-06, 
    2.55412162808696e-10, 4.42752775100864e-09, 1.83544370183539e-08, 
    1.40644381425798e-05, 9.19802926859811e-06, 1.56640876196013e-06, 
    2.3963880517679e-06, 3.98385717129097e-06, 5.02669171617889e-07, 
    7.16726118618548e-07, 2.37747878744227e-06, 8.84949190118096e-07, 
    4.59319852069082e-07, 4.11196375286188e-07, 5.36772335543265e-07, 
    5.37408512605712e-07, 1.55137433646588e-07, 1.27143359732163e-07, 
    6.00895491777692e-12, 5.16431712680987e-07, 6.3228215319751e-07, 
    4.65267583611069e-07, 1.48500429240728e-06, 1.02957234388746e-06, 
    1.27389031560563e-06, 1.13317951191781e-06, 1.65414925684047e-06, 
    2.86312300522922e-05, 4.66900833449119e-05, 6.04591071681495e-07, 
    2.15389994518784e-07, 9.55671356513325e-08, 7.15481329986545e-08, 
    6.15602152381135e-05, 7.47051507044139e-05, 0.0001352295876083, 
    0.00014565979369297, 1.65495558942236e-06, 3.57474904690889e-09, 
    2.08027009529737e-06, 5.47454153307968e-07, 1.11557500617463e-06, 
    1.83412738837323e-06, 1.66040980545174e-06, 1.49147822462467e-06, 
    7.37538629229135e-07, 7.17323374911848e-07, 2.82573764582952e-08, 
    4.39325851345988e-06, 9.11911645945188e-06, 2.38776330496446e-05, 
    5.28802604328172e-05, 4.64104919753443e-05, 5.84648080709306e-05, 
    6.51192826655336e-08, 5.09463565351854e-20, 3.75452944566068e-05, 
    7.1764179566627e-05, 1.06676485994456e-05, 1.10391335065113e-06, 
    2.26484028630395e-20, 4.8584514422151e-18, 2.67343306207962e-20, 
    3.65018510765836e-21, 1.19951839514452e-11, 1.24445488570001e-08, 
    1.91866847933857e-07, 5.03870149979217e-09, 8.29525445851281e-09, 
    1.79369297017551e-07, 5.26524926719568e-08, 5.30139660886767e-09, 
    2.91409454509302e-08, 4.2606864048675e-06, 7.65414319927035e-05, 
    0.000176245676851285, 8.35625257952895e-05, 1.08288675216065e-06, 
    1.57664612635516e-06, 2.6868515030434e-06, 3.01314344490923e-07, 
    1.34682134447943e-07, 6.90720000090813e-08, 8.36549936185513e-05, 
    0.000206372689237282, 6.05446753559413e-06, 2.17262845041327e-07, 
    1.58374103998207e-09, 1.70395234822847e-10, 3.84703243665766e-06, 
    1.6169001691567e-05, 5.05543436556533e-06, 5.71608415012517e-07, 
    1.1825355340185e-06, 6.96083693890651e-07, 2.09698354276068e-06,
  7.03385837612126e-10, 1.07099003432548e-05, 7.15863873187884e-06, 
    0.000221325195037774, 0.00018252012471391, 3.3777177303541e-06, 
    3.45501822555841e-11, 1.5768879276623e-18, 1.23206101324462e-23, 0, 0, 
    6.04163871020913e-17, 3.29560908685171e-12, 1.30606532470618e-11, 
    6.72945771011075e-19, 2.22533271007699e-17, 5.04581509878332e-17, 
    1.90982739109902e-17, 2.99014406627375e-10, 8.43938749103269e-21, 
    6.64546467640231e-24, 0, 7.37252019646649e-13, 2.18532459440608e-17, 
    3.98446119193225e-17, 1.49928498688135e-18, 1.00909435116759e-20, 
    1.8200541954916e-17, 1.07403078633396e-05, 1.87630829688726e-05, 
    5.9993363011644e-06, 2.14558332378315e-17, 9.55971110064531e-12, 
    3.89804936001635e-09, 4.0997977681354e-06, 1.38914328696262e-17, 
    3.02601631451141e-09, 0, 0, 1.88639823246563e-18, 4.56917886943483e-09, 
    6.79022465695744e-09, 2.53299940375603e-05, 7.33410862708191e-05, 
    0.000411789482955805, 0.000432898895519654, 0.00023030834429321, 
    6.7386277381132e-05, 5.81818860087688e-06, 4.00694693422255e-05, 
    6.77788860483995e-10, 1.30729314317067e-05, 1.73689520669772e-05, 
    1.81194703643158e-05, 1.58254732961314e-05, 1.80397310944508e-06, 
    9.66622318320954e-06, 1.53166204646705e-06, 2.6526619239663e-06, 
    1.84199923754954e-06, 1.49502001923098e-06, 1.49644495963346e-06, 
    1.46763502894062e-06, 1.66318684771482e-06, 5.83105606922747e-06, 
    5.01472071409053e-06, 7.04184563973144e-06, 7.10080156004267e-06, 
    2.71290864997787e-06, 3.1568066268152e-07, 9.26922692358123e-07, 
    9.03054830401602e-07, 7.55456137856532e-07, 8.65290338978933e-07, 
    3.24424795384936e-07, 1.26835736173455e-06, 4.00285546248785e-05, 
    4.96887770325399e-05, 3.92374151416628e-07, 1.68420775411739e-06, 
    2.36147245179285e-07, 5.44459760339134e-08, 1.37965087089864e-07, 
    1.02347409470572e-07, 1.80459685389465e-07, 1.06832446014613e-08, 
    1.2378024963014e-07, 2.12422216960156e-08, 7.08298381052632e-07, 
    5.87538783434176e-07, 3.21547784441719e-06, 1.86635866052562e-06, 
    2.58306993045326e-06, 3.63522513943815e-06, 2.87828257765063e-06, 
    4.86384783420059e-05, 5.28183086178075e-05, 3.24322981102527e-05, 
    2.86763695981569e-05, 5.21301370253325e-05, 7.70279958607016e-05, 
    0.000263814057702826, 0.000169569831394646, 0.000108247935328878, 
    7.99452194700016e-05, 1.44357661101942e-05, 7.49751246079992e-05, 
    0.000224803236071685, 5.9795197832362e-05, 8.9321204936238e-11, 
    2.34643685348034e-24, 2.11341507196747e-12, 4.4083759616883e-09, 
    9.66407770435546e-09, 1.16257561595106e-05, 2.7617187275346e-05, 
    1.29677062781795e-05, 1.2178191744581e-05, 4.18095683068177e-06, 
    1.5400219335803e-06, 1.64528766377896e-07, 3.30426047719313e-05, 
    0.000217901623896204, 0.000329133186647288, 9.79724667818929e-05, 
    6.37884074160833e-09, 1.70742725263507e-06, 1.70285344773782e-06, 
    9.88457016344252e-06, 1.16278004743091e-05, 8.1813541456863e-07, 
    3.14419484879375e-06, 0.000201771422396146, 9.22576942666835e-05, 
    1.23749104579969e-09, 6.75473132584462e-08, 9.39940796200047e-10, 
    1.32903208460998e-06, 5.82956988753919e-06, 9.05502483024873e-06, 
    6.8358139307853e-07, 6.55114693647462e-06, 2.06756436941615e-06, 
    2.66554082599967e-06,
  6.98173029975317e-08, 4.76477920586762e-06, 4.2216126421807e-09, 
    4.70933945232379e-05, 6.69553009376244e-05, 6.37780921668357e-06, 
    5.48612955121496e-05, 7.33729313332058e-05, 4.01213915179167e-05, 
    1.61744535066717e-06, 1.45667225126969e-07, 3.11643918444467e-19, 
    6.96131249298252e-13, 1.74309498172376e-09, 5.34948624723601e-11, 
    3.31472179571699e-17, 5.16777839189056e-16, 9.69354572974829e-16, 
    4.89267312399467e-16, 4.2254096204521e-18, 4.56951283908031e-25, 
    1.00911589898813e-18, 6.82862884920548e-17, 2.07056460645264e-16, 
    5.60924415925376e-17, 4.51661669823117e-25, 2.66369435427576e-18, 0, 
    4.00016957815967e-07, 1.47829768500404e-05, 2.01901773935226e-05, 
    2.21719681965905e-08, 4.95835001732372e-07, 7.71512111355768e-05, 
    7.36772857926196e-05, 7.62520260453595e-08, 2.98254679072145e-17, 
    2.89465196158273e-11, 6.13068361668051e-07, 2.27536217255129e-12, 
    2.16162509534333e-07, 6.22625415995752e-09, 1.51480561775136e-06, 
    1.76575215938747e-08, 2.1437723117655e-05, 0.000228941687746164, 
    0.000420586441195556, 0.000280878566904153, 0.000120051404661341, 
    1.25278659035175e-05, 3.43121645643859e-06, 2.04838203190791e-05, 
    1.12194433228619e-05, 2.07871246769799e-05, 1.85793437040597e-05, 
    8.33562017363235e-06, 1.05394800213844e-06, 5.34779983714363e-07, 
    2.94396690963731e-06, 2.4684659041625e-06, 2.68711281406321e-06, 
    6.68295301655057e-06, 1.20349002605204e-05, 5.13628904670473e-06, 
    7.81532347547033e-06, 6.52265474511031e-06, 8.78970321911686e-06, 
    1.70231270189742e-05, 3.11453832912481e-05, 1.11596903103088e-05, 
    1.3222384691672e-06, 1.71477384064227e-06, 1.8749780702553e-06, 
    4.93983140365381e-07, 1.22040979796996e-06, 6.98639716105841e-07, 
    7.13746198314814e-07, 2.39572500286149e-05, 3.85405038582948e-05, 
    3.65626102643311e-06, 3.34780285792204e-06, 2.12120219632966e-08, 
    2.56767242014978e-14, 5.70871242117568e-08, 3.89909965215288e-08, 
    3.88991290994993e-09, 5.02985656689412e-08, 4.6836978964539e-07, 
    6.84047930940088e-07, 7.65214179188996e-07, 1.90765109833953e-06, 
    1.76895350811166e-06, 1.20745625346494e-06, 2.42958606753005e-06, 
    1.51865053565901e-06, 0.000285907005229586, 0.000132405473839768, 
    8.81818871124832e-05, 5.32446452363668e-05, 8.61302835141659e-05, 
    0.000286502259070523, 5.38463995656778e-05, 3.42109926686242e-05, 
    2.78942740612299e-05, 5.7096506603346e-05, 0.000147609732812483, 
    0.000327406172359957, 0.000164104171687065, 9.35838078922088e-06, 
    2.08722822529561e-11, 4.35684703275086e-07, 5.28490702975118e-07, 
    3.34193929041571e-08, 3.19670198297459e-06, 1.9133827541973e-05, 
    4.49737836365515e-05, 0.00014457046687456, 0.000315239801186612, 
    0.000188072172284885, 6.52893421603009e-05, 5.33508565060881e-05, 
    0.000178770326265354, 0.000259512026140362, 0.000184194424931131, 
    4.70008090780257e-12, 6.09642802682283e-06, 4.94153886696585e-06, 
    1.17739329196437e-06, 9.7146181852676e-06, 1.09513846915696e-05, 
    3.03588644496718e-06, 0.000113289429336367, 0.000115271284380734, 
    0.00012441335264614, 1.39856929255818e-05, 1.07077267891557e-06, 
    8.38797185563769e-06, 1.10467402334062e-05, 2.78469356017841e-06, 
    1.83535121045113e-05, 1.75549924183213e-05, 2.8349064636457e-06, 
    9.8459334202794e-07, 1.59238254236077e-06,
  2.27391514989051e-08, 5.29008025658997e-10, 8.73548063785178e-12, 
    3.79032810819692e-05, 3.63801397857858e-05, 4.5877324983617e-06, 
    4.86025971045486e-05, 7.35756441378824e-05, 7.52907929151668e-05, 
    2.13555267556028e-06, 1.75870873786485e-06, 7.42203617312533e-06, 
    3.57968149439041e-05, 0, 2.46827263149572e-11, 1.67131813867806e-21, 
    1.03961062547845e-22, 0, 0, 1.37025488405069e-10, 6.23734445439971e-11, 
    7.72408056509267e-10, 2.67002037069306e-08, 1.90416696022996e-08, 
    4.5011068649297e-12, 7.18685796524477e-17, 8.71609496536307e-10, 
    6.74067956795634e-09, 1.48675260364727e-09, 6.76201983964147e-09, 
    6.58817724289129e-16, 3.50047889976321e-08, 4.42504588286996e-06, 
    0.000108823121640689, 0.000150987486937158, 0, 4.28811917478234e-18, 
    4.21225395374395e-17, 2.162843327373e-12, 0, 2.54822264264445e-11, 
    2.81917499453116e-10, 7.20058889885628e-09, 2.86657901250055e-10, 
    2.32631866264225e-09, 2.50125229565693e-05, 4.08892216384282e-06, 
    0.000235762959626749, 0.000294405013262133, 0.00015485488523801, 
    1.08425151641361e-05, 1.95593911296305e-05, 3.66256635365209e-06, 
    7.46361279882358e-06, 8.54977776170618e-06, 2.45218630459787e-06, 
    1.16449446220604e-08, 3.52022155371227e-08, 2.59669697527919e-06, 
    3.77122992342082e-06, 3.78367207171343e-06, 3.4818793695061e-06, 
    2.83770288355801e-06, 2.26872527421835e-06, 3.43883572412808e-06, 
    3.03857802164167e-06, 2.21331733519604e-06, 3.70908678769239e-06, 
    9.23255575285648e-06, 2.54583544352167e-05, 4.30654864053852e-06, 
    5.95900360408536e-08, 8.25337243860426e-09, 1.8699662122035e-21, 
    1.59970207535514e-07, 5.39824701231165e-07, 8.91768128188823e-08, 
    2.95212565453963e-07, 3.09775988501424e-05, 3.60390301288512e-05, 
    3.29976397753479e-06, 2.85940585340841e-06, 1.31558351772093e-06, 
    4.64240850677241e-08, 2.18905581013725e-07, 1.11747026903721e-07, 
    3.83743036743668e-07, 9.16926741096015e-08, 0, 7.16638406717055e-07, 
    1.17834200763331e-06, 1.59463111998288e-06, 1.61490131951134e-07, 
    2.71246995764222e-08, 0.000102830084531713, 0.000214856008676211, 
    0.000324532466226425, 0.000177891806236482, 0.000267405233090809, 
    0.00044458809701085, 0.000288181563850501, 9.99369098473916e-05, 
    1.99746131183312e-05, 1.96493849354061e-05, 7.15941067798763e-05, 
    0.000134253642126164, 9.62432769778954e-05, 3.38551415072969e-06, 
    6.49631199650414e-06, 2.23960246351999e-05, 4.56755501482918e-05, 
    3.10560825949967e-05, 1.11308632658314e-06, 7.54828861594033e-06, 
    8.84010289982664e-06, 7.05955646626722e-05, 0.000232351800846181, 
    0.000476983868073862, 0.000564595203585006, 0.000353100116767797, 
    0.000225603113028521, 0.000258054375763673, 1.64647222333344e-05, 
    2.87370065886351e-12, 3.39664060237155e-07, 4.04109930137536e-06, 
    1.50491326185382e-06, 2.61563916452595e-06, 1.25032094158164e-05, 
    4.42153703391818e-06, 6.39244650366697e-07, 4.78993645926756e-05, 
    0.000191996784747236, 0.000187315004206971, 0.000100872994684223, 
    1.01772492470194e-05, 1.16915623472584e-05, 1.0985892745659e-05, 
    1.55437869632062e-06, 9.99682312660552e-06, 1.88980698622448e-06, 
    8.3558722946274e-07, 2.39074294906361e-07, 2.02659020167325e-06,
  1.23560929510314e-08, 1.80594701579717e-06, 9.51771123039167e-06, 
    0.000124815644609357, 4.58502773185849e-12, 3.758776810562e-10, 
    1.50026860249691e-19, 1.226744363505e-05, 1.88965554086573e-05, 0, 
    2.80189703573111e-05, 0, 0, 0, 0, 0, 0, 2.94454460820827e-12, 
    7.28103273543218e-11, 1.08691180028172e-09, 3.46353691081073e-08, 
    2.00662255801308e-07, 4.89457800204947e-06, 4.76948320547484e-06, 
    9.87117135774006e-06, 5.64812811250699e-06, 1.30854673492049e-08, 
    3.74018664023126e-09, 9.95467987791859e-16, 5.00949373068732e-11, 
    8.6697428729822e-06, 1.52459837442173e-07, 4.3542882882683e-08, 
    0.000172729899085066, 4.69416336007896e-05, 2.15879591018703e-05, 
    1.78036248614561e-05, 1.53112251935648e-05, 7.36201358776221e-05, 
    1.44622419523854e-05, 1.34555780808736e-12, 8.71111448979849e-23, 
    1.76936292209132e-11, 0, 4.23742508638205e-12, 3.81531103641655e-10, 
    3.39419957107843e-08, 2.40674611773699e-08, 6.48329998246331e-05, 
    0.000186523243636584, 0.000107538153143374, 8.88781007958852e-05, 
    1.12447682710284e-05, 2.97903429271357e-06, 5.50957956983242e-07, 
    4.63794312088356e-08, 2.74318054315625e-23, 7.34531287895991e-21, 
    3.84475691889789e-06, 5.96575133465417e-06, 4.93833911827951e-06, 
    6.74737526339223e-06, 5.20695268475896e-06, 5.31721886834791e-06, 
    1.91408518177241e-06, 3.01091440600559e-06, 4.60704426302596e-06, 
    8.90664130255969e-06, 3.36693421602189e-05, 0.000156687887780193, 
    6.62471476913805e-05, 1.21953441878415e-07, 8.33291759771573e-10, 
    1.68639430725748e-11, 0, 1.90154675933959e-06, 6.68701491949019e-07, 
    1.58697271477537e-06, 1.03500716766695e-09, 2.33608262167065e-05, 
    3.1553576899453e-05, 3.8130637680883e-06, 1.37716110268482e-06, 
    1.02680705206193e-06, 6.50680459710941e-07, 1.3548018334637e-06, 
    1.46672303767152e-06, 3.80330602881545e-09, 6.42653665978462e-08, 
    2.89852076368812e-07, 7.45070688977499e-07, 1.25912570312508e-06, 
    4.31853566991075e-09, 3.4907705166954e-06, 0.000118811343931281, 
    0.00015739367389334, 0.00023715937458167, 0.000173632059746061, 
    0.000268868356353856, 0.000213636561682454, 0.000296734714642879, 
    0.000288858591274175, 0.0003093481489073, 0.000137257024985159, 
    0.00015807302585481, 0.000188954011127991, 9.42026841212422e-05, 
    0.000119955726415422, 3.44497247440476e-05, 3.67452943414541e-05, 
    1.40248493819086e-05, 2.90833704516921e-05, 2.90660227455158e-25, 
    1.19515352897271e-05, 3.4522973632958e-05, 3.81434937500979e-05, 
    0.000103045026461047, 0.000251350837319811, 0.000375301995652356, 
    0.000200796396658531, 1.42497047054204e-05, 3.74042267086208e-08, 
    1.28361332882633e-06, 4.87329821246144e-07, 3.12128077065699e-07, 
    1.1773802475215e-06, 8.68502375648393e-07, 1.95709655255339e-06, 
    3.42707682654705e-07, 7.28164369291273e-06, 8.32851319943122e-05, 
    0.000285275811358447, 0.000323105513958434, 0.000243108855514073, 
    7.51853757403298e-05, 1.47562614843054e-05, 1.56066738236008e-06, 
    6.43622227381428e-06, 2.91418710674867e-06, 1.02589312619972e-05, 
    1.32635597033502e-05, 1.06325676029719e-08, 6.67258896732791e-08, 
    2.46422793246743e-15,
  1.57678260969578e-06, 2.11867663725741e-11, 1.72853517890566e-05, 
    2.1488812278175e-05, 1.00113016107938e-18, 4.1907710944385e-29, 
    1.81432203879529e-05, 4.61861789497242e-05, 4.43992721899252e-05, 
    2.99881138605622e-05, 0, 0, 1.67351227187505e-11, 0, 0, 0, 0, 
    3.42113626054192e-11, 4.72766826881508e-10, 1.25107050860163e-08, 
    4.19987500932856e-06, 1.53329752151584e-07, 6.64164824394916e-06, 
    7.95894573907916e-06, 2.99233909212138e-05, 6.44182741072355e-07, 
    4.63981823276534e-10, 3.14431037178164e-06, 1.09212951507339e-07, 
    4.07331598346547e-06, 1.37902157414365e-05, 1.86359873370753e-09, 
    5.54936653051117e-05, 0.000191339866921115, 0.000128728814525662, 
    7.30818344161732e-05, 3.64367573095798e-05, 4.06140150377649e-05, 
    4.1834958586311e-19, 3.54223982103026e-06, 3.57356162592624e-13, 
    1.39218861186479e-10, 1.02496211576073e-19, 3.33148029651375e-11, 
    7.22309092278097e-09, 3.82320557736137e-09, 3.48236700658787e-10, 
    1.7598577675921e-11, 2.51414053947244e-11, 1.36954338748852e-17, 
    0.000254216250882968, 0.000116291603861428, 0.000112817291765875, 
    1.37337657643606e-05, 5.9704836628326e-08, 6.77534316943727e-09, 
    1.31078923532243e-09, 1.70597403147649e-07, 2.76189077346152e-06, 
    6.10555392879673e-06, 8.49918272292987e-06, 1.42933907367735e-05, 
    1.7679878026072e-06, 9.85717553677217e-07, 1.4284967337075e-06, 
    9.81537980115193e-07, 2.97655232260177e-06, 9.66950932807678e-06, 
    7.38676790686658e-05, 0.00038386429072483, 0.000453146959065327, 
    7.98226300645879e-05, 4.85796154221824e-09, 2.07810959464116e-10, 0, 
    1.23814146767286e-06, 1.78829714513238e-07, 5.79875700346835e-07, 
    1.16946567032625e-06, 1.18726520705301e-11, 8.04089301567072e-06, 
    1.85577188478287e-05, 4.97201203921546e-06, 3.47074549395466e-07, 
    5.32770698288183e-07, 2.70644981350706e-07, 2.01549122514505e-06, 
    1.17882896078555e-08, 2.62778417281562e-07, 1.08638320326137e-06, 
    4.78583124199609e-07, 2.03247102644063e-07, 5.10729307092068e-09, 
    1.09751210026698e-05, 3.6179748394874e-05, 8.43813602309161e-05, 
    8.35854361713369e-05, 0.000176937158784398, 0.000177654591214252, 
    0.000112022411885257, 6.88221756068628e-05, 1.81202016965531e-05, 
    2.4995191214381e-06, 2.68117410730287e-05, 5.23113223979105e-05, 
    8.83393898851941e-05, 0.000120719440993832, 3.13943153241342e-05, 
    0.000124630816623263, 0.000160581732909774, 7.62825637388167e-05, 
    4.93702455449096e-11, 1.42495760154685e-21, 1.79924338059773e-05, 
    3.87023861328445e-05, 4.46125814887319e-06, 2.66529229199425e-06, 
    1.09645199197003e-06, 8.13985668526082e-06, 8.07863144749756e-06, 
    1.22552436148677e-06, 6.54197190200567e-06, 6.43820079856291e-06, 
    2.26151894692873e-06, 1.34699208048643e-06, 6.51553466978441e-08, 
    2.0308262239324e-06, 6.64260770997276e-06, 2.37374182107678e-05, 
    0.000123343195806541, 0.000269570251405238, 0.000314040857806301, 
    0.00021668395713842, 2.99658026091753e-05, 4.57650295452692e-06, 
    5.81245734776977e-06, 2.41118735406501e-06, 3.22367476319498e-06, 
    1.3495759655721e-06, 5.13290432075608e-06, 1.69501045090456e-05, 
    3.0938775884796e-07, 2.42742684995345e-06, 3.61454261410694e-10,
  1.29982047835401e-09, 1.25255436570559e-05, 4.29408898931924e-05, 
    3.61078845771405e-05, 5.04440446513189e-06, 7.92421803100939e-19, 
    3.83146070781841e-05, 6.23481509860332e-05, 6.13406868421099e-06, 0, 0, 
    5.02538284155546e-12, 3.30294262611836e-10, 0, 0, 0, 0, 0, 0, 
    4.2602914795717e-11, 2.57304266497226e-09, 3.41191050679573e-21, 
    2.16036377237237e-17, 5.80109650707898e-16, 1.02245518961604e-17, 
    3.69603444004058e-07, 3.56467683174136e-20, 2.47940202397406e-11, 
    5.79827828853664e-10, 6.53848757252359e-10, 2.52098343502156e-13, 
    2.98610227221562e-06, 2.89356724127521e-05, 2.14771743652399e-06, 
    5.04830729404295e-05, 2.64014568519168e-05, 2.14627755785901e-06, 
    9.03294933620206e-20, 4.81593185461706e-19, 4.94969138656428e-19, 
    6.15530541393134e-06, 9.4744561374836e-06, 4.00270579572762e-05, 
    5.30101678198034e-05, 6.89072341832274e-05, 1.44535017309706e-05, 
    1.78463860299124e-05, 1.67962061783205e-09, 4.14832925414253e-11, 
    1.94367408835994e-12, 6.36504566405462e-05, 0.000249066968191575, 
    9.64862583985003e-05, 7.24102000013715e-05, 2.53229625039562e-07, 
    5.72416033362917e-08, 6.07646903140051e-09, 5.45550333051786e-07, 
    6.7017152463161e-06, 1.00990746059256e-05, 1.67419462246343e-05, 
    2.27089376723258e-05, 2.24248210623249e-06, 4.57810902404923e-07, 
    3.59275176249551e-06, 3.47843232916021e-06, 1.57397432247712e-06, 
    3.91373877391781e-06, 1.10943610131329e-05, 0.000115723728836357, 
    0.000352720994338739, 0.000322131564689193, 8.21380611221757e-05, 
    5.63606375828167e-10, 2.25528108666059e-10, 2.14048985253192e-08, 
    1.02374737136768e-06, 8.71682148503574e-08, 3.01395250242769e-07, 
    9.82261059172038e-07, 2.46991742840105e-06, 1.94840171940705e-07, 
    1.26389919002564e-05, 9.75073732756612e-06, 2.38105662477922e-06, 
    5.74150607607797e-07, 9.83603110588108e-07, 1.37523739614067e-07, 
    1.53511709541535e-06, 1.84951627614356e-06, 1.80369063210053e-06, 
    9.24557161926453e-06, 8.45406349083106e-06, 9.93113827596285e-06, 
    5.45857067940439e-05, 2.36270350040444e-05, 2.55522884969221e-05, 
    0.000106128418301494, 5.94562098935008e-05, 9.73298976060814e-06, 0, 
    2.0964788522444e-10, 1.97010384264802e-10, 2.34473129291174e-10, 
    6.25596179067367e-06, 5.3189296491371e-05, 5.08387955106939e-05, 
    3.32571405789889e-05, 7.96108847574605e-05, 4.45489630347188e-05, 
    2.84348209119575e-09, 2.42695413984571e-12, 2.01582731067043e-20, 
    1.75073652349539e-05, 2.58193505793754e-05, 5.25811378221793e-06, 
    7.03281158313176e-07, 4.39447202411041e-07, 3.97240284969741e-06, 
    1.00862265562288e-06, 1.26126839096107e-05, 7.50314387125792e-06, 
    6.13401884152245e-06, 1.16428105432402e-05, 9.5565960441074e-06, 
    1.05240146476169e-05, 6.23993307877825e-06, 6.5240660939695e-05, 
    0.000161425423585163, 0.000266600688348522, 0.000248083343055218, 
    0.000102460494258075, 1.29667878454683e-06, 1.22771996339548e-08, 
    3.26469003150098e-06, 9.83613820298183e-12, 2.26628428078416e-06, 
    6.601888586e-06, 3.80455321524322e-06, 6.36048952091455e-07, 
    2.12522629406429e-11, 4.93674760726653e-09, 2.76769347106785e-07, 
    6.56856008923473e-06,
  4.30893009217189e-07, 5.5135630626622e-05, 0.000111617411922943, 
    0.00010568982702937, 5.11937589382883e-20, 1.08390451504685e-11, 0, 
    2.18899684539039e-13, 1.1172935235489e-05, 5.4393967589421e-06, 
    3.03370741353295e-10, 8.93617981776276e-10, 6.82747317591808e-12, 
    2.7459823909471e-19, 8.19084893199332e-20, 2.30764311329386e-20, 
    2.00561485942468e-19, 0, 0, 2.8815211132934e-11, 6.2862532396442e-09, 
    8.64746924089395e-09, 4.26960031690521e-08, 3.87753485823677e-13, 
    6.49512200793515e-10, 3.50973584105096e-25, 1.63944060505048e-20, 0, 
    3.63921547699248e-19, 3.29255746335614e-11, 4.66802946949653e-10, 
    1.34042285503142e-06, 1.01095030566434e-06, 1.53022567604147e-05, 
    2.0387681727546e-06, 2.66916273081348e-07, 1.59518075539024e-10, 
    2.9096151385209e-08, 8.43565713582235e-08, 3.07369301853625e-09, 
    4.57742241433752e-17, 1.15031806504659e-07, 4.40335169951918e-05, 
    0.000152566529646754, 0.00019511934720943, 0.000244100036668692, 
    7.71230547366347e-05, 1.99750089519153e-05, 1.02893276666327e-09, 
    2.11854755149676e-10, 2.2670528518958e-05, 0.000218439612037844, 
    0.000135758951433728, 0.000117861013759621, 2.84589057304515e-07, 
    7.31153802879361e-09, 3.47677052535374e-10, 8.47474619517233e-08, 
    1.09887846565981e-05, 1.68658451780464e-05, 2.25472750607679e-05, 
    2.74992222645265e-05, 3.5428153274234e-05, 4.90245773261616e-05, 
    3.49772729168975e-05, 1.51889272745732e-06, 3.51800349309584e-07, 
    2.64770585781392e-09, 5.71322267712824e-09, 8.21148999221756e-07, 
    3.4148197603535e-05, 0.000156893003560519, 0.000197564969522555, 
    6.30767828069325e-05, 7.21653372943729e-10, 5.68946104393128e-11, 
    1.34916818572304e-07, 6.24683057305623e-08, 1.65200750087996e-07, 
    3.194962275586e-07, 3.08978247993377e-06, 1.36931751820101e-05, 
    1.21862575132156e-05, 7.51755947781289e-06, 1.76529112752022e-07, 
    3.92652429397525e-08, 8.39309503548861e-07, 1.76455300108142e-06, 
    4.16196908226299e-06, 5.77927289510222e-06, 6.22385869488804e-06, 
    8.09692112933088e-06, 1.42246431597265e-05, 1.04887463200641e-05, 
    8.8509518810538e-06, 4.73246799880749e-06, 1.26060813046766e-11, 
    1.04509505605391e-09, 7.42691010022122e-19, 0, 0, 2.19026512395155e-18, 
    1.07886306282577e-09, 7.40265633116989e-07, 5.5330484397214e-08, 
    6.52156185218475e-05, 4.54505309883313e-05, 5.86031649231502e-06, 
    1.6823177733288e-10, 1.91597706202284e-09, 5.6699111657804e-09, 
    8.41392016263593e-09, 1.07473341415954e-12, 2.60904425362131e-05, 
    1.3837015078126e-05, 8.06934816185155e-06, 1.30471554383208e-05, 
    5.4824023024218e-06, 6.30631131939216e-07, 2.10904098519598e-06, 
    3.9034151372104e-06, 1.13135593610845e-06, 5.47848595886602e-07, 
    3.00234512394077e-07, 1.28828382342208e-06, 7.3213414307364e-06, 
    4.65734289934824e-05, 0.000124926733176808, 0.000154845305474536, 
    0.000118931266691978, 1.33208964004681e-05, 3.6109113007625e-07, 
    1.05800038741087e-07, 2.82714995291334e-07, 1.36787542844855e-20, 
    9.46408900081245e-06, 5.9186818982767e-06, 8.19870050251724e-06, 
    4.55870667824776e-06, 5.43478881242748e-11, 1.14209736684084e-08, 
    5.26856491007339e-07, 4.81214531645781e-15, 8.79755657515757e-06,
  2.65169982120063e-06, 3.51017271448204e-05, 0.000118597038972023, 
    4.85432133454742e-05, 4.06767378765654e-10, 1.54783283934763e-09, 
    5.15167597551006e-08, 7.23401629951638e-06, 3.19013811748122e-06, 
    1.50689240007227e-06, 6.09498863209792e-06, 1.88303302238731e-09, 
    5.84596349139732e-08, 6.02733340711192e-11, 5.71676858792636e-09, 
    1.22617314362165e-19, 2.62038557108276e-21, 1.06059883530139e-23, 
    8.50686314823784e-20, 1.00355949489603e-18, 2.11833122380531e-19, 
    7.15755616017593e-11, 5.86619798327881e-19, 1.88645178935822e-08, 
    1.14195811578553e-09, 8.19365990743782e-12, 7.06541598949379e-10, 
    1.41845562960227e-11, 1.03168651316845e-12, 6.13542707015942e-12, 
    1.19248958985956e-09, 7.46571211806448e-06, 2.70759322103225e-05, 
    1.8951814442061e-05, 1.20366055183403e-06, 4.79451382584181e-09, 
    2.28034460569291e-11, 2.4630354197796e-07, 2.82397745150817e-29, 
    1.07523373412821e-18, 1.23336125049916e-18, 3.36315191161282e-20, 
    1.471848762817e-05, 4.44991603486272e-05, 6.77571875932415e-05, 
    7.76765969439983e-05, 9.23638305009282e-06, 2.4882528098082e-07, 
    3.22594188499012e-10, 3.61773502715721e-18, 6.09353752446009e-09, 
    2.86096740129726e-08, 1.24744379326171e-08, 0.000127796782529013, 
    0.000111831041931907, 4.73464631200147e-05, 4.36381305661539e-05, 
    6.09386405741161e-07, 2.10285368764406e-05, 0.000157067511629997, 
    0.000342982048635407, 0.000369911403678772, 0.000335265825892252, 
    0.000183897916446605, 3.18415210955653e-05, 2.95275782754539e-09, 
    5.161164082166e-10, 0, 0, 0, 5.86969060921822e-09, 2.57169941355107e-05, 
    0.00010051755190491, 0.000186741701434365, 7.40516719221773e-05, 
    2.71405519035922e-06, 1.86482194545303e-07, 5.39713466538744e-09, 
    2.95233054129521e-08, 7.68694333879183e-07, 9.15403087757735e-06, 
    1.37947773786536e-05, 4.85202367856561e-05, 1.49206708887409e-05, 
    5.91212302487645e-06, 2.94745433894158e-05, 1.22507065779909e-05, 
    7.37315183414993e-06, 5.74411514360872e-06, 1.56350823347153e-05, 
    1.40786863467516e-05, 3.5513494022354e-06, 1.32245345503564e-05, 
    8.97434362798695e-06, 6.87584957140117e-05, 7.54699485805367e-09, 
    1.62846523473839e-10, 3.10588883086896e-12, 3.81258832917865e-11, 0, 
    1.36496527153975e-19, 1.92397613814905e-05, 4.1862966960132e-09, 
    2.49029612670357e-05, 5.948939115861e-05, 1.03468465618404e-06, 
    1.05305343764996e-07, 1.4754308104645e-07, 3.88844402994881e-11, 
    1.939302220956e-09, 9.28124642447824e-08, 8.78923001150514e-07, 
    2.4879275008441e-06, 3.60824261808208e-05, 1.7947957412635e-06, 
    4.12394882260678e-06, 3.62661463568211e-09, 4.43047023764793e-11, 
    3.81447685538826e-08, 2.22332640476729e-08, 5.37014086018309e-09, 
    5.33656936014478e-06, 5.72470798038114e-06, 2.16298630067753e-06, 
    1.55106829109356e-05, 4.93152586364326e-05, 8.31409761439498e-05, 
    8.04553869403031e-05, 3.57159823559892e-05, 6.80824172838836e-06, 
    7.21165687372314e-06, 3.97811417883392e-06, 1.42910079865181e-06, 
    6.023272012856e-07, 4.31554445087641e-06, 3.98171742590336e-06, 
    1.0934825493139e-05, 1.15413409451843e-06, 1.28945024149224e-08, 
    1.54722584265683e-06, 7.13788877726401e-06, 8.27971663070003e-06, 
    1.12982650563254e-05, 2.66530951311245e-06,
  3.48658133901987e-06, 6.85229919516103e-06, 9.09672154098113e-05, 
    4.31797347988715e-05, 2.87344023092703e-05, 4.74171026763616e-05, 
    1.94644123588482e-07, 1.68157891322834e-06, 1.71822225134648e-08, 
    1.36021274168868e-08, 6.93765525269072e-10, 8.36908902359607e-18, 
    8.87099613969636e-08, 2.5279903620099e-07, 3.42499852172106e-07, 
    9.02499050640047e-09, 6.58059666655275e-10, 3.20052238384052e-21, 
    4.41595882601619e-21, 4.59383739313568e-11, 2.09453519070301e-10, 
    3.97580836828478e-24, 3.89680340055965e-23, 1.37441910795088e-08, 
    3.8570665251088e-12, 3.97006861126253e-10, 9.72203207771449e-10, 
    3.77611753677841e-11, 0, 0, 2.50659639205111e-09, 7.32032294943861e-05, 
    0.000119591203189423, 3.94596599244527e-05, 9.51349975870961e-08, 
    3.95442519497653e-10, 2.42933129295047e-10, 1.4176326353595e-12, 
    3.41014709721191e-20, 0, 0, 0, 5.61772291850138e-25, 
    2.96715076380434e-24, 4.03164435130938e-23, 7.47702190339157e-20, 
    2.03966363410444e-11, 1.62245295877071e-21, 2.04090375927822e-23, 0, 
    3.49401346979642e-07, 1.11952556986579e-06, 4.41499172971822e-06, 
    0.000118162999319301, 2.59606989973302e-05, 3.31968438679525e-05, 
    3.22668160982632e-05, 4.06907256539074e-05, 8.41979521839982e-05, 
    0.000284383070420946, 0.000391288875448192, 0.000239703027853001, 
    2.90473105345148e-05, 4.89730555502472e-24, 2.45197771890422e-12, 
    4.12541042410104e-12, 2.44749808813193e-10, 2.76825646037999e-10, 
    5.38345861764286e-10, 4.21208020452091e-10, 3.33331924893564e-11, 
    1.8970627287338e-10, 2.02704914121611e-07, 6.01840966818409e-07, 
    1.29627423025439e-07, 2.12200954388099e-07, 1.58402809693543e-06, 
    1.11023872716492e-05, 1.89002865249469e-05, 1.81337674248092e-06, 
    2.30888073868699e-05, 4.06166067672831e-05, 2.92634328890866e-05, 
    4.04123295214663e-05, 1.58928657407181e-05, 2.54968796281348e-05, 
    3.66115980009221e-05, 2.71999855914697e-05, 4.10180777405503e-08, 
    2.29550924067794e-05, 5.77095921923353e-06, 1.0791089470627e-05, 
    7.13475263537129e-06, 6.79972074957226e-06, 4.49454841607022e-07, 
    2.62119127927121e-10, 1.16353546267039e-08, 8.71463420093929e-21, 
    3.62364183859557e-14, 7.71423372656126e-11, 3.47695712339161e-08, 
    1.57520077821195e-05, 6.6093116378716e-08, 7.0875719616197e-09, 
    4.40455237837901e-06, 4.04012775077997e-05, 4.58546748990981e-08, 
    2.10671761408497e-09, 5.87864963253504e-10, 2.77515490074391e-08, 
    3.5083805783855e-07, 4.51099743505519e-07, 1.19366893263099e-07, 
    1.60952214109129e-07, 1.72688690074107e-07, 1.28397664018016e-06, 
    2.94195568893249e-07, 8.73337648593937e-10, 2.43148543475733e-08, 
    3.79952598459462e-08, 1.67531403303807e-09, 3.73021829808479e-11, 
    3.9335650075107e-07, 2.45228969668854e-10, 2.59068832368577e-05, 
    4.4603418678276e-05, 7.83650802978934e-05, 0.000109415850728412, 
    7.63969870238896e-05, 4.10981793405593e-05, 1.41000817373892e-05, 
    9.45331191146844e-06, 1.35326520636513e-05, 1.25240971048889e-05, 
    6.95299343536284e-06, 5.82187641344712e-07, 4.1927110391137e-07, 
    1.2871101847607e-06, 3.96459127941573e-06, 2.96742561612862e-06, 
    1.02676627020877e-05, 1.24058946603938e-05, 7.58019395124123e-06, 
    3.6308767189738e-06,
  3.14792657910741e-06, 2.19634244345467e-06, 1.26079418110311e-05, 
    1.37421303977314e-06, 3.23516804408785e-06, 7.78349854665956e-05, 
    1.86554071786065e-05, 4.76200388886072e-09, 6.73335969887225e-10, 
    1.30504437400036e-10, 7.38704563529852e-11, 2.88829275398895e-10, 
    1.67306611063338e-08, 2.20378700438891e-08, 1.59152159125614e-07, 
    5.39936083972306e-07, 4.00101809571656e-05, 0.000133054925278701, 
    8.47363820866848e-05, 7.04598336864949e-06, 4.84503445029536e-08, 
    1.29982328178417e-10, 1.02392075982431e-10, 2.02254429836216e-12, 
    9.95910697978839e-20, 2.48192203338211e-14, 2.63865890937695e-10, 
    1.42689167090412e-11, 0, 5.81548618490032e-11, 7.60931353546982e-13, 
    9.8397577170242e-05, 0.00030661714548332, 0.000110118289331685, 
    7.25623608333624e-10, 1.63238728625918e-10, 2.21573703405055e-11, 
    3.73708612955349e-10, 1.23050181381254e-20, 2.1282711515792e-05, 
    5.51513314142584e-12, 1.17232100719794e-18, 1.99416322880436e-12, 
    2.84336169905265e-07, 8.49285084776577e-08, 5.72923997452288e-12, 
    1.0298862287003e-24, 2.7206849213074e-07, 4.25573972815511e-06, 
    8.7900011201775e-06, 2.4227304174535e-05, 3.87370743958209e-05, 
    3.10748658916821e-05, 0.000105586440530583, 2.55800329642983e-05, 
    3.47171331931406e-05, 3.52875176584218e-05, 1.49368741535154e-05, 
    1.35459500588024e-07, 5.81784937082016e-08, 6.76144072985185e-09, 0, 
    1.1716478916042e-12, 6.3334607247218e-11, 1.57854610373014e-09, 
    8.63820770788893e-09, 1.12521498504613e-07, 2.24290957961366e-07, 
    3.23183879018042e-07, 3.67504873683485e-07, 1.79512217020745e-07, 
    1.87482980833174e-08, 4.08081056767061e-08, 3.99364496596543e-11, 
    2.19744686476075e-15, 3.36605778456062e-11, 9.08397726160923e-11, 
    4.15899783378386e-11, 1.15512017646882e-05, 1.90432584429041e-05, 
    1.35955415205372e-05, 2.2624425922515e-05, 2.99174366245782e-05, 
    3.45659494644601e-05, 5.16391374555357e-05, 6.3886532114956e-05, 
    6.88036776328401e-05, 0.000135288992951608, 5.2605428132756e-05, 
    7.31494629021764e-05, 6.64940723101532e-05, 4.02305941087773e-05, 
    3.53162715062374e-06, 1.958551208766e-05, 3.1200418102714e-08, 
    1.19525667188218e-10, 9.42420925833434e-21, 6.44015915579674e-10, 
    5.54994152857335e-10, 6.58353049465474e-12, 2.26345633070361e-07, 0, 
    1.16680894788373e-09, 3.81472153353289e-11, 7.22651970503626e-06, 
    7.04660960919463e-05, 2.6906361623621e-07, 4.78846956524927e-09, 
    1.80445178097964e-11, 7.72809064040691e-10, 2.37975851246674e-07, 
    4.27457090663036e-07, 4.22173901799721e-06, 2.15750186117137e-06, 
    6.43687061561834e-07, 6.008134633874e-07, 1.33295052904433e-06, 
    2.08215650603037e-06, 3.9985565168742e-07, 1.45629596198894e-06, 
    1.97572769382675e-07, 2.23137666342189e-07, 7.30045623102192e-10, 
    1.61094170525673e-08, 2.29257007635876e-07, 0, 0, 0, 
    3.11392335642965e-06, 6.21921568068489e-06, 2.01235696151521e-06, 
    5.55801261395902e-07, 1.97206804550038e-06, 5.05850785550139e-07, 
    3.09848449961676e-07, 7.93812783888036e-07, 7.27083853511746e-07, 
    4.36053844426847e-11, 1.12800104075177e-09, 4.02715207065617e-07, 
    3.96384553302204e-06, 4.65755028799753e-06, 8.6438843983095e-06, 
    1.19140806920848e-05,
  5.46658209075642e-06, 4.26669008441941e-06, 9.46646971869749e-06, 
    1.62634965016019e-05, 1.56783301285619e-05, 1.35668545199753e-11, 
    3.09585803081526e-05, 6.07305004184511e-08, 1.00110447479171e-08, 
    4.42960505210462e-08, 1.63767607654113e-08, 2.00686800175523e-10, 
    3.39772076628024e-11, 3.35354069736779e-09, 2.83443208809886e-05, 
    9.3477899808895e-05, 9.8382569851002e-05, 0.000205293011882791, 
    0.000186362838010834, 7.21301343683024e-05, 1.77030448770136e-06, 
    1.48433954456715e-09, 3.17141878498131e-09, 9.16453387221995e-14, 
    5.06238144889668e-11, 1.16535079976632e-07, 4.11519859286991e-07, 
    1.86511164418413e-09, 2.7438096981125e-20, 7.933870058183e-21, 
    1.53681263007626e-14, 4.92663204105421e-07, 0.000343347079429502, 
    0.000292550524639128, 9.80395011927039e-09, 1.49073903136963e-08, 
    1.72116651665879e-08, 2.76356518020874e-09, 1.31769886648513e-17, 
    4.26086918691114e-07, 8.76341870646949e-10, 3.55344929974569e-37, 
    3.91385430451684e-19, 0, 1.92485750604724e-20, 5.5375717443339e-16, 0, 
    1.40974601936649e-11, 2.0174075277757e-10, 2.01167208362579e-07, 
    2.97664179665876e-05, 2.09385842697213e-06, 5.45028735989125e-06, 
    4.25909822207703e-06, 1.87632118780075e-06, 2.75000294174588e-07, 
    3.46850979557017e-07, 2.68109357134934e-07, 1.12428524209373e-07, 
    1.07367726894331e-11, 9.10708667560049e-14, 2.33181110671759e-11, 
    2.74793651598181e-10, 3.43586909555319e-09, 9.07712662084841e-08, 
    6.8657571410873e-08, 7.54486107816486e-07, 5.84709579738655e-07, 
    9.21794094588256e-07, 7.47855430936244e-07, 1.68696162693711e-07, 
    2.26726972309254e-08, 7.3976598073859e-07, 6.79159554316453e-08, 
    8.17312896343491e-09, 2.22867089103598e-09, 5.10869813871216e-19, 
    1.80173625897389e-08, 9.94975336105031e-06, 1.07845076632009e-05, 
    8.09827893396795e-06, 2.00931400743026e-05, 3.3925511349529e-05, 
    5.15529165636693e-05, 7.00238062003087e-05, 5.48844800498449e-05, 
    0.000127340293432734, 0.00012288692330142, 8.62929822200855e-05, 
    5.37198620239434e-05, 1.96329717621692e-05, 2.84779532357508e-05, 
    2.28073547676438e-05, 1.20523982966247e-06, 5.26689099134525e-06, 
    1.51865927431454e-06, 2.0592993811041e-05, 1.58437137151341e-09, 
    2.07038319279523e-06, 1.10956862539783e-06, 1.59313908346958e-07, 
    3.19775144138379e-08, 1.54400333917253e-09, 1.61513495351716e-11, 
    1.85208940853707e-06, 6.09661657818212e-05, 9.29693337401319e-07, 
    6.86445612532732e-06, 3.41172649122578e-06, 3.65846795754272e-05, 
    6.17837063876468e-06, 9.66247081344846e-07, 9.04139157116245e-07, 
    7.06825179359848e-06, 1.68944402602835e-06, 1.43897172580951e-06, 
    7.55539803346688e-08, 8.36755652445704e-08, 2.50504989271873e-08, 
    5.39113977784383e-08, 1.58628356644394e-06, 3.42422096568204e-06, 
    7.90697670287469e-08, 1.84591543020919e-08, 5.88839878596234e-10, 0, 
    7.0779767682745e-12, 0, 1.24007051201611e-09, 0, 5.66425191494303e-07, 
    5.16430210569578e-06, 4.73703221861627e-06, 8.00015623403027e-08, 
    3.86603992165127e-09, 8.9741015859491e-09, 8.31801018323598e-09, 
    1.89060184838112e-09, 9.39867895963468e-12, 6.33851874479286e-09, 
    7.01429191431578e-07, 5.07181276506039e-06, 2.55908602272306e-06, 
    6.96971527452644e-06,
  6.83761372900598e-06, 9.02693974109408e-06, 4.16713471179835e-06, 
    3.49680206183306e-06, 1.29954739190978e-05, 1.17149639419154e-05, 
    1.41174815230148e-06, 2.92303057352499e-06, 1.21778480752981e-05, 
    5.44169611337758e-05, 0.000128916711312486, 0.00015599350783627, 
    0.00013451681872919, 0.000117649591707018, 2.31268262262981e-05, 
    6.66194109012268e-05, 0.000121758949319801, 9.81750919962107e-05, 
    4.37979591880132e-05, 9.95347772549068e-07, 1.91595831349214e-10, 
    2.03945488922041e-07, 5.32447712968825e-11, 2.42644622640342e-09, 
    2.06824182523963e-07, 1.61030743159363e-06, 2.8740760789355e-06, 
    2.26018862002634e-08, 3.94068780902412e-10, 3.986181140522e-11, 
    4.15508016780946e-22, 1.22697042521769e-08, 3.64337401387564e-05, 
    0.000278051397165234, 3.84566171597509e-05, 3.16376016093914e-08, 
    1.59790338432189e-08, 1.56478915028398e-09, 5.95569808650272e-17, 
    1.15312738260831e-17, 4.54715598410525e-17, 0, 0, 0, 0, 
    5.60062616754451e-18, 2.03980666369373e-16, 1.9743972697572e-21, 
    3.78517655244465e-15, 9.35927690496115e-16, 3.1617949290158e-09, 
    1.36498536494996e-07, 3.04427638115515e-07, 3.20595437577155e-08, 
    9.83020242699962e-23, 3.98699488514839e-17, 0, 0, 0, 3.9203367890466e-12, 
    6.24891864072373e-11, 1.43135268050071e-09, 3.84630328867821e-08, 
    4.72770003992294e-08, 2.58609115595547e-06, 2.53946234186918e-06, 
    3.21878655350013e-06, 4.72198569965841e-06, 9.15467555832456e-06, 
    1.22276330839212e-05, 9.72207537842591e-06, 5.44616764692587e-06, 
    2.85611091085889e-07, 8.7133861254725e-09, 6.41125395216335e-07, 
    2.11946103788835e-07, 1.40837526503422e-10, 8.93410249411238e-09, 
    2.04535121480844e-06, 1.65808871997099e-05, 5.12149750033447e-05, 
    1.51478096655275e-05, 2.06133032633182e-05, 1.07764425170734e-05, 
    7.67010947585902e-06, 7.14779313178863e-06, 5.82831318867787e-05, 
    9.89201944072688e-05, 0.00012406095842286, 4.11062563493284e-05, 
    5.08988065827348e-05, 6.09150063474668e-05, 4.2471166008832e-05, 
    4.67846446348191e-05, 5.09504176056103e-05, 4.38686361896627e-05, 
    4.85396495921105e-05, 1.25559541239112e-05, 8.59242616009672e-05, 
    6.45258149066746e-07, 1.65340436594523e-07, 0, 3.17285991567445e-11, 
    3.38472665719725e-10, 1.56604576336062e-18, 7.20261130615085e-05, 
    2.50873520210385e-05, 1.33518779319944e-06, 2.66586426196628e-05, 
    3.43387067279006e-05, 4.58870015508188e-06, 2.52810298311483e-09, 
    6.25741793030236e-07, 1.10505047058785e-06, 2.67049610041119e-06, 
    5.76918668939121e-08, 2.41833345994584e-10, 2.7021809324967e-12, 
    7.80140614480222e-11, 1.49890135573635e-11, 5.85093156203523e-07, 
    1.7994190648381e-06, 1.55539416404197e-06, 6.56978079830452e-17, 0, 0, 0, 
    0, 6.30337004402862e-11, 5.54083079038442e-09, 0, 0, 
    4.11628625504118e-11, 0, 5.74399883997191e-09, 1.48052508319522e-08, 
    6.62384905464581e-08, 9.3138320736334e-08, 5.30652622271995e-08, 
    1.32174706982394e-08, 3.0619647871931e-06, 6.95537656279862e-06, 
    6.45145041806955e-06, 8.52572274018239e-06,
  9.90952095239631e-06, 6.54568257232674e-06, 1.99466789179577e-06, 
    1.07272999936892e-08, 2.00479555634024e-06, 1.77218331854235e-06, 
    1.4799718570381e-05, 4.69369331178984e-05, 8.97675387719308e-05, 
    0.000168657096555134, 0.000269423528595714, 0.000341360136490718, 
    0.000309653762803721, 0.00021680962766355, 8.71664199730216e-05, 
    3.66362221640629e-06, 2.7716030522131e-07, 5.58713653825015e-07, 
    1.48333865800642e-06, 9.3709621740795e-07, 3.29694905514308e-06, 0, 0, 
    2.05008353485781e-06, 2.16628364281134e-06, 5.20884404804247e-06, 
    5.36093557109977e-06, 3.77850644691222e-06, 7.74263972976041e-06, 
    7.93154365406986e-07, 1.01805274398544e-10, 6.89739524447652e-10, 
    3.69707536446147e-10, 5.27552994564753e-07, 0.000109463828110862, 
    3.95333030660507e-06, 2.92406134049027e-07, 2.41476536918592e-10, 
    2.83525418325207e-11, 2.09128984279623e-10, 5.64674460062887e-20, 0, 0, 
    0, 0, 0, 5.07789114214996e-17, 5.44719300732592e-25, 0, 0, 0, 0, 0, 
    4.31851510817365e-15, 1.19849876319045e-11, 1.86674462287943e-23, 
    6.12913521063649e-24, 4.64714592327775e-24, 0, 9.21826174377693e-11, 
    1.05473782098108e-09, 1.55424516624533e-08, 3.36285462675922e-08, 
    2.73846730695479e-07, 4.16056123857805e-09, 1.79452152630352e-07, 
    4.42771603889278e-09, 3.10113015856079e-06, 3.00300501498509e-05, 
    5.97490576078509e-05, 5.62466109808995e-05, 3.47136626566813e-05, 
    2.57743917075049e-05, 1.8485592422382e-05, 4.19678978543306e-06, 
    1.05693978525153e-07, 8.70465892326819e-09, 2.35038209672952e-11, 
    3.06065200545355e-08, 2.81622343634166e-06, 9.59762206957026e-06, 
    8.70298095921324e-06, 7.12197411540962e-06, 7.68756832810535e-06, 
    5.39235482728893e-06, 2.64237536989738e-05, 1.69433585814117e-05, 
    6.75591792327666e-05, 1.54375830770874e-05, 1.64384414277422e-06, 
    2.21721752328226e-05, 3.42326421465868e-05, 4.36278748351213e-05, 
    7.79470446980074e-05, 5.88094517023049e-05, 5.65954451537854e-05, 
    4.03992082331462e-05, 9.89461541799821e-06, 1.77573049856881e-05, 
    6.39037687258383e-20, 8.77823818681925e-23, 1.04631646210108e-09, 
    4.82465931979371e-12, 1.43613238419448e-10, 8.96540563918047e-07, 
    4.09558879025521e-05, 2.97326499521481e-05, 7.7334343090735e-10, 
    9.59338035558159e-07, 4.57245130338845e-07, 4.86328376333769e-07, 
    9.0594632192939e-10, 1.49542277687243e-08, 1.0948625300987e-08, 
    5.00716928223746e-08, 3.06211014138171e-10, 0, 7.26625800020863e-12, 
    5.29671618326315e-10, 9.48609556392381e-09, 1.31796460614931e-06, 
    3.19030407432749e-07, 4.03094031351084e-09, 0, 0, 0, 0, 0, 0, 0, 0, 
    7.18291340788076e-12, 0, 0, 8.09539166059592e-18, 5.56024026462429e-11, 
    5.04992322156681e-10, 1.0343034908289e-09, 1.04499183472308e-09, 
    3.8205075931562e-08, 6.05231200912237e-06, 8.21262189097853e-06, 
    7.78297892267506e-06, 7.11442904070625e-06,
  7.94482964687799e-06, 1.05818595807025e-05, 6.92721434122127e-06, 
    2.20304180729355e-06, 2.57163754047482e-06, 2.54720673709667e-06, 
    1.4626680836016e-06, 3.11849816725706e-07, 4.76415351672581e-06, 
    3.19419422364956e-06, 8.50994110449046e-06, 3.98078146431402e-06, 
    3.41230903223218e-06, 1.82472166572016e-06, 1.66046183622392e-06, 
    1.68513710248926e-06, 2.92425567461385e-06, 2.90682472446885e-06, 
    9.93387632651175e-09, 2.34311914746303e-06, 1.49565572456986e-08, 0, 0, 
    0, 1.1233865711196e-07, 9.08754607188715e-10, 1.09163757004061e-06, 
    3.57480896840007e-06, 5.08092762275264e-06, 5.58742294457342e-06, 
    8.30823754145843e-08, 7.93150910284947e-17, 2.00799761671271e-12, 
    1.15173410991344e-09, 5.70694442579523e-13, 2.13873827130347e-05, 
    1.10766145036568e-05, 1.01727770151948e-11, 1.24752905814094e-08, 
    6.96790533701946e-09, 0, 1.78723765235809e-16, 2.1706684747668e-19, 
    3.49414343931143e-19, 5.99156163380456e-21, 9.41305835561574e-17, 
    1.07266512855603e-16, 4.95638194246643e-19, 3.92709824582086e-20, 0, 0, 
    0, 9.05249706172829e-19, 9.65695113306282e-24, 2.71633906497413e-21, 0, 
    0, 1.9972044419903e-23, 1.66753961119714e-21, 1.52569655225161e-10, 
    1.99668073224272e-08, 6.99589349645846e-08, 2.83348346605748e-07, 
    5.40347338257353e-07, 2.23855105478424e-07, 2.39269971584674e-06, 
    3.97686261083654e-06, 2.43609290280745e-06, 4.38284872234243e-06, 
    2.73449777315838e-05, 2.22371383121796e-05, 1.33999104088985e-05, 
    2.78414674586035e-06, 2.01094982576771e-06, 7.80316815227718e-07, 
    9.53584628572494e-07, 9.35976956796647e-07, 4.12040874930795e-07, 
    3.42984276851155e-07, 1.67634342039268e-07, 1.39995425518102e-08, 
    9.79796964782955e-10, 3.61941234199731e-09, 4.124003424252e-08, 
    1.24434315670388e-08, 6.62316507197787e-09, 2.69762414283889e-10, 
    4.72833054405513e-21, 1.80686438427712e-17, 1.67818750136844e-16, 
    8.39047508406157e-23, 2.02004081001519e-07, 7.06155319483982e-06, 
    1.13517225858135e-05, 7.42746016498763e-05, 4.02659900278179e-05, 
    3.28039313878301e-06, 1.7178983481314e-06, 8.78343050635543e-10, 
    2.46153823834044e-08, 9.40001637750774e-09, 1.16060082791725e-11, 0, 
    1.66480449911538e-10, 3.21216789812618e-08, 2.03461800661196e-07, 
    1.56034311425528e-10, 1.26302250583631e-10, 1.60502676341578e-10, 
    2.23469766351947e-09, 1.93693562406005e-08, 1.13129808650407e-10, 
    1.50707185287476e-09, 2.85316021537389e-10, 1.09086015398882e-19, 
    1.2431606187911e-19, 5.19525013166613e-11, 4.05277900169682e-10, 
    4.18629993503129e-08, 1.34029823238306e-06, 4.02126229609908e-06, 
    2.59311513228615e-07, 3.34233768514126e-10, 0, 0, 0, 0, 0, 0, 0, 
    7.03137017351673e-12, 0, 0, 0, 0, 7.2837663314416e-18, 
    1.20088320653985e-09, 3.03648080191461e-08, 1.04018187455177e-06, 
    4.30790852529628e-06, 5.01572406474352e-06, 5.04062203384408e-06, 
    8.81435105550319e-06, 6.4707826036567e-06,
  4.48823871878553e-06, 4.25699673189664e-06, 7.36248335092801e-06, 
    5.16909544278691e-06, 9.24734538669174e-07, 4.63386777589027e-08, 
    4.36772452030676e-07, 3.28849802295743e-07, 2.42367072226454e-07, 
    3.17022582257407e-07, 1.07824587433959e-06, 8.15991225583306e-07, 
    2.18007115759142e-06, 5.31498236759083e-07, 2.36454805265477e-10, 
    7.32841820732862e-10, 0, 0, 2.58436616581087e-11, 0, 0, 0, 0, 0, 0, 0, 
    1.36033993318203e-06, 1.29656015454819e-07, 7.48456436649949e-07, 
    2.11972159274586e-07, 7.70512360154971e-08, 4.82185088959828e-09, 
    2.25361830330645e-10, 2.98815265796528e-07, 7.77220451571552e-07, 
    9.69630404546927e-09, 2.47090945739556e-08, 6.35492377389522e-06, 
    1.13584184586149e-05, 5.83658058479216e-08, 9.34211178782244e-08, 
    1.35114469452173e-10, 6.45872182343128e-11, 5.33587794795176e-11, 
    3.58186636320865e-11, 1.10903502222241e-10, 8.98694531152436e-10, 
    4.13344310340219e-10, 1.60515832236383e-11, 0, 2.80004247750974e-12, 
    2.35484024103376e-17, 2.16356425509119e-11, 3.66982213694095e-12, 
    4.8974087933712e-14, 0, 0, 0, 3.20635078671608e-25, 3.71131390455224e-11, 
    2.40716046181344e-09, 2.12645266345235e-08, 1.9009109913049e-12, 
    1.04901152908355e-07, 7.17086978928141e-08, 6.07539774970581e-08, 
    7.61013980707175e-07, 1.89315721857348e-06, 1.53786648635789e-06, 
    3.88338163793464e-07, 1.15074778493399e-06, 1.09674133343985e-07, 
    9.38530488403343e-08, 1.05738755989212e-09, 1.41443559488513e-08, 
    4.51563794938897e-08, 5.56865178592206e-08, 5.46461522429875e-08, 
    3.51049019321285e-08, 1.93694437004014e-08, 1.10817681631257e-18, 
    3.93168759775055e-11, 2.85138799971227e-11, 6.05950753872551e-11, 
    1.10129998013261e-11, 1.66714532038677e-10, 1.97339332300748e-11, 
    1.5593924237862e-07, 4.26636950021627e-06, 1.94327721413691e-05, 
    1.75195306760444e-05, 1.05637658027632e-05, 4.83026610452284e-06, 
    4.89844334494397e-05, 1.51426461452056e-05, 6.31442535853452e-10, 
    2.59373324081161e-25, 2.72689529232228e-23, 1.74552390845823e-19, 
    1.09889534964255e-22, 6.64509237713057e-17, 0, 0, 4.51026108051466e-15, 
    7.25409440982313e-10, 3.11123216598768e-08, 0, 1.94656509658127e-25, 
    3.17182974462803e-08, 2.16192518647992e-10, 8.50503825761461e-10, 
    1.37146179768348e-10, 3.18104697370757e-08, 1.65059707887871e-06, 
    2.99195168073111e-06, 2.29320244378274e-06, 3.27084092615083e-06, 
    3.25888219520128e-06, 2.86199840994035e-06, 9.68798850786339e-07, 
    1.39917703584854e-07, 3.10855649414214e-09, 1.21952798336501e-19, 0, 
    2.58599801935055e-20, 0, 0, 0, 0, 0, 5.02080389415882e-09, 
    2.28332300578961e-11, 0, 0, 0, 2.70415706485787e-19, 
    3.77413937183131e-11, 1.30210755750138e-09, 1.1260169591193e-08, 
    1.14899608197013e-09, 9.19042582262238e-08, 1.0177921180622e-06, 
    3.57288039116778e-06, 4.53662317698875e-06,
  7.84324421214815e-06, 6.47351465985394e-06, 5.63856181549398e-06, 
    1.07897378084321e-05, 2.35945041376735e-06, 3.97410066820352e-07, 
    4.6038162270231e-10, 9.42085488305693e-12, 1.25103243202131e-10, 
    2.16668943632856e-11, 3.24461791718072e-13, 1.24925431291318e-10, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.85840395116424e-06, 1.20342531264996e-06, 1.22817763446159e-06, 
    1.23028506759077e-06, 3.61276791625726e-06, 2.0562529138517e-06, 
    4.20059149235234e-06, 1.30124800703512e-06, 2.59561856297057e-06, 
    8.9179349321661e-10, 3.31241857535888e-09, 6.75117677189427e-09, 
    9.42280302499015e-09, 5.75929101743565e-09, 1.33784411915477e-07, 
    1.81848218583696e-07, 1.14483297823177e-07, 1.6789162359316e-09, 
    3.15851490729335e-10, 1.97946100749394e-10, 4.11119744094914e-09, 
    1.67600136730161e-11, 4.36283403856359e-11, 0, 0, 0, 0, 0, 
    2.45007807878877e-08, 2.40872625934154e-05, 3.83854354295185e-05, 
    3.32741795379467e-05, 9.45206868207071e-08, 4.33918793126006e-06, 
    3.77543840219439e-08, 1.0628716380262e-06, 5.20776033797687e-07, 
    3.69802428074346e-07, 3.03447685189688e-07, 2.98736043736922e-07, 
    5.56954706060778e-12, 1.74374091131095e-13, 9.08410634039723e-10, 
    1.04341916951086e-10, 5.37325016225859e-11, 2.11960590002637e-11, 
    3.71559209768771e-09, 4.63061092775752e-12, 5.59162334449801e-11, 
    7.88527057068838e-12, 8.90731305278729e-13, 6.90240364727005e-19, 
    3.25015618953588e-07, 5.24246211485717e-06, 6.50036926233511e-06, 
    4.83598000843489e-06, 3.52967476019809e-06, 3.03855775045551e-06, 
    2.32925530955756e-06, 1.14170321820151e-06, 3.0610816808154e-08, 
    6.68786844086064e-17, 3.99788733993233e-15, 3.59278164660044e-10, 0, 
    9.87625477871923e-23, 5.90043352253548e-20, 1.48232873629775e-24, 0, 0, 
    0, 0, 2.54744914492937e-22, 0, 4.91215462622722e-18, 0, 
    9.6026836164417e-12, 8.75356694425673e-11, 2.81621638185804e-09, 
    6.97287199946878e-20, 2.14512763213096e-07, 8.17804582170856e-07, 
    1.07997954905727e-06, 1.06355842465781e-06, 4.42346240023882e-07, 
    1.12217759964993e-06, 1.27570359437041e-07, 4.07886322746445e-09, 
    2.10211072676731e-09, 2.14572019251141e-12, 1.26343091976868e-18, 
    1.79383486203778e-11, 8.44139028796295e-12, 0, 0, 0, 
    3.60752042412932e-10, 0, 0, 0, 0, 0, 0, 0, 4.06576305849195e-16, 
    1.08241930353405e-11, 1.57633142923695e-10, 1.30865891933864e-10, 
    1.08978574412403e-09, 1.76441055011173e-09, 1.99773905220019e-06, 0,
  4.73253455768324e-06, 6.70232710092965e-07, 1.51449533982468e-06, 0, 0, 
    9.38732144432759e-11, 1.02988862038066e-11, 8.70000225163446e-12, 
    6.23629098444684e-11, 2.03935159818783e-11, 7.6121604185994e-12, 
    7.946394273504e-12, 0, 0, 8.0642993805713e-07, 2.34574331766495e-06, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.25846872228423e-07, 
    2.46836620376924e-06, 0, 0, 0, 8.64941021048804e-10, 0, 
    3.59458918091861e-07, 4.34476150230221e-08, 0, 0, 0, 
    7.54667989295789e-07, 9.19366865012041e-07, 0, 8.73882205247058e-09, 
    2.14288440428758e-07, 2.62802451108485e-08, 6.16767337905143e-08, 
    1.42038011300614e-07, 3.71143612646309e-07, 4.13718169137205e-07, 
    9.7106891777901e-08, 2.86993553380598e-12, 2.3100903137508e-10, 
    3.50665636445777e-10, 0, 0, 0, 8.60881687150075e-26, 
    4.35464599205989e-14, 3.72775718324358e-06, 3.0568661468822e-06, 
    3.4494510969196e-05, 8.15112683660113e-06, 1.45015017659148e-06, 
    2.50914402259133e-06, 1.48618479852106e-06, 5.96426659072838e-07, 
    1.53045348828011e-08, 7.97822277015046e-09, 3.03882914252759e-08, 
    2.23813738053334e-09, 6.14447112696778e-13, 1.32657973927094e-10, 
    8.01751346553484e-12, 1.3946357016032e-09, 3.44256774144038e-08, 
    3.20920914660814e-13, 1.14077724626332e-13, 2.21031550955363e-23, 
    1.45316299390211e-23, 9.68241690198127e-20, 5.31533235625236e-21, 
    9.07106528029065e-09, 7.21242755494708e-09, 5.18752167496719e-09, 
    3.8414358754133e-10, 1.87492107455726e-10, 0, 9.96761211560965e-09, 
    4.10430787170469e-09, 0, 0, 2.7491823649997e-17, 8.72976223410606e-12, 
    1.72728464513733e-13, 1.0803708126117e-13, 0, 0, 0, 0, 0, 0, 0, 0, 
    3.40238768209862e-21, 0, 2.95765113312303e-11, 5.73383194219492e-10, 
    3.78808403380401e-17, 1.15716940506607e-08, 4.83703058589539e-08, 
    1.81839721501218e-08, 5.87374515404925e-09, 1.11323141636169e-09, 
    6.81921090935728e-09, 2.11821428562345e-09, 1.73041133996367e-10, 
    1.46503116009825e-12, 0, 0, 0, 0, 0, 0, 0, 0, 3.07352125491256e-11, 
    1.01744144869604e-10, 2.34823896235933e-10, 0, 0, 1.69017587852181e-12, 
    1.42534408958065e-10, 5.36118398747486e-10, 3.79881888813544e-10, 
    3.04965280208336e-09, 4.76329294165419e-10, 7.13189647650617e-11, 
    4.00713947591205e-10, 2.25376930309519e-06, 8.44406497905465e-06,
  5.53937099871576e-06, 1.72241789550133e-06, 3.68196453994309e-07, 
    9.26314510569164e-07, 0, 0, 0, 0, 1.0367692117103e-10, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1.89979236792779e-06, 1.80887060224243e-06, 3.78173442794504e-07, 
    1.95366965773902e-08, 6.53326294109382e-09, 1.33480501244356e-09, 
    1.26917571106978e-09, 2.80727417601165e-08, 1.43889770240357e-07, 
    6.62960857401438e-07, 1.75964079634619e-06, 0, 2.05546688724583e-08, 
    4.16995484388376e-07, 8.60375796710827e-07, 2.00047413387041e-07, 
    9.0896968012013e-08, 1.0983339220182e-08, 6.07569668055212e-11, 
    2.74755150286832e-25, 4.24058063124863e-24, 9.10100975920425e-07, 
    1.11968714845349e-06, 5.6832685110809e-06, 1.40713852659238e-06, 
    3.91863384927253e-06, 1.04975293209647e-05, 2.60721057239358e-06, 
    1.29300013042921e-08, 1.83790447131982e-06, 5.11963512920361e-10, 
    9.52008417094291e-08, 3.54695377807458e-09, 1.47045035344184e-08, 
    2.64746180866908e-09, 1.66937819050533e-18, 4.01123940321364e-18, 
    1.56706275296917e-22, 0, 0, 0, 0, 0, 0, 3.9319753228471e-18, 
    5.39755160275861e-18, 0, 2.6210111295403e-22, 0, 3.26997403258497e-12, 
    2.55860081969703e-23, 1.19553874560592e-17, 3.94750474645037e-20, 
    1.28919763847178e-17, 1.6914956870684e-19, 2.99547808259082e-23, 
    1.20086509891213e-21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.8549284327652e-11, 
    4.38079086398799e-10, 4.27640526540119e-09, 2.31467400913789e-11, 
    1.54455137642739e-19, 1.49734473921377e-09, 1.12770162595335e-10, 
    6.91827049052517e-10, 2.37147350587802e-11, 3.27203139639224e-10, 
    5.05796873371607e-09, 4.24933312474542e-10, 6.55597020088952e-11, 
    2.73044668660442e-12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.70465404254939e-24, 
    2.81983083773681e-11, 2.26949711747813e-10, 1.15478977585409e-19, 
    4.02175133035734e-09, 7.45879305820739e-09, 9.02202749508973e-09, 
    2.37584697379806e-12, 9.30426914617711e-09, 3.35611801978357e-10, 
    5.66475934350862e-10, 7.40813597906665e-08, 8.59491446693361e-07, 
    2.86075564119528e-06, 4.71221175888781e-06,
  5.86309157288254e-06, 5.7849760377578e-06, 8.36035439732266e-06, 
    7.60789724821144e-06, 4.6203649770551e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3.98346247411701e-06, 2.46353828024539e-06, 1.4388413455606e-06, 
    2.1915681703319e-06, 3.09391299559918e-06, 4.13983553963611e-06, 
    3.46775000604553e-06, 2.07991917138669e-06, 6.09748948578318e-07, 
    4.67311107305165e-07, 6.15245110108357e-07, 1.03593859731181e-06, 
    1.32402148008752e-06, 1.14837115814627e-06, 6.33137902757438e-07, 
    5.779727170547e-07, 1.01975876410911e-06, 1.53970560112911e-06, 
    1.61246965393285e-06, 2.34419708584667e-07, 3.90057780365212e-08, 
    5.8701793789282e-09, 2.24047487956567e-08, 1.56377525034378e-07, 
    6.70799571633578e-07, 1.93571469224683e-06, 0, 0, 0, 
    2.76592739678557e-06, 5.03561916778372e-05, 7.1399512685441e-06, 
    4.70680535246267e-07, 6.31254110660303e-07, 1.58662627487225e-13, 
    8.51196847060098e-17, 8.00856520448788e-09, 5.15470874075863e-07, 
    6.93505175614493e-08, 1.54337859712178e-07, 1.91069105134121e-10, 
    7.06260159166687e-12, 0, 9.72617257148625e-14, 0, 0, 3.6134563264941e-11, 
    0, 0, 0, 1.52684307928854e-08, 5.00088018931927e-11, 
    1.23824365416398e-17, 3.65710278636847e-21, 9.11781842688346e-22, 
    6.48681683194014e-18, 0, 2.28451496318845e-18, 0, 0, 
    8.58889297578977e-21, 1.56413564615197e-23, 3.73043619196666e-17, 
    1.72944216214558e-18, 0, 0, 1.14953300836707e-18, 0, 0, 
    1.43740076433268e-11, 4.36001703111088e-10, 5.35812348447159e-09, 
    1.16877028174227e-08, 0, 0, 3.84103999959876e-18, 1.11901054173809e-18, 
    7.30973116843696e-08, 7.30979648106687e-08, 3.7553617079639e-08, 
    5.87593818959419e-09, 8.01499829800373e-10, 8.69664145140657e-11, 
    4.34220513087687e-09, 1.73109435187936e-21, 6.53986645666218e-21, 
    3.78220298861198e-22, 5.46836450119027e-11, 0, 0, 5.99424586998337e-25, 
    1.76399510813903e-21, 1.39674848148565e-12, 8.45885186228108e-09, 
    8.53089214349161e-09, 9.3219137955294e-11, 7.67768297316681e-11, 
    2.31526685764632e-08, 1.45511764289434e-07, 3.71493314054539e-07, 
    4.58893143967647e-07, 7.93549117931599e-07, 9.8460379290312e-07, 
    1.31993761608544e-06, 1.14078107420776e-06, 1.90111681744252e-06, 
    4.82360774491628e-06,
  5.1669656955627e-07, 7.47219348624612e-07, 1.62701656614095e-06, 
    2.59278737947299e-06, 2.76970611996587e-06, 3.10207640577511e-06, 
    2.61822592532095e-06, 5.11436733289339e-06, 3.30895278331554e-06, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1.34476580442528e-06, 3.63968584460466e-06, 
    8.09688940390112e-06, 7.04725158185479e-06, 6.07677981545671e-06, 
    4.62417900003901e-06, 5.60477184562511e-06, 5.80690952035983e-06, 
    4.177805298617e-06, 2.95442792472946e-06, 4.32675181198278e-06, 
    3.1019984838506e-06, 2.74044427605754e-06, 1.92497042501556e-06, 
    1.67325126139063e-06, 2.69431848155298e-06, 8.75568770359376e-07, 
    2.68353074690154e-06, 2.94339104544553e-07, 0, 0, 0, 0, 0, 
    1.30236102198209e-06, 1.12288238940552e-08, 1.87537769431715e-05, 
    6.9373215443033e-07, 2.36628189269179e-07, 1.30150521199966e-07, 
    1.02581697014393e-16, 2.6122033663847e-07, 2.6302093639328e-06, 
    8.76699097147653e-06, 2.40491669314303e-05, 4.2104719271324e-05, 
    4.82512224808259e-05, 4.50855200595578e-05, 3.77999943287298e-05, 
    2.63059256783393e-05, 1.5410865257386e-05, 5.73574862605591e-06, 
    8.21003466184352e-07, 0, 0, 0, 0, 0, 1.75245585527211e-20, 
    1.1147730707313e-19, 0, 3.39184337089513e-23, 1.12925507584136e-19, 
    4.17484172348242e-09, 7.94545449986342e-19, 1.02430108888221e-19, 
    1.89989624387204e-22, 1.19276491211927e-20, 0, 0, 0, 0, 0, 0, 
    1.41351565057608e-17, 2.33787678739733e-09, 2.48976782272685e-09, 
    5.61075485305489e-09, 2.20386134605259e-08, 4.00076996543847e-08, 
    4.59988206992596e-08, 4.13341390722547e-08, 7.86062192050199e-10, 
    2.63321443586543e-09, 9.02776896237219e-09, 2.53074254802853e-08, 
    3.25759698884961e-09, 1.98969948726633e-18, 4.00520046195739e-22, 
    1.91082908436524e-10, 3.35724209341869e-10, 2.6636770446103e-20, 
    3.33748102817324e-10, 4.17101105887544e-17, 1.43208455537074e-08, 
    8.01713780653764e-11, 6.58963590354728e-23, 2.05737073817543e-20, 
    1.8685745128055e-12, 4.72060905469184e-11, 4.7930406508358e-08, 
    3.58994514026132e-07, 5.8241543649509e-07, 8.11815882693239e-07, 
    5.85058121001939e-07, 7.11672704788316e-07, 3.99336644042829e-07, 
    4.55543922033409e-07, 3.99083921031506e-07, 4.61569556011025e-07, 
    3.95199926556369e-07, 4.6899687365473e-07,
  2.6892214769164e-07, 2.50508328950353e-07, 4.88260504531944e-07, 
    1.26923738627642e-06, 3.0719367321513e-06, 6.21310472439664e-06, 
    8.71933005284622e-06, 1.20978089610913e-05, 6.50142105395912e-06, 0, 0, 
    0, 0, 0, 0, 0, 0, 5.51199128128882e-06, 4.54561993869871e-06, 0, 
    7.94928975369533e-06, 3.60038385694625e-06, 0, 1.68408187744971e-06, 
    8.91933053664929e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.48299615203571e-06, 3.70984508464277e-06, 5.69483476116206e-06, 
    8.87568702952781e-06, 2.38245056862875e-05, 4.91986735252894e-06, 
    1.77413024296454e-06, 6.40993904589349e-07, 7.6162261982876e-07, 
    5.12765155069173e-06, 1.07007528565034e-05, 1.75330705808738e-05, 
    2.95011505534274e-05, 4.63013204515993e-05, 5.71585136716022e-05, 
    6.63909976057335e-05, 8.01948059771796e-05, 8.54091599495557e-05, 
    8.94818113777771e-05, 8.56866019307901e-05, 7.78495208229767e-05, 
    6.89290801180222e-05, 6.01901382464884e-05, 5.13131735327362e-05, 
    4.2315233952703e-05, 3.3632650434652e-05, 2.61155424774181e-05, 
    1.93205982168854e-05, 1.37026898016994e-05, 9.29378173526483e-06, 
    6.20703624680743e-06, 3.95314951627439e-06, 2.26027472423564e-06, 
    1.161988679667e-06, 4.04823991211393e-07, 5.24920746180289e-09, 
    1.88287831379312e-12, 1.57811646243063e-12, 8.94853173563114e-13, 
    7.319912527544e-13, 6.06570564658842e-13, 4.75898734215605e-13, 
    4.81935660749036e-13, 1.28776382176929e-12, 3.60171513358676e-12, 
    7.38021434212413e-12, 9.49225345939256e-12, 2.20212806920975e-11, 
    6.72209849858581e-11, 8.83227137211686e-11, 1.10321984232649e-10, 
    1.57200383003875e-10, 9.45218991926999e-10, 1.47894434643046e-09, 
    1.26317032919171e-09, 1.49165289358711e-09, 3.15210094236235e-08, 
    1.5068378754502e-06, 1.60105994431928e-06, 1.83268445527397e-06, 
    1.76802331420152e-06, 2.1023940160217e-06, 1.23734416863738e-08, 
    1.29579285302928e-08, 1.33778520347457e-08, 1.43587586543676e-08, 
    1.50790025766725e-08, 1.37714401550552e-08, 1.16171661848293e-08, 
    1.08787563693547e-08, 8.7803774610885e-09, 4.84605295342148e-09, 
    9.11454602244042e-09, 4.13614241575916e-09, 7.39678782061544e-11, 
    1.61990626252717e-11, 9.20379328916303e-08, 1.13570016600503e-07, 
    5.31166390687251e-07, 5.52995646694255e-07, 7.75480969030341e-07,
  1.84771844984617e-07, 4.67309892598242e-07, 1.27437369676956e-06, 
    1.63352608302489e-06, 1.72313189447549e-06, 2.17929046265735e-06, 
    3.1761116976214e-06, 4.52851244367535e-06, 7.47780650552601e-06, 0, 0, 0, 
    0, 0, 0, 0, 2.78629769804893e-06, 5.03780392430006e-06, 0, 
    2.96013941791592e-06, 3.04709394965895e-06, 1.47954235821009e-06, 
    4.58137153820443e-06, 3.38123262733936e-06, 2.82771710798551e-06, 
    3.85965646922721e-06, 3.35940907478846e-06, 3.55308390799919e-06, 
    3.51920374093871e-06, 3.84032655477573e-06, 3.8839054247175e-06, 
    4.22667568539721e-06, 4.29718556107905e-06, 4.50025654004033e-06, 
    4.63253471465105e-06, 4.7313761962841e-06, 4.87934814579482e-06, 
    5.35452561748697e-06, 5.74778653875434e-06, 6.10451498961382e-06, 
    6.53277980219437e-06, 6.46646510994618e-06, 6.72159959316242e-06, 
    6.83964077835864e-06, 7.23802666723848e-06, 7.28427013457656e-06, 
    7.51192855884416e-06, 7.68804819327109e-06, 7.80400111050718e-06, 
    8.19903856058117e-06, 8.4816079294242e-06, 8.85768827304556e-06, 
    9.33929460571647e-06, 9.88434847366396e-06, 1.03149436668772e-05, 
    1.0656810421896e-05, 1.09036975337741e-05, 1.10208905699246e-05, 
    1.06963650532053e-05, 1.02179026463098e-05, 9.31162253118178e-06, 
    1.5398539337679e-05, 1.34157468906167e-05, 1.01603817859176e-05, 
    6.7974495343253e-06, 9.41014902604985e-06, 3.97459954948465e-06, 
    1.49160079011437e-06, 8.61701877895989e-07, 6.70947648307356e-07, 
    6.36510505114757e-07, 0, 3.16333743029731e-06, 4.50714900479953e-06, 
    5.58194945431134e-06, 7.13261454019253e-06, 1.0973185371007e-05, 
    1.39717226166102e-05, 1.81827515315308e-05, 2.22324965599547e-05, 
    2.61518256439057e-05, 2.97566418610838e-05, 3.32776746825536e-05, 
    3.67030162395329e-05, 3.89576172995579e-05, 4.07945085787317e-05, 
    4.21334744406686e-05, 4.25399067817573e-05, 4.139684031477e-05, 
    4.0878488548239e-05, 4.10840304255028e-05, 4.03322999109126e-05, 
    3.95581916361883e-05, 3.84400035107721e-05, 3.71155513153975e-05, 
    3.57384485270955e-05, 3.43754824014763e-05, 3.27074856062147e-05, 
    3.07973330517606e-05, 2.88428272017397e-05, 2.6549561506559e-05, 
    2.42728382133569e-05, 2.18240620758498e-05, 1.96878066857387e-05, 
    1.84408677981566e-05, 1.59438526997308e-05, 1.31040216663374e-05, 
    9.95378846097462e-06, 8.39096769807208e-06, 6.95173984289581e-06, 
    5.8886112764092e-06, 4.97546849397568e-06, 4.03479694118884e-06, 
    3.32460182242774e-06, 2.58043906208516e-06, 2.05295648209054e-06, 
    1.53221129822274e-06, 8.76787969065635e-07, 6.63275648378244e-07, 
    4.31499288381239e-07, 2.01558279537113e-07, 3.55828402004161e-07, 
    1.56823990616179e-07, 1.87794626648602e-07, 2.43746307825004e-07, 
    2.69060552514759e-07, 3.97884451687218e-07, 1.12890319520763e-07, 
    1.21436874385845e-07, 1.03014430271763e-08, 1.1639719890929e-08, 
    1.0600410209076e-08, 1.06510564708755e-08, 1.3409973015057e-08, 
    2.08508204140243e-08, 2.97375280742884e-08, 3.77342719343924e-08, 
    4.10182918291255e-08, 2.8709885353652e-08, 2.48073491336731e-08, 
    1.02896438844643e-07, 2.19525038993119e-07, 3.59834206656777e-07, 
    2.52554550307956e-07,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3.34921335714216e-09, 7.41259084466957e-09, 
    1.08626143236844e-08, 1.37496598917243e-08, 1.56111843070411e-08, 
    1.65496678218322e-08, 1.67290990929163e-08, 1.59959301348059e-08, 
    1.44059654520563e-08, 1.20703482146009e-08, 9.02064302995467e-09, 
    5.41729757514403e-09, 1.55225796267597e-09, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.68886274015136e-09, 
    7.57144096812027e-09, 1.22356672141639e-08, 1.6368837890504e-08, 
    1.99648497330377e-08, 2.30025383638465e-08, 2.5253241413785e-08, 
    2.66289941667525e-08, 2.7046041905214e-08, 2.65450039056276e-08, 
    2.50209379039731e-08, 2.28343689142069e-08, 2.12990439006454e-08, 
    1.9556993937746e-08, 1.72248784974974e-08, 1.40425397499025e-08, 
    1.00766306925013e-08, 6.68640255957172e-09, 3.30990730579823e-09, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2.21966948884756e-09, 9.3966249726325e-09, 
    1.65144388436339e-08, 2.34238691302324e-08, 3.03094373485659e-08, 
    3.75572210024623e-08, 4.55575864641448e-08, 5.39723896205946e-08, 
    6.30210760051932e-08, 7.10588013456901e-08, 7.75950681610926e-08, 
    8.2719956922955e-08, 8.69045721735424e-08, 9.00762685499005e-08, 
    9.22199450298662e-08, 9.28051300007852e-08, 9.22550116759142e-08, 
    9.06650770596901e-08, 8.82544290486902e-08, 8.49603201057507e-08, 
    8.00064691515345e-08, 7.34242642859841e-08, 6.47152762084138e-08, 
    5.42172576615155e-08, 4.34564069750756e-08, 3.32573203390668e-08, 
    2.37937845983198e-08, 1.48567335331236e-08, 6.94512817056443e-09, 
    2.38695797066465e-10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0 ;

 fprec =
  8.03798132669413e-11, 8.10150881960469e-11, 8.16341368258176e-11, 
    8.2722052376085e-11, 8.4164320609457e-11, 8.46434207585672e-11, 
    8.59677761122404e-11, 8.62806070189787e-11, 8.64973186594349e-11, 
    8.66251992163868e-11, 8.478940424093e-11, 8.4686320747227e-11, 
    9.08880003669685e-11, 9.06309148790172e-11, 9.02807171616317e-11, 
    8.98561134149865e-11, 8.18404146076789e-11, 8.11907587479925e-11, 
    7.57088860233054e-11, 7.49426997928475e-11, 7.4188780650487e-11, 
    7.34386155156715e-11, 7.10574304601552e-11, 7.03743949973172e-11, 
    6.49618777339904e-11, 6.443867163873e-11, 6.40339698482086e-11, 
    6.38011232446294e-11, 6.26523733901874e-11, 6.2728714062462e-11, 
    5.52427736605869e-11, 5.57011866958146e-11, 5.63258852504738e-11, 
    5.70906254109403e-11, 5.79726246184514e-11, 5.89392784725355e-11, 
    6.80720152983794e-11, 6.89733028685816e-11, 6.9862683904449e-11, 
    7.07343714706078e-11, 7.15580384180345e-11, 7.22928333678613e-11, 
    6.78972476156948e-11, 6.84668342369521e-11, 6.88957708468683e-11, 
    6.91511472496285e-11, 6.92409388866102e-11, 6.91788891764388e-11, 
    6.66292211039014e-11, 6.62233220372802e-11, 6.56597960461204e-11, 
    6.49596683248158e-11, 6.41565993923239e-11, 6.325578952753e-11, 
    7.26833814365169e-11, 7.18628959036842e-11, 7.10363835726583e-11, 
    7.02362133782705e-11, 6.94709989125897e-11, 6.87418289868192e-11, 
    5.9796415868313e-11, 5.91858297472003e-11, 5.87334133500398e-11, 
    5.84480746858527e-11, 5.83325003685044e-11, 5.83886806565502e-11, 
    5.27011641318232e-11, 5.31849534049138e-11, 5.38396844755598e-11, 
    5.46559371911278e-11, 5.55841789103204e-11, 5.66009398614857e-11, 
    5.0150804306743e-11, 5.14474491533171e-11, 5.27200397305069e-11, 
    5.39513099025591e-11, 5.46481784716864e-11, 5.57332257328956e-11, 
    6.98960697066841e-11, 7.0577006644755e-11, 7.37638123100718e-11, 
    7.41545587777418e-11, 7.57750967490082e-11, 7.58231164216734e-11, 
    1.035096985381e-10, 1.04190619898294e-10, 1.04115945664549e-10, 
    1.0393245158236e-10, 1.03648908612614e-10, 8.56455103641916e-11, 
    1.02771612056344e-10, 1.02500916876385e-10, 1.02070071190117e-10, 
    1.0165328336092e-10, 1.01259740054516e-10, 1.00885718935932e-10, 
    8.31940429304965e-11, 8.28090067090647e-11, 8.25027767145666e-11, 
    8.23079045049218e-11, 8.22157694201503e-11, 8.22297716622098e-11, 
    7.27966316038992e-11, 7.31156868478972e-11, 7.35665198245542e-11, 
    7.41193746089658e-11, 7.47402397902212e-11, 7.54116112630524e-11, 
    6.21328342396089e-11, 6.31395270242067e-11, 6.41398637145774e-11, 
    6.51175433842178e-11, 6.60315566651871e-11, 6.68575182471701e-11, 
    6.75835076277687e-11, 6.81650211920518e-11, 6.85883969695973e-11, 
    6.88445262711246e-11, 6.8934144230579e-11, 6.88537753855942e-11, 
    6.8603670658248e-11, 6.81799969631173e-11, 6.75983196686e-11, 
    6.68896446542481e-11, 6.60645618925067e-11, 6.5135806693188e-11, 
    6.41354337395428e-11, 6.30975254229162e-11, 6.2048970556205e-11, 
    6.10172388432163e-11, 6.00394602536041e-11, 5.91345223374824e-11, 
    6.14557846655984e-11, 6.08293271779521e-11, 6.03369851634626e-11, 
    6.00073306463975e-11, 5.98505676099334e-11, 5.98388202223692e-11, 
    7.31314660767495e-11, 7.33738480436644e-11, 7.37459404082931e-11, 
    7.42017623490394e-11, 7.47534160264954e-11, 7.24292189446495e-11,
  0, 2.66024079763018e-11, 9.63802274128126e-11, 2.47323772925662e-10, 
    5.63322371959029e-10, 1.52240639144163e-09, 3.20073583866983e-09, 
    5.28804944774369e-09, 8.44609097483169e-09, 1.15301421307861e-08, 
    1.30917220921147e-08, 1.51367085824616e-08, 1.53111807976175e-08, 
    1.39809105528015e-08, 9.46699769289928e-09, 5.97697218759231e-09, 
    2.19671420417693e-09, 9.70908434339036e-11, 2.14464856893811e-11, 
    1.63463700183267e-11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6.3201246307701e-13, 7.89062556255672e-11, 1.2492309177955e-08, 
    1.83560124271343e-07, 5.23932871118919e-07, 9.14584714848565e-07, 
    1.28338196675714e-06, 1.46247170055283e-06, 1.63328860419225e-06, 
    1.75291150526498e-06, 1.80177140099065e-06, 1.88312755544416e-06, 
    1.88116612016139e-06, 1.81620451984371e-06, 1.79281200980339e-06, 
    1.71564876213794e-06, 1.69456955127426e-06, 1.64569273003764e-06, 
    1.59569577698272e-06, 1.52543755631422e-06, 1.43257488356768e-06, 
    1.28305890854256e-06, 1.1689358915061e-06, 1.10254925204855e-06, 
    1.04577871571763e-06, 9.65453627302507e-07, 9.36486390446543e-07, 
    9.40153683174036e-07, 9.76637347427504e-07, 1.0613129796608e-06, 
    1.10650427927476e-06, 1.09508155258698e-06, 1.14069106115446e-06, 
    1.16849845734651e-06, 1.22888490362904e-06, 1.35231806292592e-06, 
    1.48193213022155e-06, 1.61583614180959e-06, 1.72441537421121e-06, 
    1.81659738655972e-06, 1.79429461965971e-06, 1.75697886080914e-06, 
    1.76355577547972e-06, 1.81399853297437e-06, 1.87477924119005e-06, 
    1.90258643880914e-06, 1.88201348474349e-06, 1.88709574316305e-06, 
    1.85373160258291e-06, 1.84924761113678e-06, 1.85001694774152e-06, 
    1.86452046067135e-06, 1.88980103812682e-06, 1.93117054967065e-06, 
    1.89768199493061e-06, 1.78208751972878e-06, 1.48558147474699e-06, 
    1.08666008357265e-06, 6.44573678219862e-07, 2.61386382631949e-07, 
    4.43939609548882e-08, 6.18184500923194e-10, 2.09623979509354e-10, 
    1.08889143773514e-10, 4.85827251787003e-11, 1.34026074822707e-11, 
    8.4535112821009e-13, 0, 4.7685867431265e-13, 0, 0, 0, 0, 0, 
    2.6392756668339e-11, 1.70434787362171e-11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 7.67553413647131e-11, 1.82192998704726e-10, 7.90521222311683e-10, 
    3.36427819961081e-09, 1.43598090690947e-08, 3.4516305806081e-08, 
    7.82694062669174e-08, 1.34056957403254e-07, 1.83243040637917e-07, 
    2.23852484720436e-07, 2.53906757552814e-07, 2.48831152890745e-07, 
    2.13094093189118e-07, 1.66493046608696e-07, 1.31563551529084e-07, 
    8.19029570971176e-08, 1.93128596039349e-08, 3.70210091659387e-09, 
    1.7227943728053e-09, 1.09447946641268e-09, 7.0834983810011e-10, 
    4.29010225212328e-10, 3.06655468536951e-10, 3.47539845657401e-10, 
    3.38742215249648e-10, 4.85466889031082e-10, 3.64620852458082e-10, 
    9.52544030093629e-11, 1.66692078401755e-10, 2.92697721148054e-10, 
    1.32583848897177e-10, 3.11770825692173e-10, 2.67248862346997e-10, 
    1.64841390956226e-10, 1.26529373501816e-10, 0, 0, 0, 0, 0, 0, 
    5.17202732353462e-12, 1.09972106780769e-08, 2.09597429320271e-07, 
    3.56695503026104e-07, 4.3577892764228e-07, 5.73497859642151e-07, 
    7.27129188469437e-07, 8.44614556881376e-07, 9.7637786270827e-07, 
    1.04120863523806e-06, 1.08600932334679e-06, 1.07644672425871e-06, 
    9.94897678189406e-07, 9.07476526790881e-07, 8.79536665324649e-07, 
    8.79527059213502e-07, 8.53849147293353e-07, 8.39125411195396e-07, 
    8.27618091797947e-07, 8.53468348478095e-07, 8.67273538346184e-07, 
    8.92987113333343e-07, 1.15667189467255e-06, 1.59077253276831e-06, 
    1.40151488324539e-06, 1.36815139352636e-06, 1.3128785234707e-06, 
    1.39615761418734e-06, 1.60293425701201e-06, 1.69398757245791e-06, 
    1.52848427355552e-06, 1.19602446418751e-06, 8.17607487297085e-07, 
    3.8935853059017e-07, 1.13684209490509e-07, 2.27244259333007e-08, 
    2.90406739640841e-09, 3.16981520150625e-09, 2.29746365179637e-09, 
    1.86192288221996e-09, 1.35620782709528e-09, 1.0773046723429e-09, 
    8.34328080137434e-10, 6.25912064515525e-10, 4.6149771273274e-10, 
    3.34997442361936e-10, 2.44156297225637e-10, 1.85724945005074e-10, 
    1.57851359983489e-10, 2.19503814477971e-10, 2.5823767006057e-10, 
    3.07876201660583e-10, 3.11910204372877e-10, 3.20835569091014e-10, 
    1.61106267318606e-10, 1.19405383744953e-10, 6.36105482758847e-11, 
    1.52901115598899e-11, 1.0288978175264e-12, 0, 0, 1.73284541915277e-10, 
    4.22626319926777e-10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3.93941894651764e-11, 3.1012088037321e-12, 0, 0, 0, 4.27822380776187e-11, 
    9.28774376213442e-09, 6.24843993383959e-08, 1.89664903333448e-07, 
    3.14731786093255e-07, 4.36676073761323e-07, 4.18111782686996e-07, 
    4.27403987178922e-07, 3.75623661864583e-07, 2.5460351936268e-07, 
    2.11052705422109e-07, 2.1722978820632e-07, 2.28136595890714e-07, 
    2.12798130083536e-07, 1.89091518016288e-07, 1.68640589942016e-07, 
    1.53775358574831e-07, 1.47279917408205e-07, 1.47032919070514e-07, 
    1.53599628589648e-07, 1.59239550930936e-07, 1.54408066317394e-07, 
    1.28160523446871e-07, 6.49222737445074e-08, 2.18935581316435e-07, 
    1.31566424975094e-07, 2.47464513455246e-07, 1.73064688402475e-07, 
    7.800927210176e-08, 3.23539287847901e-08, 1.32222136393583e-08, 
    3.44063884089341e-09, 1.49992752933593e-10, 2.54903881999459e-12, 0, 0, 
    0, 0, 1.09112523818453e-11, 1.26672099241155e-07, 5.00421803203397e-07, 
    4.4423788583743e-07, 4.85399560773121e-07, 3.7061982824748e-07, 
    4.58557320926325e-07, 4.70123192688078e-07, 6.50448653724326e-07, 
    5.10916814839047e-07, 4.24183887654289e-07, 4.10200923112099e-07, 
    4.47146630556202e-07, 5.47365900645139e-07, 6.54208422262141e-07, 
    6.52123799552194e-07, 3.790019915695e-07, 4.98754852805623e-08, 
    2.94637497079601e-09, 2.68581772266883e-09, 2.17641057949269e-09, 
    3.30019463792106e-09, 4.30590318444857e-09, 4.69200537437448e-09, 
    6.66121895375631e-09, 8.10840996932106e-09, 7.21947293014419e-09, 
    8.26357030548698e-09, 6.47378570071233e-09, 4.77423972573326e-09, 
    1.64898070419914e-09, 6.62424292980586e-10, 7.80734017312372e-11, 
    4.20091924419669e-11, 1.34501988494713e-11, 2.96123855834135e-12, 
    2.17157876527803e-13, 0, 0, 4.14412137096495e-13, 0, 0, 0, 0, 0, 0, 0, 0, 
    3.86224638974057e-12, 6.42436975918542e-11, 1.13124604911962e-10, 
    1.19931736650976e-07, 3.90856303498109e-07, 5.82272248057498e-07, 
    6.22136992766728e-07, 5.31115867467716e-07, 3.57188307034119e-07, 
    1.2885685733229e-07, 3.96758137761553e-09, 3.16059207154655e-11, 
    5.12780666828606e-10, 1.23680538360094e-09, 1.24381876631924e-10, 
    7.46813480043053e-10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 7.17207278726641e-12, 0, 6.96551228982796e-12, 
    2.55790827448145e-13, 2.91983307543704e-10, 4.50427276080941e-10, 
    6.44050266635266e-10, 4.6304255349248e-10, 2.07843832446347e-10, 
    2.11709160787522e-10, 1.25625703453728e-09, 2.66794283251647e-09, 
    3.6848439211805e-09, 7.42841149488179e-09, 6.7857804784092e-09, 
    5.37827317096988e-10,
  3.86145894312219e-07, 2.42747277800048e-08, 3.81941538135005e-10, 
    2.53050383364707e-13, 0, 2.20675956841403e-12, 5.53620782084061e-10, 
    2.70395632162309e-08, 1.36843603822729e-07, 4.05880818941365e-07, 
    6.68525627640613e-07, 7.11728966114611e-07, 8.63095813729043e-07, 
    9.88202024017468e-07, 9.5839542607537e-07, 8.87213868321006e-07, 
    8.17667833327013e-07, 7.74740061207446e-07, 7.60825083592568e-07, 
    7.56384338245764e-07, 7.44145505469672e-07, 7.31590876781675e-07, 
    6.45435603458055e-07, 7.02287569698101e-07, 7.28458987080062e-07, 
    5.95281534701724e-07, 4.56694351351882e-07, 5.76624492557851e-07, 
    4.72843616252655e-07, 4.53657173397433e-07, 4.58479632104455e-07, 
    4.31227390187974e-07, 4.05452172569701e-07, 3.46437769198304e-07, 
    2.72310846908171e-07, 1.41102188964338e-07, 5.36479484713841e-08, 
    3.43657327681072e-09, 1.88507791130794e-09, 2.35775030477505e-09, 
    2.57270730077723e-10, 0, 0, 0, 9.83643485040778e-10, 
    4.48247470188116e-08, 4.32202047231971e-07, 3.87315395089768e-07, 
    3.75512515559755e-07, 4.94698531875802e-07, 4.33758423499185e-07, 
    6.25742307281343e-07, 6.22410884033327e-07, 5.39996733433196e-07, 
    5.82186619186883e-07, 7.21670204860872e-07, 8.64408258955598e-07, 
    9.49099691368838e-07, 9.50800629086091e-07, 1.02408463022734e-06, 
    8.38597389558559e-07, 4.84482484499837e-07, 1.59688508981674e-08, 
    1.86829533419848e-10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.51608796015419e-09, 1.69342287565561e-11, 5.83847772989069e-11, 
    4.76901382338608e-11, 2.72007639698151e-11, 6.27997712943015e-11, 
    1.3835405628764e-11, 3.74118547845916e-14, 1.61874299732722e-11, 
    9.24914698512908e-12, 9.04385708594249e-11, 1.43910975284674e-11, 
    4.19936131295449e-10, 1.27287692537181e-06, 5.92780768893242e-06, 
    9.02075355186016e-06, 1.1813257688543e-05, 1.37718961624436e-05, 
    1.41087696846355e-05, 1.23056203472694e-05, 5.60517950060909e-06, 
    1.52165091448823e-08, 2.12977471885047e-08, 2.66288176955852e-07, 
    1.22298154087743e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5.57418882593053e-11, 0, 0, 0, 0, 0, 0, 3.85103768567546e-11, 
    2.25326535116904e-11, 6.58615858568958e-11, 6.47364075883818e-10, 
    3.20062197613512e-09, 2.06666036440499e-08, 8.21605024498008e-08, 
    2.77138432617251e-07, 6.96246973378664e-07, 1.16253425728815e-06, 
    1.55171489403869e-06, 1.94106066252501e-06, 2.2959715264608e-06, 
    2.28904555886704e-06, 2.23558350882906e-06, 1.78910050489561e-06, 
    1.09599618817304e-06,
  3.74198638025562e-06, 2.59243724066425e-06, 2.33899366765797e-08, 
    1.10389036421216e-11, 4.314442629767e-10, 4.90977594059522e-09, 
    6.27882599292957e-09, 3.87679411318006e-08, 8.19005995904265e-08, 
    2.05240833704299e-07, 2.88495084981449e-07, 4.98543963943989e-07, 
    4.90160974839975e-07, 4.10304645783038e-07, 3.20505867963572e-07, 
    3.10849000599997e-07, 4.37105421060422e-07, 6.10430934066238e-07, 
    7.30809786233614e-07, 7.51051078803722e-07, 9.02210620712917e-07, 
    1.04467145767849e-06, 1.07752792775915e-06, 1.07012746353523e-06, 
    9.40300793407081e-07, 7.41074678383203e-07, 6.23858996769417e-07, 
    4.11371533499936e-07, 2.41399634667766e-07, 1.75819179187294e-07, 
    1.68139770269741e-07, 1.939605159451e-07, 2.43006682126297e-07, 
    3.32256824434336e-07, 4.05533300880297e-07, 5.32871725726465e-07, 
    4.22388841744657e-07, 2.71252495271868e-07, 1.52116254260884e-07, 
    6.80447525210572e-08, 7.11349454783319e-09, 1.34444396311876e-10, 
    9.03248433018167e-10, 2.32238184030166e-09, 3.21723589876736e-10, 
    3.52176637932501e-08, 1.51276243846503e-07, 4.92497974483755e-07, 
    3.34991868184046e-07, 3.45955279512889e-07, 4.25548572450915e-07, 
    4.46059215431175e-07, 5.75621225188669e-07, 7.72662737740167e-07, 
    1.01874431769463e-06, 1.13456335000004e-06, 1.12696179191636e-06, 
    1.13769811303933e-06, 1.25112717411204e-06, 1.18318578594574e-06, 
    1.28304702922242e-06, 1.21877544621488e-06, 6.4107143090692e-07, 
    2.02847546772733e-08, 1.96412595342633e-12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6.15966889728531e-12, 1.66988303367947e-09, 2.47149735356354e-08, 
    9.53500665992034e-08, 6.48909179455262e-08, 1.91178282684516e-07, 
    7.43179367041107e-07, 9.91716156934606e-07, 7.28016053831054e-07, 
    1.64893653177809e-07, 3.82522424331688e-09, 4.21519542093067e-09, 
    8.44127946411861e-10, 5.5256045143038e-09, 4.10348103235144e-09, 
    5.91851295617275e-09, 1.32268193781067e-08, 2.11041525745793e-08, 
    2.87594141114035e-08, 8.15037974250153e-08, 5.10252070020926e-07, 
    4.7832849120514e-06, 7.9052282408641e-06, 1.01818253099902e-05, 
    1.20372359522092e-05, 1.4621946769176e-05, 1.27819848828793e-05, 
    1.5555894000118e-07, 1.18337960634483e-11, 5.13156477381847e-11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 9.07274068123529e-11, 4.09717347825893e-09, 
    6.98282984934388e-08, 5.13225424954672e-08, 2.01079434164555e-09, 
    2.46327998300362e-09, 1.4593908415803e-08, 2.0788471423262e-09, 
    4.87225634180975e-09, 3.96477351647708e-08, 3.73036406769574e-12, 
    1.25193562426349e-11, 3.23213173573897e-08, 2.00349302601069e-07, 
    2.26290849481416e-07, 1.77947915429427e-06, 2.85488022814429e-06, 
    4.94961051653858e-06, 6.20297701490809e-06, 7.74932528139623e-06, 
    9.28312975497673e-06, 1.05045807996374e-05, 1.07410645857205e-05, 
    9.71464927124912e-06, 9.29378029588717e-06, 9.48409872436659e-06, 
    8.14030906159833e-06, 6.08977565898001e-06, 4.96726206528542e-06,
  2.5408451603371e-06, 1.88288774508109e-06, 2.33429339990212e-10, 
    6.17606383382238e-10, 9.55827246142353e-08, 2.20215158220269e-07, 
    4.08661412774173e-07, 1.35114782511887e-06, 2.04658460258819e-06, 
    1.84072577774804e-06, 1.34449295545976e-06, 9.93316022184905e-07, 
    6.92904389315931e-07, 7.60955577477862e-07, 6.75431686728777e-07, 
    5.3148732549114e-07, 5.34633017134423e-07, 8.37243549306869e-07, 
    1.15265328139551e-06, 1.54403549048034e-06, 1.95767764502787e-06, 
    2.20395257934116e-06, 2.36206111453036e-06, 2.43301646561843e-06, 
    2.30801452564482e-06, 2.07009908053957e-06, 1.64368350089277e-06, 
    1.3000804383768e-06, 1.11335767300477e-06, 1.05287262524172e-06, 
    9.06272830869457e-07, 8.04568902518284e-07, 3.88542299988057e-07, 
    1.40189678148115e-07, 1.43298313941273e-07, 9.52723650127411e-08, 
    7.38253428069428e-08, 4.07175190118113e-08, 5.12745845408582e-08, 
    3.85146898290159e-08, 9.90490190429327e-09, 3.01484926571563e-09, 
    1.17298384451481e-09, 1.56293191711676e-08, 2.58646743745536e-08, 
    4.91292785136612e-08, 4.88352116443532e-08, 1.50060069778252e-07, 
    5.12999978399965e-07, 4.01166093252789e-07, 4.20327998716032e-07, 
    5.13620634254314e-07, 6.98359070138159e-07, 8.07075284939556e-07, 
    9.35328441493778e-07, 1.02176340117204e-06, 9.19370230549082e-07, 
    8.63360972145817e-07, 8.30150434046837e-07, 7.14585086231648e-07, 
    6.59860063188872e-07, 4.55190121047024e-07, 2.06977869174597e-07, 
    3.54168470841036e-08, 5.9830497823655e-12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.65299442182828e-11, 0, 4.73309078496417e-06, 5.05715412595497e-06, 
    7.29097291427596e-06, 1.1259529020184e-05, 1.17796432034706e-05, 
    9.02823075128367e-06, 6.01090732401232e-06, 3.62923349068973e-06, 
    2.39637803504391e-06, 1.96087032447534e-06, 2.35673284325964e-06, 
    2.19154745090815e-06, 3.46705973743149e-06, 4.2271726413432e-06, 
    4.19561689233693e-06, 6.15772917431773e-06, 7.83339024064326e-06, 
    7.93463077499575e-06, 1.72074265545034e-05, 2.3354582011329e-05, 
    3.2615082326294e-05, 4.24061873795981e-05, 5.16487717637419e-05, 
    5.56136664806418e-05, 5.12594365561002e-05, 4.32651297529107e-05, 
    3.08697648656904e-05, 7.23226863010705e-06, 2.53771917069182e-12, 0, 0, 
    0, 0, 0, 0, 0, 5.06833854429573e-10, 1.12392229553152e-07, 
    6.51051713893382e-07, 1.1218329870489e-06, 1.15805198784299e-06, 
    1.04148932340519e-06, 1.36487674254862e-06, 1.34461560318668e-06, 
    9.85191529018061e-07, 5.59044048610489e-07, 4.52479519250648e-07, 
    7.5719633823066e-08, 0, 0, 1.44055452252413e-09, 4.81261378243961e-08, 
    1.6279128096796e-07, 3.00872240249769e-06, 6.31956697793956e-06, 
    1.22041548759421e-05, 1.42952985591855e-05, 1.67763298137348e-05, 
    1.58757995064764e-05, 1.47703214272674e-05, 1.31933029056461e-05, 
    1.13204501920351e-05, 8.59826093342867e-06, 7.12956326188321e-06, 
    6.35156948205403e-06, 5.3957266378016e-06, 3.56396432714242e-06,
  0, 2.01785480771983e-10, 6.36632207266154e-08, 1.2198560817146e-07, 
    1.48503286207275e-07, 3.24453282913562e-07, 8.37729280850818e-07, 
    1.0620246467538e-06, 9.52702149412422e-07, 9.76871036945163e-07, 
    9.40099282354693e-07, 7.54113736217175e-07, 5.3714281472686e-07, 
    6.30384529743124e-07, 4.88899951573786e-07, 5.34387626514022e-07, 
    7.11263515083444e-07, 1.1363145159675e-06, 1.51205319062922e-06, 
    2.17173390882243e-06, 2.68931619436589e-06, 3.21465095947171e-06, 
    3.84130908004575e-06, 4.8560547051222e-06, 5.38471728098322e-06, 
    4.66425050134733e-06, 3.06347043230615e-06, 2.53056941365516e-06, 
    1.66497509915167e-06, 9.8983725493118e-07, 2.27766773589975e-07, 
    2.14155128777098e-08, 5.13022154170221e-08, 8.18236972647802e-08, 
    9.33019339154269e-08, 8.26458057431512e-08, 1.09493239052554e-07, 
    5.98376059187789e-08, 5.04015265489138e-08, 3.87336502757861e-08, 
    1.9249150842814e-09, 8.71826237168342e-09, 6.86753045572307e-09, 
    1.15218602741228e-09, 7.84311939564248e-09, 1.80390816751223e-08, 
    1.84381338379122e-08, 3.26281318958771e-08, 1.13590739191394e-07, 
    2.34336191423505e-07, 2.33570337223469e-07, 2.76644299240109e-07, 
    3.47242939912728e-07, 4.50637746655256e-07, 5.18607426333196e-07, 
    5.15116566391405e-07, 4.83537772135283e-07, 3.74272675859897e-07, 
    3.6603809682468e-07, 3.7949002647493e-07, 3.856524193761e-07, 
    3.0319186471436e-07, 1.92753043038855e-07, 2.58706962728804e-08, 
    1.65822515249822e-09, 0, 0, 0, 0, 0, 0, 1.64114568175022e-09, 
    3.40140064935623e-09, 1.10137226567938e-10, 1.96802118587826e-09, 
    1.0106587560832e-10, 0, 1.23710320531403e-07, 2.53104095194656e-06, 
    3.72844854712229e-06, 7.93640301506728e-06, 9.87042293114508e-06, 
    7.45157552623871e-06, 6.91405743106284e-06, 9.44307149756502e-06, 
    1.24442152377809e-05, 1.67030933610242e-05, 1.9314749051305e-05, 
    2.02987929783604e-05, 2.29252856762169e-05, 1.81775165883059e-05, 
    1.67004597638479e-05, 1.901914248835e-05, 1.98532227284241e-05, 
    2.39855178430371e-05, 3.24268372671235e-05, 6.20249269574776e-05, 
    9.49685386207851e-05, 0.000133228881237494, 0.000163888702071398, 
    0.000178743693444565, 0.000186029949946519, 0.000163418807432557, 
    0.000119058889048658, 5.35890893500709e-05, 1.43179850085986e-08, 
    7.24536546041748e-12, 0, 0, 0, 0, 0, 0, 1.19143695761098e-10, 
    9.30043808055186e-08, 2.02025654087943e-06, 5.12472014655821e-06, 
    6.60293113114939e-06, 5.85551192782672e-06, 3.37582614706259e-06, 
    1.82437162811196e-06, 7.75203129574755e-08, 8.35328015422305e-08, 
    1.11174939767053e-06, 1.82540303955186e-06, 4.60857549840946e-06, 
    8.41697256835053e-06, 3.26133617851005e-06, 2.73032030383176e-08, 
    9.83168754709393e-07, 1.51334138124763e-06, 9.49589040215164e-06, 
    2.15976484133512e-05, 4.29312818211218e-05, 6.19635202601453e-05, 
    6.58914314264796e-05, 5.8055298398655e-05, 4.69474220871565e-05, 
    3.17011335585553e-05, 1.92765221685197e-05, 8.35422637833873e-06, 
    2.79089540097953e-07, 3.35641119399015e-08, 7.39959816056592e-12,
  1.76376454759093e-14, 0, 2.47272480104122e-10, 2.19978447336498e-10, 
    3.15885252301346e-10, 8.57143782419023e-08, 2.55590762417411e-07, 
    4.6117024059383e-07, 7.73190764632384e-07, 1.32223415455241e-06, 
    1.89246314675627e-06, 2.25924806031013e-06, 2.25378750986885e-06, 
    1.79381682250588e-06, 1.32482071381981e-06, 1.22364837117016e-06, 
    1.57289067321165e-06, 1.46231002444613e-06, 2.07392571067803e-06, 
    2.6690752647358e-06, 3.97779926399557e-06, 5.53103674162784e-06, 
    7.82612750410114e-06, 1.13960276920228e-05, 1.62862432335218e-05, 
    1.906422038347e-05, 1.52187609989222e-05, 7.16468747622816e-06, 
    3.09928379682919e-06, 3.43245699187602e-06, 3.5235616403437e-06, 
    1.69380569857461e-06, 4.01695618591516e-09, 3.15180316871041e-08, 
    5.22689256660537e-08, 1.9217001730716e-08, 3.77979054752081e-08, 
    3.84938241636229e-08, 3.15807727115385e-08, 1.81941669564784e-09, 
    1.0318150628011e-10, 2.95439262683577e-10, 2.58248169512708e-10, 
    4.43269166094649e-11, 4.25777648677714e-10, 1.2687305633036e-08, 
    1.26204898842463e-08, 1.47899389404185e-08, 1.56962477274312e-08, 
    1.14057735258085e-07, 2.44012807882749e-07, 1.65420602248164e-07, 
    1.58239307870281e-07, 2.31752996732212e-07, 2.6309955503638e-07, 
    2.61059781857084e-07, 3.0538136829761e-07, 2.43165279639112e-07, 
    2.43998777373237e-07, 2.29681571033401e-07, 2.78114177870981e-07, 
    2.88922860654532e-07, 2.97192360177316e-07, 7.07276275449547e-07, 
    4.22396922356923e-07, 5.49026268973375e-07, 7.05528332556746e-08, 
    2.08870808779342e-11, 0, 0, 2.31354403517006e-08, 9.67897653165722e-08, 
    7.63942263888009e-08, 9.48386739628384e-09, 2.52508772725389e-10, 
    4.42776776462799e-11, 0, 2.43184588394652e-10, 1.55217174498909e-07, 
    2.55614736769885e-06, 4.25055907911717e-06, 4.43042515479452e-06, 
    5.52131513699243e-06, 5.09838412950209e-06, 8.44126381649451e-06, 
    2.18495438757737e-05, 3.65344922195544e-05, 4.15516747742956e-05, 
    4.19087451271346e-05, 3.54467355752022e-05, 2.01068666987206e-05, 
    6.99601794698484e-06, 7.7330705792023e-06, 7.38285543444761e-06, 
    5.46109268392479e-06, 4.32694976641668e-06, 8.32566177415133e-06, 
    6.84812224733632e-05, 0.000103123004101213, 0.000131067964330168, 
    0.000189979523078585, 0.000249169011871363, 0.000277203641759034, 
    0.00024912522963449, 0.000208666488134986, 0.000125965101356228, 
    1.12135377065907e-05, 3.91859217724155e-10, 0, 0, 0, 0, 0, 
    3.91030673682837e-15, 6.27411868079774e-07, 4.57000522946548e-06, 
    5.15863024276503e-06, 4.85816726758775e-06, 2.63062140540646e-06, 
    1.42971025059449e-06, 8.49840054276965e-08, 9.47436336457247e-10, 
    5.2740539712082e-07, 6.91727179682089e-06, 1.95448733364573e-05, 
    3.91158933742065e-05, 5.55395244556252e-05, 6.15175965122744e-05, 
    6.19319308071323e-05, 5.30664401452351e-05, 3.76720949989436e-05, 
    2.3575451101745e-05, 9.75975675663425e-06, 1.66564023207846e-05, 
    4.10019299521148e-05, 8.12546499163751e-05, 0.000108088000124265, 
    0.000110283807778402, 8.15711473889921e-05, 4.3989900220416e-05, 
    7.26370812458344e-06, 3.10536224461646e-09, 2.37176273969907e-11, 0,
  0, 0, 0, 0, 0, 0, 3.15217072695814e-09, 3.03648419891308e-09, 
    4.62222552430397e-09, 2.52988813449196e-07, 1.09780816239383e-06, 
    2.44278067743237e-06, 4.60788404410928e-06, 7.2648626917751e-06, 
    6.81645620811939e-06, 5.09797497411721e-06, 3.02928777275783e-06, 
    1.33134658759944e-06, 6.44086620360769e-07, 1.09651667296855e-06, 
    2.6157490772481e-06, 5.35045962662102e-06, 9.4332532187584e-06, 
    1.3401762141645e-05, 1.98881628719886e-05, 2.75003827322782e-05, 
    2.84822417747579e-05, 2.90831256931521e-05, 3.10312828246227e-05, 
    2.48081957387125e-05, 1.7135675697346e-05, 1.14518480570428e-05, 
    2.8576463711234e-07, 2.98642561644688e-11, 1.73808982872206e-09, 
    9.8896766103859e-09, 3.7856658866142e-08, 2.76051282010391e-10, 
    1.14777275764676e-09, 2.37445625687217e-11, 0, 1.06584778307565e-12, 
    5.31800402512676e-14, 0, 7.76759543601636e-12, 2.50953806206495e-10, 
    4.56539940280224e-11, 2.17413314550572e-10, 2.37447955533735e-10, 
    2.99127158477532e-09, 1.14291306241403e-08, 7.16677832224392e-09, 
    2.95889693814696e-08, 5.42055160938891e-08, 1.54344932684586e-07, 
    8.60963367645845e-08, 3.6635938629164e-08, 3.29139457050336e-08, 
    2.92738423969922e-08, 7.84897355822947e-08, 2.36251367899371e-07, 
    2.69334018878857e-07, 7.67402726193731e-07, 1.61196345651234e-06, 
    2.81990470230118e-06, 4.47346231901063e-06, 1.44101025396316e-06, 
    2.33914304996735e-09, 1.84347119148995e-09, 7.59124567763991e-08, 
    9.76030277154139e-08, 1.15184066396667e-07, 2.72284253637574e-08, 
    2.85995253552909e-10, 2.87221136563499e-09, 0, 0, 0, 
    4.03834708275609e-10, 1.15524385645233e-07, 7.74519352362545e-07, 
    7.46558457566614e-07, 2.59298020452055e-06, 2.06175124985237e-06, 
    3.99376639720294e-06, 3.88448030783549e-06, 1.00235941603535e-05, 
    1.86757863474329e-05, 2.16723153679425e-05, 2.10144940798172e-05, 
    6.57082615274446e-06, 9.12089080778825e-07, 3.88859904525819e-07, 
    1.11908841011936e-07, 2.40786940298684e-09, 6.11657040062773e-12, 
    1.33656349936581e-08, 4.38539467896794e-05, 7.37289403275112e-05, 
    5.97181662813851e-05, 5.80341675589929e-05, 6.67105613780013e-05, 
    0.000103210222472748, 0.00018025275011566, 0.000255008370911955, 
    0.000275541533520231, 0.00021748129149135, 0.000127560683263669, 
    2.90318138017244e-07, 5.25673889254821e-12, 0, 0, 0, 0, 
    5.39346156705874e-09, 2.99254697554859e-07, 2.842206165857e-07, 
    6.32357730970009e-08, 3.01155809102827e-08, 1.15759926044568e-08, 
    2.50393228734289e-10, 3.14083518612147e-08, 1.43702828737573e-05, 
    3.04701584885777e-05, 5.60779111964367e-05, 5.39664708741576e-05, 
    6.4425031892759e-05, 7.21300246055221e-05, 6.83393325115788e-05, 
    5.86798310625284e-05, 4.28491363099215e-05, 2.02554931065491e-05, 
    8.63345208853238e-06, 5.39177822821421e-06, 1.58677972775867e-05, 
    4.92534285232487e-05, 8.98462587570028e-05, 0.000137724457467389, 
    0.000140828199401418, 8.23242880242754e-05, 1.49991192622013e-05, 
    5.07440767349428e-07, 0, 0,
  0, 0, 0, 0, 5.70047577806184e-12, 8.6584704055949e-07, 3.7282139274007e-07, 
    4.27950068286704e-06, 8.32703282868672e-06, 1.01903474585327e-05, 
    8.49638182239653e-06, 8.20113682490123e-06, 1.45798635468624e-05, 
    2.08482225697273e-05, 1.848915609614e-05, 1.46744287450249e-05, 
    1.26217283451541e-05, 1.18537700360418e-05, 6.48221109157449e-06, 
    1.82134782407082e-06, 1.36320250400962e-06, 2.12636571691351e-06, 
    3.94004473327122e-06, 9.81092145743704e-06, 1.73811190123986e-05, 
    3.48458542522009e-05, 6.48734673785835e-05, 0.000101899080380379, 
    0.000106534172725722, 7.54377061252292e-05, 4.60290914179081e-05, 
    3.62850511764199e-05, 1.53602599314959e-05, 2.36748670498079e-09, 
    3.92106036074854e-12, 3.27759453670236e-10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2.90471415882699e-10, 3.31759028871021e-10, 
    9.63444420835367e-10, 6.10933746567363e-10, 1.37144887328986e-08, 
    8.65446312891219e-08, 1.67008892948445e-06, 3.01720691134017e-06, 
    3.50437995099724e-06, 2.87899035553549e-06, 4.27151267281076e-06, 
    9.17862897942758e-06, 1.29644090022971e-05, 1.08365485438451e-05, 
    6.6591670450398e-06, 2.40773739757943e-08, 5.7624923772445e-08, 
    8.67439335329665e-09, 1.56864520118973e-08, 2.58852866887328e-09, 
    4.2437742940917e-10, 0, 0, 0, 0, 0, 2.31617213959868e-09, 
    3.22143072143571e-07, 1.1498704268909e-07, 2.67647332819956e-07, 
    5.54843777728788e-07, 1.96391108866937e-06, 3.44811069660027e-06, 
    2.01906989679103e-06, 3.05889558687757e-06, 1.18912975685693e-05, 
    1.14086760427307e-05, 1.1302116085478e-05, 3.738288833704e-06, 
    7.57210055261814e-07, 4.54099786369628e-08, 3.65030668351793e-10, 0, 
    1.01229298626742e-05, 0.000127102566800397, 0.000150212972628077, 
    0.000131580800224794, 7.80300241244346e-05, 3.91554227080727e-06, 0, 0, 
    0, 5.02481595495971e-05, 0.000138798543610765, 0.000192702600442522, 
    0.000184559472682925, 0.000157235886274269, 4.77723886187648e-07, 
    3.10185002927313e-09, 0, 0, 0, 2.58306026207486e-10, 
    1.63499235764233e-09, 6.56180811185718e-10, 8.77385272465819e-11, 
    3.32818017377934e-11, 6.94455706881775e-10, 3.94170708368273e-10, 
    7.74523788406961e-06, 3.92397536009587e-05, 4.95919256925488e-05, 
    1.86641810381323e-05, 7.79935812259008e-06, 1.1052999073307e-05, 
    3.03823037334125e-05, 3.10727722753922e-05, 2.14739890218938e-05, 
    1.00267890683344e-05, 3.92007079242374e-06, 3.06356916074307e-06, 
    5.13637971211935e-06, 7.23608870327646e-06, 2.59584687653522e-05, 
    4.34487126076321e-05, 5.42648145133273e-05, 5.00641471636431e-05, 
    3.04440322143981e-05, 2.14565154508298e-05, 1.87579047953996e-07, 
    9.94173979103836e-11, 0,
  0, 2.44690601807315e-07, 7.90782956278899e-06, 2.35560752901937e-06, 
    9.45477513981201e-09, 5.37575803804223e-10, 4.36732713914751e-10, 
    1.00603147638014e-07, 2.18853726556301e-06, 4.79281461927873e-06, 
    1.16429165196965e-05, 2.69661327694071e-05, 1.84224704176254e-05, 
    1.54638666423565e-05, 1.79717202093476e-05, 1.50759106989999e-05, 
    2.16085539548943e-05, 3.34476238644029e-05, 3.53334535427621e-05, 
    2.63204820321869e-05, 2.23661435948423e-05, 1.11028914465276e-05, 
    6.85970898605857e-07, 1.3584206444618e-07, 3.05477653557606e-06, 
    1.3505301493024e-05, 3.31954213096881e-05, 5.32282538683964e-05, 
    6.9804216063165e-05, 9.77872127513258e-05, 0.000130175698683823, 
    0.000126097973609751, 0.000107065962972792, 1.61048115308411e-05, 
    4.42935176285059e-09, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7.1325570895872e-11, 1.57432537040729e-10, 7.6085102430871e-08, 
    1.9584946098998e-06, 4.24367988254581e-06, 4.98437429691564e-06, 
    2.67097485938452e-06, 1.58016187763631e-06, 1.79202080646859e-06, 
    8.75453227205225e-06, 2.2622522889222e-05, 2.78371257934694e-05, 
    2.7126488919564e-05, 2.12659069122316e-05, 1.69090564171339e-05, 
    1.74679147406211e-05, 2.39725491480026e-05, 3.75314893380416e-05, 
    4.88429477535832e-05, 5.22184887495293e-05, 5.38013048092657e-05, 
    5.79065084790352e-05, 6.36260323751463e-05, 4.74521559475367e-05, 
    2.67357856790021e-06, 1.8026504656516e-06, 1.03664473968562e-06, 
    3.5393563919957e-07, 1.51966934358463e-07, 7.05786998942495e-08, 
    6.99491408608747e-08, 3.11570643623317e-07, 6.92806310124263e-07, 
    1.78101340489424e-06, 2.86110473886863e-06, 2.3371622491679e-06, 
    4.62259243297915e-06, 5.44005586509862e-06, 1.72695024115355e-06, 
    1.68452081558513e-06, 3.54211733184505e-05, 0.000178436482560605, 
    0.000236111184019254, 0.000184579059599743, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.000114108908189907, 0.000132399631251293, 0.000113698919807751, 
    7.32102528859778e-06, 6.39830319514008e-08, 8.03264434823229e-10, 0, 0, 
    2.31925723875996e-11, 0, 0, 0, 9.02024873552121e-11, 
    2.55237459712478e-07, 1.06917701988579e-05, 2.89309008316102e-05, 
    1.52869236591204e-05, 4.1618693539301e-06, 1.56955045159889e-06, 
    7.9880655101217e-06, 3.40103231525733e-05, 3.8441476969592e-05, 
    1.60862486395588e-05, 4.20547306275891e-06, 2.0120083838911e-06, 
    4.43097303948744e-06, 1.12200425846925e-05, 1.27274294978106e-05, 
    3.17922654711581e-05, 3.04456427913604e-05, 1.30878498875611e-05, 
    8.45899648152049e-06, 4.77679892143541e-06, 5.18167962096348e-06, 
    3.73762854724797e-06, 2.20599111615483e-07, 6.08645778773315e-10,
  1.13732790543258e-05, 9.91127034589773e-06, 9.71502085948754e-06, 
    3.60412663774183e-06, 1.01602745467899e-05, 4.43965818724295e-06, 
    7.99998681836682e-07, 8.88729166530008e-06, 1.35011193313804e-05, 
    1.29853039045992e-05, 1.97265685656815e-05, 1.95172543874507e-05, 
    1.37628095096658e-05, 1.36794633868959e-05, 7.74553302477647e-06, 
    2.47374900651903e-06, 5.21829419735148e-06, 7.2983436424434e-06, 
    1.91090889313594e-05, 4.61377861876032e-05, 2.8620778542105e-05, 
    3.13894240603132e-05, 2.01019302015926e-05, 5.70149764933989e-06, 
    9.27598313372707e-09, 2.06107227993367e-08, 7.46290444417962e-08, 
    1.76953736168416e-06, 1.28454433568371e-06, 4.57623345581108e-06, 
    2.01790566798314e-05, 6.51592007662475e-05, 0.000157187913597677, 
    0.000172733730339512, 9.8326054036108e-05, 2.85662897523097e-08, 
    3.50763785763091e-11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.71166428823897e-12, 
    7.98545523996314e-10, 5.64189996363781e-14, 0, 0, 0, 0, 0, 0, 
    7.12464791411109e-11, 7.05286494106522e-11, 1.27212492388532e-07, 
    3.16948042658419e-06, 1.65504905008653e-06, 1.20219835278401e-07, 
    1.41808492981901e-06, 8.02862927723536e-06, 1.4094189089556e-05, 
    4.29883523986989e-05, 6.21051938175018e-05, 5.79059858834026e-05, 
    4.52190470131364e-05, 3.88239054149036e-05, 2.45884671312229e-05, 
    1.54693978100439e-05, 1.53131236908787e-05, 2.15477744699541e-05, 
    3.25986022716847e-05, 4.83523204005209e-05, 5.9519918421734e-05, 
    5.71750328993159e-05, 7.83654885921909e-05, 0.000130607753163649, 
    0.00015714227545568, 0.000163425432491092, 8.79784643962726e-05, 
    1.02917292724137e-05, 2.80854283788843e-06, 2.79534129782383e-06, 
    2.11559511763223e-06, 7.10159655829171e-06, 1.31360537758312e-05, 
    1.31460670819223e-05, 1.04836844994951e-05, 9.01378072846832e-06, 
    1.19689634078724e-05, 7.31413487180228e-06, 7.18073449230695e-05, 
    0.000238969976977267, 0.000296156684066131, 0.000116413146146392, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3.05036586184294e-05, 4.5073701609443e-05, 
    3.01474099061873e-05, 2.08279461820092e-06, 2.12418495124551e-06, 
    2.05858440697827e-06, 3.79513638379332e-06, 5.55472895567891e-06, 
    7.9301219599222e-07, 1.55859465690301e-06, 1.16787756937699e-07, 
    2.19430686862651e-10, 1.93532337114916e-09, 2.77738120956313e-07, 
    5.4710738671858e-06, 2.67360515914377e-06, 1.50882792670299e-06, 
    2.38585289753678e-06, 3.88111155221897e-05, 5.5364025019857e-05, 
    3.52031696062135e-05, 1.45367290106259e-05, 2.61746556338599e-06, 
    4.89107018626315e-06, 1.56723118965513e-05, 5.02423454449554e-06, 
    7.10101970348467e-06, 2.10801612841075e-05, 4.21800006105464e-05, 
    1.83974764621527e-05, 3.14644832488858e-06, 1.04463149256778e-06, 
    3.1240996848876e-06, 2.20842722595916e-06, 3.48146676359898e-06, 
    2.1794054494789e-06,
  1.04277186072811e-05, 6.09471790467508e-06, 7.8908262088188e-06, 
    7.67502806356401e-06, 7.1477125829977e-06, 1.10002570511146e-05, 
    8.15562370617294e-06, 2.23268210896937e-05, 1.97327903199552e-05, 
    2.44561294208642e-05, 2.5774805894166e-05, 1.29438987686425e-05, 
    3.51912684204972e-05, 3.702515818452e-05, 1.68738129931804e-05, 
    3.21914842202482e-05, 2.95039323537438e-05, 2.73146420550759e-05, 
    1.79870465961752e-05, 2.72364191231766e-05, 1.98412216003526e-05, 
    1.42884918528261e-05, 1.0880737970852e-05, 1.39267931748767e-05, 
    2.32450789170635e-07, 1.14663101157973e-07, 9.53964120251952e-08, 
    1.43846799808744e-08, 1.07504360921258e-08, 3.41161480251189e-09, 
    1.52752329519306e-09, 5.47971710349368e-08, 1.60231168488134e-05, 
    8.93908118308898e-05, 0.000182870601780817, 0.000115333603467054, 
    3.12477763257255e-07, 1.11029590231901e-07, 3.04226786624661e-09, 0, 0, 
    0, 0, 0, 6.28402600358223e-12, 4.42392916653042e-08, 
    2.32710938880108e-06, 3.66100171100183e-06, 3.10207681733843e-06, 
    5.19430095937286e-06, 1.25822597438394e-05, 1.0385884233925e-05, 
    1.14174908109563e-05, 9.86482839800915e-06, 1.08080019040246e-05, 
    1.06165256983919e-05, 1.15853582941702e-05, 5.72404665679472e-06, 
    1.10514264938687e-05, 1.41794517683578e-05, 1.19184807706432e-05, 
    1.49613714150006e-05, 3.42586610462761e-05, 3.2131760643937e-05, 
    1.91087280945197e-05, 2.28716884079827e-05, 4.25113403939767e-05, 
    2.10672119049732e-05, 1.74237211586799e-05, 1.7075693311858e-05, 
    1.73478464670433e-05, 2.1317494027008e-05, 3.75393761256753e-05, 
    4.50838156756665e-05, 2.09498181316524e-05, 1.62240488834666e-05, 
    1.15277840571113e-05, 2.3396110127422e-05, 0, 0, 0.000199273073017639, 
    0.000199492694804503, 0.00014187446280185, 1.54020850637163e-05, 
    4.80381979229212e-06, 1.18576617103822e-05, 7.29182811295478e-06, 
    2.11881762546907e-05, 6.03449903634108e-06, 1.18936829693098e-05, 
    7.58969299464601e-06, 9.27233805092727e-06, 3.45016658556371e-05, 
    0.000241869986645921, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.89093924070067e-07, 2.85478398960337e-08, 0, 0, 0, 0, 
    5.16207157555824e-06, 4.2516651312521e-07, 2.36655565045712e-06, 
    1.7741870716132e-06, 6.97186348071551e-06, 1.76582879761075e-05, 
    2.13743737373704e-05, 2.41823961341392e-05, 1.46475173984885e-05, 
    7.92836624700181e-06, 3.31076400134341e-06, 1.09512922701126e-06, 
    7.74974208108342e-08, 1.3217032401004e-06, 2.52667844802577e-05, 
    5.71210373265352e-05, 3.74015515781814e-05, 2.68271117124386e-05, 
    7.70806083869362e-06, 2.16787609314403e-06, 1.00849531436719e-06, 
    2.09557001054378e-05, 1.78965856060558e-05, 9.02508993467196e-06, 
    3.13170210632146e-05, 5.38741770677441e-05, 2.53018606358579e-05, 
    4.57398894546047e-06, 1.16222436631725e-06, 1.63432256235592e-06, 
    2.62191664418638e-07, 9.95968087544162e-06, 1.43067546327519e-05,
  3.49742280640581e-06, 8.49404892478714e-06, 4.91074028092756e-06, 
    8.08163311608442e-06, 8.30112849899816e-06, 1.29522515569455e-05, 
    1.6913943641686e-05, 1.45260573313872e-05, 1.69303680190835e-05, 
    2.19752272114435e-05, 2.0771153114183e-05, 3.68178465053717e-05, 
    3.27102021871478e-05, 4.50188074703225e-05, 5.18097169666768e-05, 
    3.76563933764471e-05, 4.12834197427034e-05, 3.57830004207352e-05, 
    4.91397408625614e-05, 3.0693451701203e-05, 3.48308921797316e-05, 
    2.35978623302159e-05, 3.02741448949933e-05, 3.32003974904352e-05, 
    3.2451453345587e-05, 3.8370720369069e-05, 1.00375429240636e-05, 
    1.02809964083668e-05, 8.34089001780985e-08, 6.46228204842609e-07, 
    1.12143060569264e-06, 2.2454137916234e-07, 3.86590421180602e-06, 
    1.26711482479577e-05, 9.99539377041327e-05, 0.000176562159565878, 
    5.83670521736693e-06, 7.3234278585262e-06, 9.34482260742486e-06, 
    1.85998601467761e-06, 1.13981438004737e-06, 1.09907750765286e-06, 
    1.017448730238e-06, 4.01808140067848e-08, 8.12614373528839e-07, 
    1.65904124237599e-07, 6.39278974178569e-06, 2.39260415468279e-06, 
    4.73913902861878e-06, 1.06836308293685e-05, 1.36703132972357e-05, 
    2.33286024500832e-05, 2.43537343027982e-05, 3.67708964948827e-05, 
    4.38325460780656e-05, 5.54043928071728e-05, 5.5724041589132e-05, 
    3.69758666797254e-05, 2.372434300027e-05, 1.18484729400275e-05, 
    1.12468723947536e-05, 1.30442775555363e-05, 1.42013126286163e-05, 
    1.80259841336854e-05, 2.154646249564e-05, 2.01664414249208e-05, 
    2.54546752388908e-05, 3.38011219450552e-05, 6.53037806104312e-05, 
    7.16313106664362e-05, 6.56262858717275e-05, 5.9164297980608e-05, 
    5.13501381826877e-05, 6.77593279423231e-05, 3.75208734894965e-05, 
    2.24138002529703e-05, 3.98456061627081e-06, 1.41666367278401e-06, 
    2.03863446966359e-06, 0, 0, 0, 0.000196969478086502, 
    4.23424102129078e-05, 2.19437763532767e-06, 3.90763744954992e-07, 
    4.48226811648401e-06, 7.65816017418961e-06, 1.76614906577189e-05, 
    4.81305593952291e-06, 5.34880016391693e-06, 1.00137625124069e-05, 
    0.000145513913153486, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.73003488242418e-07, 
    1.31154968953709e-07, 4.3242900678806e-08, 2.16681925474532e-07, 
    4.93858569024871e-07, 4.94168021048321e-07, 0, 0, 0, 
    6.62944082894743e-06, 8.49419030985026e-07, 4.64555255725142e-06, 
    1.79787018468294e-07, 1.14968842254776e-06, 3.97452408087404e-06, 
    1.44199491320263e-05, 1.53649893371617e-05, 1.48762529463534e-05, 
    1.59970963209723e-05, 1.25999647978371e-05, 1.01180502465069e-05, 
    6.5966634585515e-06, 2.10261170335296e-05, 4.64478074303805e-05, 
    2.58453964463262e-05, 1.53931708950141e-05, 1.19594253359297e-05, 
    1.38159865825189e-05, 1.27751460871017e-05, 1.54976489655825e-05, 
    1.63885399948866e-05, 1.78184300879726e-05, 1.78727346145954e-05, 
    1.44004781237126e-05, 3.09880385334334e-05, 7.52092446623835e-06, 
    4.0151569450565e-07, 2.78302009290764e-06, 2.35924629200013e-06, 
    7.74582171139226e-06, 7.97598872939251e-06, 5.96531547215835e-06,
  2.54406015876995e-05, 2.4994020991672e-05, 1.79858839071164e-05, 
    1.63240215502741e-05, 1.80547471386483e-05, 2.40166301665894e-05, 
    2.36487662608824e-05, 2.20224386183992e-05, 2.67464608458594e-05, 
    1.85815302500495e-05, 3.54428136368707e-05, 5.38564254817353e-05, 
    4.09775367417804e-05, 3.46827674500641e-05, 5.80560155830359e-05, 
    4.2669630726658e-05, 5.59436052485072e-05, 8.9943540348297e-05, 
    2.95652838175625e-05, 4.12540944036568e-05, 2.60647533078967e-05, 
    3.5000192977718e-05, 3.5476196435028e-05, 2.74048661468995e-05, 
    1.11325627764079e-05, 1.0475056636872e-05, 1.08511016264965e-09, 
    1.4410493506541e-06, 3.22318326880546e-06, 1.66591497673863e-05, 
    1.79214026958417e-05, 3.09642779412076e-05, 1.00982796361512e-05, 
    4.19045807229718e-06, 2.30477172987414e-05, 0.000157374351065974, 
    7.4182946076282e-05, 1.1284023936051e-06, 5.24905459632118e-06, 
    6.5753744893008e-06, 4.8021825683199e-06, 2.97389556287588e-06, 
    4.83208674252834e-06, 8.41237016379573e-06, 1.09119975620691e-05, 
    1.41982018545005e-05, 8.84896937753043e-06, 1.94724702574909e-05, 
    3.02742324924636e-05, 2.53739079617557e-05, 4.15744904455523e-05, 
    5.72446093418177e-05, 5.70374510329838e-05, 6.94908516124792e-05, 
    6.63175885597701e-05, 7.35440425796724e-05, 5.51531366902186e-05, 
    2.39802905758268e-05, 6.84413375878111e-05, 8.59181742993784e-05, 
    6.82080992961724e-05, 2.90950822237167e-05, 1.16848707470643e-05, 
    4.16382295928332e-06, 2.35756139210397e-06, 4.21573217424382e-06, 
    1.26581296758147e-05, 3.33415138268955e-05, 3.72903213173261e-05, 
    8.01163422240326e-05, 6.72311093530647e-05, 7.71785616941286e-05, 
    7.06300447617253e-05, 6.92209044701049e-05, 4.29758145727125e-05, 
    2.44711081367138e-05, 3.75088770390219e-05, 0, 0, 0, 0, 0, 
    0.000126306451201048, 7.87934393749867e-05, 7.89305530864711e-07, 
    1.13068082695331e-06, 2.09263327787156e-06, 1.63545491734524e-05, 
    9.72980775859647e-06, 7.75508360592491e-06, 6.35664365916494e-06, 
    1.19827133864366e-05, 1.13971361057151e-06, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.79611920403974e-07, 0, 2.80314663826527e-06, 2.09810518776083e-06, 
    1.37641770800738e-06, 8.41689344006561e-07, 6.69192613428807e-07, 
    1.52214914078034e-07, 0, 2.12902526437127e-07, 2.35199534982284e-06, 
    5.24983629346882e-06, 5.91156056873588e-06, 5.31327787858255e-06, 
    1.75575828399287e-06, 9.54151956586585e-07, 3.39423510684817e-06, 
    7.25162998796316e-06, 8.73640004851104e-06, 7.69793997687295e-06, 
    7.91297878467119e-06, 4.43969324450188e-06, 1.88300027204984e-05, 
    1.76659396192032e-05, 1.14591667093456e-05, 8.27573930865495e-06, 
    2.01636181517811e-05, 2.29463507511123e-05, 3.08406125669337e-05, 
    2.13441495520898e-05, 1.13266466268003e-05, 5.71733448295295e-06, 
    1.13808257666177e-05, 1.13314443848801e-05, 9.65606277888937e-06, 
    8.27953428937635e-06, 4.0309883560463e-06, 5.12748840220261e-06, 
    3.11805613914146e-06, 4.18771995294782e-06, 4.11904344929976e-06, 
    6.78080632884105e-06, 1.47095223170244e-05,
  3.40710767233097e-05, 1.21955013126964e-05, 9.45260568691357e-06, 
    1.55565595765257e-05, 1.79027199147641e-05, 1.79306225575649e-05, 
    1.1293377707426e-05, 1.62153154673852e-05, 1.95090638828123e-05, 
    2.71726157866453e-05, 1.77922870829216e-05, 2.69974021465155e-05, 
    3.74355034840709e-05, 3.60633613709388e-05, 4.32680454379841e-05, 
    4.59947398365703e-05, 5.11640171946492e-05, 6.11033664820947e-05, 
    3.7093767924467e-05, 4.65026979915636e-05, 4.81022013521543e-05, 
    3.922006635475e-05, 4.03768307297477e-05, 3.17430943958159e-05, 
    8.41506038499045e-06, 5.4732036714926e-08, 1.37023551407967e-06, 
    5.14382497713137e-07, 0, 0, 0, 0, 0, 0, 0, 0.000144832309833647, 
    0.000172472864819653, 1.86896546946409e-06, 3.05996153777484e-08, 
    2.82062024264675e-06, 8.85266198741337e-06, 1.21411676661402e-05, 
    1.15989065918073e-05, 5.47567627559789e-06, 1.39046015553104e-05, 
    3.76246381437201e-05, 2.69484999969982e-05, 3.84893207519417e-05, 
    5.25516907515826e-05, 6.37140753651095e-05, 7.10046764087238e-05, 
    4.82920279673149e-05, 6.00181896315481e-05, 3.32174173847973e-05, 
    1.50543538035923e-05, 1.27950747196947e-05, 6.74085469640214e-06, 
    1.78717363303569e-05, 1.22712857772093e-05, 0, 0, 3.21593481004825e-08, 
    0, 5.26023018252708e-06, 4.07864306295162e-06, 4.50741312111418e-06, 
    4.64206739747876e-06, 5.9238519060089e-06, 2.48471349673792e-05, 
    3.45843475702989e-05, 3.81865312077113e-05, 7.01505548766318e-05, 
    6.1246924454523e-05, 4.76407480584243e-05, 6.5640651330846e-05, 0, 0, 0, 
    0, 0, 0, 0, 0, 8.31210236009149e-05, 8.96510114203856e-07, 
    6.18483960015657e-06, 5.28744891510383e-06, 7.64556131321241e-06, 
    1.20926748919792e-05, 7.43732534517717e-06, 9.0051708451927e-06, 
    1.59517935510774e-05, 0, 0, 0, 0, 0, 0, 0, 0, 9.4942382673643e-07, 
    8.97653610159176e-07, 7.45109102669588e-08, 1.15937395110541e-06, 
    1.38107410660083e-06, 4.87820672408472e-06, 4.74710758475118e-06, 
    5.83802985399571e-06, 4.44997107384827e-06, 0, 0, 0, 
    1.06089781824069e-05, 9.11543139081127e-06, 7.73454929165731e-06, 
    7.77673623345587e-06, 6.58452630603091e-06, 1.51186870627928e-05, 
    6.89315386238283e-06, 8.07530112315318e-06, 1.69756445068991e-05, 
    8.67586151712576e-06, 2.1484286347404e-05, 8.83153288522283e-06, 
    4.77482819048549e-06, 1.38782426298723e-05, 7.60467655313399e-05, 
    0.000108629631312457, 9.7887208507685e-05, 0.000153546957997988, 
    0.000162780714989192, 0.000132314389194757, 3.34846448291315e-05, 
    9.70140274933255e-06, 9.45326687262067e-06, 6.13045979080999e-06, 
    3.96331705579616e-06, 4.37671838288727e-06, 6.2596932552236e-06, 
    4.53430730655095e-06, 3.79440748315158e-06, 8.664844511288e-06, 
    1.24962534122981e-05, 1.8914059132129e-05,
  8.25011788066986e-06, 1.06215069136554e-05, 4.88058373083411e-06, 
    8.44766758888839e-06, 9.06059426857081e-06, 1.42579777414772e-05, 
    1.56540508138404e-05, 1.63805183052856e-05, 1.33429303120198e-05, 
    2.14264014858661e-05, 1.09253110582776e-05, 1.49267561650075e-05, 
    2.36493718842149e-05, 2.49400779424204e-05, 3.08158874031912e-05, 
    5.0953817837829e-05, 4.42063372925553e-05, 2.74108408446482e-05, 
    2.91415324647646e-05, 3.7700438133774e-05, 5.56927488204597e-05, 
    5.58969124903437e-05, 2.06036697840267e-05, 1.48857133634128e-05, 
    6.80890880719968e-07, 1.11908378000758e-06, 9.51996223322843e-08, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.00017450538632408, 2.18400007498623e-06, 
    3.95695939292236e-07, 4.3120893995103e-06, 7.64745819492358e-06, 
    7.86227217304881e-06, 1.61002859851414e-05, 2.96052513138135e-05, 
    2.94052517455453e-05, 1.59342229334814e-05, 4.81408285401894e-07, 
    2.95460062993131e-05, 3.68210723181314e-05, 5.11805146404098e-05, 
    6.89338627589029e-05, 5.03590635475393e-05, 1.36970147360387e-05, 
    3.24697777469381e-07, 2.04166783161065e-06, 4.67908274843475e-06, 
    1.12220774549127e-05, 0, 0, 0, 0, 0, 0, 1.202396101382e-05, 
    5.23273259489365e-06, 8.70661456509618e-06, 1.49622031526767e-05, 
    2.23785576134055e-05, 3.56069065971719e-05, 3.4506958105578e-05, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.53538677143065e-07, 
    5.06832384511424e-07, 1.38597227221785e-05, 2.18806331541369e-05, 
    2.4013025887262e-05, 1.14760850740136e-05, 7.0645930896122e-06, 
    9.71870345495131e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.96907815480166e-07, 
    2.54765618697273e-07, 1.96829673113455e-07, 2.19157622815631e-07, 
    6.65611409918195e-07, 1.89448723722541e-06, 1.56371164929989e-06, 
    3.15359691910045e-06, 0, 0, 0, 0, 0, 2.53307722687099e-05, 
    2.31428137353757e-05, 1.56620490139244e-05, 1.52637729964997e-05, 
    1.13037120001277e-05, 8.8313158224852e-06, 1.39011763226247e-05, 
    1.30301187299833e-05, 2.0392476474683e-06, 4.70141104463229e-06, 
    2.59121056466704e-06, 1.85499659981215e-06, 0, 0, 0, 0, 
    1.70197311502608e-07, 0, 0, 0, 5.46685392173029e-07, 
    2.51041358856358e-06, 3.16533590965834e-06, 3.04643125836139e-06, 
    3.91002999876719e-06, 4.46969237439838e-06, 3.80862161805997e-06, 
    4.68166143593355e-06, 3.08221956256678e-06, 6.69305912427446e-06,
  0.000179973621762878, 0.000209548950718559, 0.000173968708168649, 
    1.39295251548777e-05, 1.5527388828415e-06, 2.72459730625607e-06, 
    6.13299080724721e-06, 6.4729845900969e-06, 9.28565056384187e-06, 
    1.0412928346027e-05, 1.12806403412908e-05, 1.14438827792256e-05, 
    1.07793277719414e-05, 1.91987587954116e-05, 3.49411614759922e-05, 
    4.8429342260479e-05, 3.11100622415393e-05, 3.28378222629193e-05, 
    2.28732219110788e-05, 2.04249521055359e-05, 1.43765730314748e-05, 
    1.21561338087284e-05, 3.20131233702912e-06, 0, 4.55359188898855e-07, 
    1.90890645972302e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.6322047632234e-07, 
    8.14378695003711e-05, 2.99775833557716e-08, 3.47893554585666e-07, 
    5.18483332198352e-06, 1.1518870615067e-05, 3.62627001961828e-05, 
    3.83581991687707e-05, 3.15013459615459e-05, 1.67279794029296e-05, 
    2.78556899537384e-05, 3.31846339457686e-05, 3.35161355883889e-05, 
    2.50354353430525e-05, 1.60962994384962e-06, 0, 1.94379734760389e-07, 
    2.49738648169534e-05, 3.75079263311655e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.8305576990262e-07, 1.11357075905056e-06, 9.7473253138873e-06, 
    1.70414034904572e-05, 3.08683207148241e-05, 3.63435121172409e-05, 
    2.1786505694042e-05, 1.75917781832342e-06, 6.99289547479869e-06, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 9.21149438358073e-07, 1.05211420883205e-07, 
    2.21682660949816e-07, 5.12523730051155e-08, 1.46707445437933e-07, 
    1.53523237357856e-06, 1.10915672302718e-06, 2.10536995596735e-06, 
    7.04024513615911e-06, 0, 0, 0, 0, 2.58808889688268e-05, 
    1.82639973910734e-06, 6.0288260635073e-06, 3.54712871794014e-05, 
    5.08854827950176e-05, 3.00470411378038e-05, 2.56648076365709e-05, 
    2.07707947175671e-05, 4.04079286071899e-06, 1.24273143193903e-05, 
    7.131166914682e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.72777599223658e-06, 
    4.90972809875552e-06, 1.54375446686443e-06, 5.37487315410452e-06, 
    4.74627094638898e-06, 3.01599502071125e-06, 4.06323012136394e-06, 
    6.58001751435561e-06, 8.15097666196001e-05,
  0, 0, 0.000191827432240907, 0.000272622839900728, 3.41247506470459e-06, 0, 
    2.63235933259534e-06, 1.90505958540022e-06, 2.0647463733977e-06, 
    3.07652441512908e-06, 8.68952289451182e-06, 1.21958769452424e-05, 
    2.28585339034798e-05, 1.85916274966228e-05, 3.13574728838086e-05, 
    2.19643104848913e-05, 1.80861023271339e-05, 1.43500463857487e-05, 
    2.07381604694494e-05, 1.2681440380858e-05, 6.23287619645518e-06, 0, 
    1.92242718356057e-06, 3.00346253623629e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3.18503142370748e-06, 1.96711097133023e-06, 
    2.56283026110489e-06, 8.35081715133123e-06, 2.51554398330479e-05, 
    4.09018339634481e-05, 3.88953444664524e-05, 3.42933216610483e-05, 
    2.01066852282385e-05, 4.05621930800968e-05, 3.73775185714418e-05, 
    3.73642913528868e-05, 5.70045009425814e-06, 0, 1.34618181856586e-05, 
    2.59278811661803e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7.11878629522725e-06, 
    1.02339221666848e-05, 1.23211346372908e-05, 2.72237973636298e-05, 
    3.68293524783275e-05, 2.49346085130637e-05, 1.88838120341456e-05, 
    4.17721498271179e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.81700505722487e-07, 2.39211112269011e-06, 9.28729656321493e-07, 
    2.71718374473575e-07, 5.67877055293289e-08, 1.8382420877918e-06, 
    5.098032029796e-06, 5.96808485953891e-06, 0, 0, 0, 0, 4.167827332016e-06, 
    0, 2.18239244731299e-05, 5.05253276526972e-05, 4.8906315737841e-05, 
    3.71561029386241e-05, 1.51371916201769e-05, 9.03151168931121e-06, 
    8.21986676587191e-06, 1.06023664854343e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 9.73622185257484e-08, 6.18544523662487e-07, 3.50632624188905e-08, 
    5.25619275073924e-07, 2.35488686410606e-06, 2.79380253999946e-06, 
    1.36741675133109e-05, 8.41732425439315e-07, 0,
  0, 0, 0, 5.42995439091253e-07, 0.000209723648024664, 6.80901320082329e-06, 
    3.23009186757905e-06, 0, 1.56208096638553e-07, 2.12309500720281e-06, 
    4.51088145317754e-06, 1.21297021147765e-05, 1.08201034967524e-05, 
    2.82500593564257e-05, 2.36870882798705e-05, 2.42130799442814e-05, 
    2.00046752775852e-05, 1.04581711090263e-05, 8.96184854831579e-06, 0, 0, 
    3.64765680773665e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9.97246476840707e-06, 6.79638164492383e-06, 4.97818421038954e-06, 
    1.30556824017466e-05, 3.45325905530381e-05, 3.35756501941898e-05, 
    3.37175040690631e-05, 4.2042347801768e-05, 3.85868305613595e-05, 
    3.85665345602094e-05, 4.9095106813951e-05, 6.51578224403876e-06, 
    9.59098010406231e-06, 2.92827921197137e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.54757500861914e-05, 1.38081592762227e-05, 1.36780008434344e-05, 
    3.52665776624611e-05, 3.92865808662158e-05, 3.22242039604724e-05, 
    2.76860086769832e-05, 5.30416583432104e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1.10065085072048e-07, 3.45227407037383e-07, 2.96396922046823e-07, 
    2.76711764582466e-07, 2.71264389757606e-07, 6.98244701797393e-07, 0, 0, 
    0, 0, 2.51543960800698e-05, 5.02944641086376e-05, 2.18780819779629e-05, 
    0, 4.99264401803451e-05, 6.43480102654569e-05, 2.00445195150072e-05, 
    8.59536130241756e-06, 9.01415956148029e-06, 1.76017963710295e-05, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9.64061308257497e-07, 
    1.83159919242379e-06, 2.66016660001181e-06, 2.24713551386042e-06, 
    5.32031199070559e-06, 1.02754156131382e-06, 0,
  0, 0, 0, 0, 6.21686569518483e-06, 1.23082334321488e-05, 
    5.44920742087992e-07, 1.10104571875141e-07, 2.41550751226049e-07, 
    1.00569416140159e-06, 4.05919881935509e-06, 1.71407999825278e-05, 
    5.67662882154574e-06, 2.58097970177075e-05, 2.67203077992554e-05, 
    2.12006335090245e-05, 1.88735820714653e-05, 8.29599226549553e-06, 0, 0, 
    5.52469595113432e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.06890916613614e-05, 1.70379432214913e-05, 5.09537695062909e-06, 
    1.86820919186712e-05, 3.61970745247319e-05, 3.59449357619719e-05, 
    5.63009286274989e-05, 7.87369525075377e-05, 5.66765078597021e-05, 
    5.75504169376327e-05, 1.96512552513842e-05, 1.34293843685737e-05, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2.48972515579561e-05, 1.20875442537918e-05, 
    3.79213372083083e-05, 4.74042992030797e-05, 3.66159042365918e-05, 
    1.80291150341398e-05, 4.94001606722775e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1.27772037504187e-09, 1.48812214541997e-07, 
    4.2479463145904e-07, 0, 0, 0, 0, 0, 0, 6.54537715412643e-06, 
    1.22872660133819e-06, 0, 4.76918515720944e-06, 8.62711269440367e-05, 
    3.04531877001092e-05, 8.01035868009082e-06, 1.6236221164087e-05, 
    5.37592080593616e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4.02820396387089e-07, 1.40678199285817e-06, 3.87390898910451e-06, 
    1.05125449248266e-05, 6.47033588843146e-06, 0,
  0, 0, 0, 0, 0, 8.55200933572225e-06, 1.31448741362783e-06, 
    5.84752947820045e-07, 5.76192919614958e-07, 2.74347504051755e-06, 
    3.41028209197186e-06, 6.81655511636891e-06, 1.78529162490882e-05, 
    2.00227292007659e-05, 2.21586232426235e-05, 1.6640069141465e-05, 
    5.40903026835126e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1.73461891737545e-05, 1.33133800773399e-05, 
    1.14084245890186e-05, 2.49913749733695e-05, 2.97982958363701e-05, 
    0.000107761321656287, 0.000191268125586377, 8.45244788889913e-05, 
    2.61402915814881e-05, 2.03751983224608e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 2.50635039401885e-05, 2.87593251557526e-05, 3.94461701219153e-05, 
    3.21265019665879e-05, 2.92678650193004e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.16330750858159e-05, 
    1.13817264507779e-07, 9.346104098842e-07, 3.42173135741206e-06, 
    5.51567048272638e-05, 4.80524235740529e-05, 2.29309219793832e-05, 
    1.78121063194454e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.31207934501034e-06, 6.50852646249466e-06, 1.8796744168046e-05, 
    1.03141689143205e-05, 0,
  0, 0, 0, 0, 0, 0, 2.52629395913784e-06, 1.26977083061225e-07, 
    3.22098661983495e-07, 3.08559348413733e-06, 6.15793954984939e-06, 
    1.21257725963429e-05, 1.46346196824819e-05, 2.60346901336779e-05, 
    2.41066212895309e-05, 1.28645835145798e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.14709474744481e-05, 
    1.32683408452677e-05, 3.56071868294402e-05, 9.55330763738701e-05, 0, 
    7.97465127871369e-05, 2.0188789698881e-05, 1.8001574729269e-05, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.25901677474257e-05, 
    2.84411485480709e-06, 5.24525744933841e-06, 2.16120302195711e-07, 
    3.14817954628504e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 4.64774821272692e-06, 1.56117158417684e-06, 
    2.91421501285691e-06, 7.26728596911949e-06, 9.56367588801073e-06, 
    3.20090048082397e-05, 4.01281639292047e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.16239880234781e-05, 4.69029571769431e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.36968770582072e-05, 4.84831912892634e-06, 
    5.75384032907259e-06, 4.29310864059435e-08, 3.58727276549854e-06, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.04369321287433e-05, 
    8.11286694450742e-08, 4.41337058105951e-06, 2.37211487231815e-06, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6.18601092480298e-09, 7.92662818306066e-07, 9.78259403017388e-07, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.08685990068268e-05, 1.0338831170552e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 1.13712995611852e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.85781180688718e-06, 9.73199861561153e-06, 1.06236972368015e-05, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 9.97063217498753e-08, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1.97496499207386e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 3.63517774745988e-10, 1.66469131757289e-07, 
    3.06900055883847e-10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.83440662049897e-05, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.68901374779447e-10, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8.3594112450324e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.71909708306387e-05, 4.84681886864735e-06, 
    2.63526128506828e-06, 5.43946095779861e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 3.65198974686367e-09, 0, 0, 0, 2.55316417494151e-05, 
    3.90034896938872e-05, 3.33626317152178e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2.06551097151097e-09, 2.54787918897865e-06, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8.11045909087162e-06, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.86355914757527e-06, 7.23532495641103e-08, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5.68579367968944e-07, 1.18772674942394e-06, 1.81062763850303e-06, 0, 
    6.30600492374012e-09, 0, 0, 0, 0, 0, 1.67473345148838e-06, 
    3.16244429025617e-06, 3.44020536969159e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6.10443948311507e-07, 0, 4.82096170884795e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4.51836594765418e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.38164511488313e-07, 0, 0, 0, 7.59114582704576e-12, 
    4.69725504754114e-12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3.74572150365194e-06, 5.21759033473113e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1.67264773875341e-06, 8.64353361846325e-07, 
    1.69540759614651e-06, 0, 0, 2.33096438494365e-06, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1.11989261305424e-05, 1.62257759299853e-05, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 6.33953794222713e-08, 1.19347034443097e-07, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5.90394069090334e-07, 2.57343480093266e-06, 5.57944622728901e-06, 
    9.37163882904109e-07, 1.62921489819292e-06, 0, 4.16378721708804e-06, 
    3.14326480822256e-06, 0, 7.60302466489058e-06, 0, 3.11724374794974e-07, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.41473498151444e-10, 
    1.34452327117693e-08, 2.71346938033341e-10, 0, 0, 0, 0, 0, 0, 
    7.75925204845647e-09, 3.14242076041947e-07, 1.21085374476913e-09, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.75735411714454e-06, 
    2.34287815026196e-06, 1.8758138119651e-06, 1.96884980548296e-06, 
    1.59524545057704e-06, 1.6277752529033e-06, 2.43607710839475e-06, 
    4.19233129742698e-06, 3.59957434881826e-06, 9.77090261878909e-06, 
    1.89436731214092e-06, 6.6809585353228e-07, 1.47137700281571e-06, 
    1.90924304463702e-06, 1.04795697975941e-05, 5.79422000332082e-06, 
    9.20323449869043e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1.12375258907027e-07, 0, 0, 0, 0, 0, 0, 4.83387131007777e-09, 
    8.40326565307696e-07, 2.14844529047404e-06, 3.31035165827581e-08, 
    1.21163836286665e-11, 0, 0, 0, 0, 0, 0, 7.53839347867344e-09, 
    1.38499788854371e-07, 1.55234523645567e-07, 0, 0, 0,
  5.55771479482883e-07, 1.87423949836997e-06, 1.12255802345685e-06, 
    8.14672922288628e-07, 1.61766545974479e-06, 1.16346079839973e-07, 
    1.19500317399043e-06, 1.33895779310588e-06, 0, 0, 1.8488123389793e-06, 
    5.68709954237665e-07, 3.40876526479232e-06, 2.57972812372011e-06, 
    1.37978854304867e-07, 3.28085673951823e-06, 1.96725859426783e-06, 
    3.48757802959569e-06, 3.83998095236306e-06, 6.26523384953079e-06, 
    5.87177785475132e-06, 1.5785601378837e-05, 1.65526851082951e-05, 
    3.11895529787375e-05, 6.9944952514389e-06, 2.77690035961409e-06, 0, 0, 
    8.79506113167963e-07, 0, 1.29677122267941e-08, 0, 0, 0, 
    4.36643142730547e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1.75363584850787e-09, 1.68516532870581e-06, 2.84723556715593e-06, 
    3.26724284560885e-06, 3.13607052841115e-07, 1.14306325397115e-09, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4.082807596349e-09, 6.21039842562306e-07, 
    1.03318757423385e-06, 2.81482194770936e-06,
  2.44555884718596e-07, 3.13465189839946e-07, 2.80851761189466e-06, 
    1.90075421466268e-06, 1.90375042535315e-06, 6.21643638134231e-07, 
    1.29294883789469e-08, 1.33376716845716e-10, 1.03669975022799e-08, 
    1.36567059003684e-07, 5.3750897538048e-09, 1.0993838519024e-09, 
    4.63554106143367e-07, 4.11310674961054e-06, 4.27136967964315e-06, 
    1.6468625017065e-06, 3.19645095740399e-06, 8.98521232180811e-06, 
    7.954945198483e-06, 1.51643338126393e-05, 7.29931131743812e-06, 
    2.05107622022063e-06, 5.78714310967077e-06, 6.7315283668536e-06, 
    1.35362268268774e-05, 9.88993051072126e-06, 1.94857364143705e-06, 
    1.42876634100596e-07, 1.2238018813103e-06, 9.46541108624934e-07, 
    9.92325158173772e-07, 3.74121881776992e-06, 4.11866288765941e-06, 
    3.0015942043202e-06, 2.37568016379244e-06, 0, 9.99918740980637e-08, 
    1.30132969792999e-07, 3.33374100593916e-06, 1.58565177809577e-07, 
    2.53258264466676e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 7.51443305301035e-10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 7.32200478083404e-12, 6.20728670966182e-09, 3.30768474420995e-09, 
    4.87162864830055e-11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3.87838677350531e-07, 7.28261785873129e-06,
  1.29104749368316e-06, 1.48854101225037e-06, 4.45496282470147e-06, 
    1.5971563524041e-05, 1.44831504120897e-05, 7.01933517273474e-07, 
    3.09573324015649e-07, 1.12764487274817e-07, 1.27271424911004e-07, 
    1.57155193291513e-07, 3.88342287250441e-07, 4.47525109518002e-06, 
    4.45732855956573e-06, 6.79269226926199e-06, 7.43649170146939e-06, 
    8.26625899429596e-06, 1.15260946221759e-05, 1.37741990779392e-05, 
    1.06432490053753e-05, 1.4000585166649e-05, 4.78518409856704e-06, 
    3.6165713645439e-06, 4.75670118637198e-06, 5.65915237234425e-06, 
    1.08246659228085e-05, 5.68156982871795e-06, 5.91703769190685e-06, 
    2.94141305928236e-06, 2.54634167452541e-06, 7.86851483439012e-06, 
    7.38783005084901e-06, 6.21954757243415e-06, 5.53326615932056e-06, 
    6.26223074605106e-06, 3.76529420358936e-06, 2.57124041198007e-06, 
    5.61901895514895e-06, 6.77247095816918e-06, 9.37595702216135e-07, 
    1.92576206577514e-06, 3.75551464389612e-06, 1.79107539202148e-06, 
    1.34973909819059e-06, 5.75075801475006e-08, 1.03178578350143e-08, 
    8.76281669424563e-07, 5.61324250227465e-07, 5.10016480536388e-07, 
    1.15502241731307e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.72478240390166e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6.31572288140416e-13, 5.33327429298233e-12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 1.72798213753833e-06, 3.1222272850214e-06, 6.53765575340113e-06, 
    6.26394209397733e-06, 5.7231447569049e-06, 3.34322487942096e-06, 
    1.84787761225545e-06, 2.62376477475069e-06, 3.65313520500028e-06, 
    4.59285963615587e-06, 1.18927232179664e-05, 1.17649263797921e-05, 
    1.48636914962541e-05, 1.82667586204294e-05, 2.20083974768911e-05, 
    2.70890000882114e-05, 2.90316969706909e-05, 3.08880978133474e-05, 
    3.06792900978525e-05, 3.31787916793752e-05, 2.91234704966145e-05, 
    2.8154711347085e-05, 2.37745947616023e-05, 2.20702589097132e-05, 
    1.54985404292992e-05, 1.09882707755421e-05, 8.45200804687647e-06, 
    5.83507518522708e-06, 3.76763899927703e-06, 3.70187542405111e-06, 
    5.261353969812e-06, 5.85977901621117e-06, 5.58534236459679e-06, 
    6.2637859881485e-06, 5.67568591938441e-06, 2.37585233565444e-06, 
    2.15561295363079e-06, 1.21617264929709e-06, 1.93367818289229e-06, 
    2.30062330527909e-06, 4.514642177212e-07, 0, 0, 0, 0, 0, 0, 0, 
    6.29954252857093e-07, 3.47713513128259e-06, 3.66349809662721e-06, 
    1.9577918564311e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.40255191351654e-06, 
    1.43867389359018e-05, 1.49488985642874e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 1.96594701177759e-06, 1.71853669387856e-06, 2.0201327262617e-06, 
    1.81836257844126e-06, 5.70029881841053e-06, 4.93323501020486e-06, 
    4.02815906609961e-06, 7.46803637572682e-06, 1.17318261090968e-05, 
    2.17219536634435e-05, 3.14816480224757e-05, 3.73838706677092e-05, 
    3.93206952219211e-05, 4.1242816673163e-05, 4.47156229216281e-05, 
    4.73907060839237e-05, 4.68412898246044e-05, 4.5470996092124e-05, 
    4.25127459765386e-05, 4.13934508276961e-05, 4.09479826537531e-05, 
    4.09811988640267e-05, 4.17959526274152e-05, 4.17087978674762e-05, 
    4.16836920915324e-05, 4.1315703889067e-05, 4.0595025874464e-05, 
    3.88781175693148e-05, 3.63545872429915e-05, 2.9572047783812e-05, 
    2.531815342529e-05, 2.15590352792247e-05, 1.55387015872328e-05, 
    9.21262608676566e-06, 1.2723132493446e-06, 1.83121998173514e-07, 
    2.93264979861518e-07, 9.12463799164907e-07, 1.65106100534634e-06, 
    2.89519857615692e-06, 2.34041727413205e-06, 1.19500611724679e-06, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.55066949834253e-07, 
    5.37036920702981e-06, 1.14730743188933e-05, 2.26243860677788e-05, 
    4.17413683064085e-05, 0, 0, 0, 0, 0, 0, 6.76088941689098e-11, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 9.48294321899381e-07, 2.47773155308567e-06, 0, 
    2.43429356149109e-06, 8.43800240977118e-06, 1.29383175396791e-05, 
    2.18836325642796e-05, 3.05981754025856e-05, 3.72019034705842e-05, 
    4.08387125502557e-05, 4.3390970577973e-05, 4.6148735157077e-05, 
    4.70476124975595e-05, 4.52862047738711e-05, 4.35929429896747e-05, 
    4.3451584718346e-05, 4.05466308572375e-05, 3.82797219261965e-05, 
    3.58104451798311e-05, 3.29516036936922e-05, 3.04929209650821e-05, 
    2.88261485685208e-05, 2.84746196123105e-05, 2.86430343202586e-05, 
    2.87062072664865e-05, 2.87350060717239e-05, 2.63647942883151e-05, 
    2.6207609597552e-05, 2.60561326141201e-05, 2.51927193862623e-05, 
    2.32388713321967e-05, 1.99339507133211e-05, 1.55038184967441e-05, 
    1.17329467607607e-05, 1.19070794609963e-05, 8.43137432584675e-06, 
    9.96012729802185e-06, 5.68173740003919e-06, 2.36076845312182e-06, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.34587419578136e-06, 
    5.69965434239675e-06, 1.061203816581e-05, 1.69159619668035e-05, 
    3.00786655953525e-05, 5.02233771298978e-05, 6.27075032297412e-05, 
    6.20204463461029e-05, 0, 0, 7.39693263146569e-10, 0, 0, 0, 0, 
    1.60112378023589e-10, 1.02301630599617e-09, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 1.11351503310011e-05, 2.4583979409893e-05, 
    3.15005192236713e-05, 3.81727024858001e-05, 4.74424181430072e-05, 
    5.61118855420191e-05, 6.32055858673487e-05, 6.75355624210729e-05, 
    7.06619799622631e-05, 6.50925224920352e-05, 6.42434553891323e-05, 
    6.7680902670057e-05, 5.85190369846714e-05, 6.02572816606957e-05, 
    6.01076264306371e-05, 5.46019615200309e-05, 5.22057493782202e-05, 
    4.94013961283402e-05, 4.43025615986506e-05, 3.83625775131669e-05, 
    3.22662437896279e-05, 2.76009635098834e-05, 2.44480985350999e-05, 
    2.20505525254774e-05, 2.00828430795519e-05, 1.84948002709867e-05, 
    1.71304986480441e-05, 1.57647608609056e-05, 1.45938109945346e-05, 
    1.3490762666059e-05, 1.24340521960976e-05, 1.19707411049207e-05, 
    1.14674883128258e-05, 1.12058059367871e-05, 1.09826624180809e-05, 
    1.07007273367814e-05, 1.05917164567455e-05, 1.03027186370653e-05, 
    1.00218160975844e-05, 9.79153001601763e-06, 9.65386771250605e-06, 
    9.19604965809228e-06, 8.90983026270066e-06, 8.76257121524582e-06, 
    8.95265090558398e-06, 9.97912410609202e-06, 1.15805714362692e-05, 
    1.40745705988115e-05, 1.73221169773632e-05, 2.13945272396022e-05, 
    2.6267866164633e-05, 3.27358960573571e-05, 4.06617790434764e-05, 
    4.93167280545525e-05, 5.68101928778169e-05, 6.06569406346937e-05, 
    6.27374933582179e-05, 5.86931427905157e-05, 4.93833987719731e-05, 0, 0, 
    0, 5.30043393892382e-09, 2.1297969164289e-07, 6.34754646990446e-07, 
    1.41543045686271e-08, 9.76938294476058e-10, 2.45988705235689e-10, 
    3.29223433343155e-09, 3.30925428716215e-09, 2.73205268857712e-09, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 1.26905851994172e-05, 1.82864440254873e-05, 
    2.10724595177316e-05, 2.311716734893e-05, 2.49580793800734e-05, 
    2.78002404856106e-05, 3.05713944481749e-05, 3.01427197434457e-05, 
    2.98751498451917e-05, 3.73649487452034e-05, 3.74334976033519e-05, 
    4.04794750291522e-05, 4.50877422822633e-05, 4.48974492566892e-05, 
    4.83726461085962e-05, 5.04919167377237e-05, 5.04383893307887e-05, 
    5.15784161126256e-05, 5.21424764095868e-05, 5.27659559347304e-05, 
    5.24226979782688e-05, 5.18067826176096e-05, 5.08029623037956e-05, 
    5.03503048101254e-05, 4.99704711857853e-05, 4.89450121297934e-05, 
    4.72622866204359e-05, 4.54002672273402e-05, 4.31678375778659e-05, 
    4.12773665149168e-05, 3.97425451350095e-05, 3.83114559880874e-05, 
    3.70745659065362e-05, 3.56598890891018e-05, 3.42516303684351e-05, 
    3.25789419014906e-05, 3.20127917670954e-05, 3.18568017672027e-05, 
    3.13676231815808e-05, 3.02379035792375e-05, 2.94411713480579e-05, 
    2.84331294034964e-05, 2.71526352232925e-05, 2.5273120490862e-05, 
    2.37248264070968e-05, 2.18623686752944e-05, 1.99909031412775e-05, 
    1.91239998099432e-05, 1.8341343297084e-05, 1.83178033805505e-05, 
    1.71530628730044e-05, 1.57452118805708e-05, 7.47841525570602e-06, 
    6.29589955253512e-06, 3.93389384593544e-06, 4.39257906113496e-06, 
    1.13271574331051e-06, 4.05071568033686e-07, 1.06149780536332e-08, 
    6.55574105822885e-09, 4.6776433331171e-09, 2.28747569173126e-08, 
    1.31578470648105e-06, 3.96471272110296e-08, 2.32155970715148e-09, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  1.47234229453943e-05, 1.47235447128106e-05, 1.47236489179419e-05, 
    1.47237402112704e-05, 1.47238059428397e-05, 1.47238380125672e-05, 
    1.47238373274568e-05, 1.47237961561524e-05, 1.4723707413217e-05, 
    1.47235537023291e-05, 1.47233655171609e-05, 1.47231627134321e-05, 
    1.47228983619961e-05, 1.47225985330654e-05, 1.47222840227148e-05, 
    1.47218730147211e-05, 1.47214511167197e-05, 1.47209907288132e-05, 
    1.47204778592627e-05, 1.47199899151651e-05, 1.47194126470319e-05, 
    1.47187932078134e-05, 1.47181667305983e-05, 1.47175023435023e-05, 
    1.47168202535179e-05, 1.47161204042277e-05, 1.47153981451714e-05, 
    1.47146609608766e-05, 1.47139075974292e-05, 1.47090108523382e-05, 
    1.47037743417702e-05, 1.46992877304034e-05, 1.46954314037796e-05, 
    1.46926776798372e-05, 1.46909051577129e-05, 1.46899332319629e-05, 
    1.46899262274678e-05, 1.4690830355962e-05, 1.46925366814559e-05, 
    1.46950310724014e-05, 1.46981783930846e-05, 1.47017643211482e-05, 
    1.47030938502441e-05, 1.47023517891346e-05, 1.470161453045e-05, 
    1.47008872864505e-05, 1.47001675670559e-05, 1.46994505914013e-05, 
    1.46987396918944e-05, 1.46980351718653e-05, 1.46973383295982e-05, 
    1.46966497279847e-05, 1.46959699283581e-05, 1.46952969775141e-05, 
    1.46946301311203e-05, 1.46939748974732e-05, 1.46933329553875e-05, 
    1.46927028512097e-05, 1.46920865116603e-05, 1.46914870529621e-05, 
    1.46909070608586e-05, 1.46903495671857e-05, 1.46898215505695e-05, 
    1.46859383587251e-05, 1.46800973937243e-05, 1.46746712228833e-05, 
    1.46699054061821e-05, 1.46657727806351e-05, 1.46622806797989e-05, 
    1.46596629620094e-05, 1.46580054843235e-05, 1.46573917995258e-05, 
    1.46577790196352e-05, 1.46592780173377e-05, 1.46615074891595e-05, 
    1.46630953443566e-05, 1.4664948813946e-05, 1.46674720212564e-05, 
    1.46709509081819e-05, 1.46753391531981e-05, 1.46791956085731e-05, 
    1.46831574663737e-05, 1.46875328700167e-05, 1.46878501420574e-05, 
    1.46881893439414e-05, 1.46885471884185e-05, 1.46889190742489e-05, 
    1.4689308683023e-05, 1.46897125841813e-05, 1.46901251786897e-05, 
    1.46905489537739e-05, 1.46881385953174e-05, 1.4680720507951e-05, 
    1.46736545292915e-05, 1.46669378394539e-05, 1.46603216567285e-05, 
    1.46533841429267e-05, 1.4645711202229e-05, 1.46376516136643e-05, 
    1.46289805909787e-05, 1.46213888857726e-05, 1.4615370405963e-05, 
    1.46108246068224e-05, 1.46072629671825e-05, 1.46047570243133e-05, 
    1.46033181286458e-05, 1.46034885507558e-05, 1.46048330259612e-05, 
    1.46072530370125e-05, 1.46105238586876e-05, 1.46147096206797e-05, 
    1.46206064130903e-05, 1.46281842563422e-05, 1.46379626747127e-05, 
    1.46496084251291e-05, 1.46615630307304e-05, 1.46729822446765e-05, 
    1.46836938989442e-05, 1.46939377407905e-05, 1.47032355245451e-05, 
    1.47116911245278e-05, 1.47129461544002e-05, 1.47137221588189e-05, 
    1.47144734233938e-05, 1.47151994111322e-05, 1.4715891325683e-05, 
    1.47165605109972e-05, 1.47171985402458e-05, 1.47178089185045e-05, 
    1.47183887599986e-05, 1.47189388298427e-05, 1.47194562026783e-05, 
    1.4719943468669e-05, 1.47204017286293e-05, 1.47208267555137e-05, 
    1.47212059958342e-05, 1.47215552795994e-05, 1.47218770809063e-05, 
    1.47221685312707e-05, 1.47224337494845e-05, 1.47226804836047e-05, 
    1.47229059551994e-05, 1.47231045214517e-05, 1.47232761649076e-05 ;

 gust =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.567520903586482, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.863923707191847, 0.733756783813976, 0.630804239020818, 
    0, 0, 0, 0, 0, 0.591712633423921, 0.622572206746877, 0.489097611927072, 
    0.348688489556893, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.583725301415489, 
    0.69301312657212, 0.392250163664805, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.286063969132462, 0.797307383268872, 
    0.833990727387383, 0, 0, 0, 0.596598360408889, 0.720468191688168, 
    0.8341318336326, 0.770034042730103, 0.600806573363008, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.647936207045712, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.8491476505816, 0.69857974158234, 
    0.633530610183037, 0.472758741609529, 0.409753387455471, 
    0.450877716591415, 0.537982719301844, 0.599147099831206, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.546176444612319, 0.931905034348861, 
    0.446569821815951, 0.932191751589279, 0, 0, 0, 0.708513634638037, 
    0.549200411354417, 0, 0, 0, 0, 0, 0, 0.261046516749979, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.807128170794421, 0.907660466269717, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1.12760033787957, 0.992771058177099, 0.441686940425401, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.597860048078992, 
    0.715886586333908, 0.890141348583863, 0.779023149677981, 
    0.824206739916134, 0.8099627302914, 0.771188945680824, 0.737617974930202, 
    0.722018115935177, 0.590279967700368, 0.444804805469234, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.72341065561004, 0.76245455390988, 0.909626912495379, 
    0.851595165668342, 0.805872663831493, 0.178646003559317, 0, 0, 0, 0, 
    0.601873926263921, 0.813270437071572, 0.740794660746859, 
    0.448907610205172, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.669001769030734, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.987262513201857, 1.39519914600157, 
    0.846034373420577, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0.417159951781243, 1.63837790202744, 0.677322904056793, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.498423211983762, 0.756264624117018, 0.774967073486325, 
    0.582053879109414, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.716216315473594, 
    0.82446557105626, 1.02705518699221, 1.14114030836987, 1.31400486003779, 
    1.35293034237613, 1.36885475574555, 1.31762245354609, 1.22665008408212, 
    1.36823656014111, 1.20976425289919, 1.17921567353639, 1.16512631013437, 
    1.13366320302059, 1.07841365853952, 1.01825567569862, 0.850272796791624, 
    0.358079787157632, 0, 0, 0, 0, 0, 0.483131781955001, 0.638154125579333, 
    0.724765889822362, 0.337071319350696, 0.979602133641506, 
    0.846213879572337, 0.805575972080873, 1.06276950773882, 1.08360046148108, 
    0.333319510241801, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.930579750591928, 0.980574193366367, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.534126778122204, 1.15009809756313, 0.646288278090265, 0, 0, 
    0.572154450869762, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  2.03124105824777, 2.04461880602183, 1.98783960221939, 1.89666811394517, 
    1.38507945249475, 0, 0, 1.45558884464481, 1.63846752608274, 
    1.58837871484419, 1.57751345736749, 0.978376863176956, 0.651323847767908, 
    0.525814459021158, 0, 0, 0.27908025977344, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.568036488102629, 0.789888380880534, 0.752541316516556, 
    0.508894582780804, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.599438620693438, 0.458683939090978, 0, 0, 
    1.21481896242804, 1.34292033650459, 1.29408075684895, 1.41674118212388, 
    1.28878154283541, 1.01745575536088, 0.768002976023747, 0, 0, 0, 
    0.867589519178588, 0.594550905235545, 0.396660585510924, 
    0.652151972858051, 0.911420606756386, 0, 0, 0, 0, 0, 0, 0.36751363832085, 
    0.583514830940808, 0, 1.45554893106408, 1.6835773276817, 
    1.60432405995495, 1.49190999598714, 1.73733731528312, 1.59534844382958, 
    1.77123662668138, 1.50832303330867, 0.249914175434333, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.69871031912757, 1.19639353806463, 
    1.2510842694705, 1.2669893756681, 1.61095136071027, 1.57363737550371, 
    0.627313886758247, 0.696313668352875, 0, 0, 0, 0, 0.805297726684301, 0, 
    0.610960273712287, 0.86273205123807, 0.646661404139109, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.601524012793816, 0.855107909237996,
  1.76362042118424, 1.74643678935859, 1.74169788157098, 1.74558620293004, 
    1.70671051207192, 1.70566140016455, 1.71448982252241, 1.73425343970374, 
    1.79920385251891, 1.82820991811737, 1.82953302877288, 1.77867305846294, 
    1.66759484261494, 1.56143543498608, 1.44002118682901, 1.34862484772633, 
    1.27637979526242, 1.2581504770967, 1.23971007748, 0.781545107155279, 
    0.619454479081969, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.454094596596224, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.437032797635578, 
    0.576455960821601, 0.678125400160953, 1.0870358256917, 1.55114427376233, 
    1.63155069462264, 1.69081900253045, 1.68035371584145, 1.64558018903434, 
    1.54087564685067, 1.39842436972687, 1.24699637962487, 1.4210173889625, 
    1.41797634364478, 1.34608512629001, 1.61299644643608, 2.14614102653915, 
    2.17961873599912, 1.90128301978873, 1.61138453270609, 1.12525419807575, 
    0.783204844796358, 0.629670424917991, 0.612644344678805, 
    0.629965115606735, 0.559180237542546, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.969957695432136, 1.27859280714175, 1.36407364161751, 1.4189657678994, 
    1.49634285077833, 1.56867256933381, 1.61610530548682, 1.56926994859397, 
    1.52916908217244, 1.47988406614261, 1.63054518499646, 1.35768412090921, 
    0.246082642554668, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.87385338953133, 1.28660526709388, 1.44035163837252, 1.63556932269774, 
    1.81654158325312, 1.97920288148344, 2.14875680680595, 1.97703325678506, 
    1.81211275677137, 1.46268118049255, 0.840768686312611, 0.544803239676759, 
    0, 1.06597595710345, 0.417519507128395, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1.56208715489799, 1.8093665332743,
  1.22054550242288, 1.1947498628364, 1.20277897548568, 1.2454035277378, 
    1.30225490153174, 1.36994345510533, 1.4294235067825, 1.46968704340934, 
    1.50945636943084, 1.55818608418113, 1.5854268079444, 1.60783968543764, 
    1.62357483468785, 1.58729851345338, 1.5193618854411, 1.44366832554879, 
    1.3589819100684, 1.30588006281391, 1.25993516760243, 1.18931368198685, 
    1.13111442999995, 1.0675094467406, 0.966689842410185, 0.881512386956931, 
    0.747441051138815, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.897654938141068, 
    0.504461267438067, 0, 0, 0, 0, 0, 0.548011390258895, 0.984158955955123, 
    1.23977638078745, 1.45594819328663, 1.61548229293869, 1.75089497419172, 
    1.86753091815003, 1.85912317796314, 1.82568146590722, 1.72256347611322, 
    1.60753379626224, 1.51093235955274, 1.41748345061165, 1.33371217320076, 
    1.24677375211961, 1.17915025531166, 1.19776471951628, 1.57559848812926, 
    1.84526644865141, 2.03815923900342, 2.14242071588739, 2.03615382888084, 
    1.79746889177187, 1.51907014072016, 1.33786366931516, 1.24520757222303, 
    1.17091080176744, 1.06545150007808, 0.744550120302705, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1.10878060110687, 1.29684133914425, 1.31937929009667, 
    1.34960816872341, 1.40428327586159, 1.45029280740469, 1.49128166022502, 
    1.46504828385525, 1.55835302475552, 1.48665900958673, 0.741427262648506, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.556184129116722, 
    1.05038917699098, 1.21026770887931, 1.33743450881058, 1.44213401473373, 
    1.56761900360351, 1.71113178843064, 1.84382445751067, 1.91079631778456, 
    1.87060900483614, 1.87897179282713, 1.87517707675835, 1.38623897405644, 
    0.588215721117407, 0.302584329253541, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.568684838026986, 0, 0.61933069823686, 1.39972442442225, 
    1.50442593058244, 1.33562458808126,
  0.537240811263733, 0.59353624645987, 0.657022124493155, 0.717814242940723, 
    0.781832112518984, 0.887559254050193, 0.992888149599606, 
    1.08398283537803, 1.17615201314103, 1.26704357892568, 1.34366452520633, 
    1.39271765861584, 1.40684441256711, 1.45058739125941, 1.45785564862866, 
    1.43130396640759, 1.35680474158768, 1.30475738160955, 1.29195418633536, 
    1.21602481702926, 1.13563782608782, 1.03250970707851, 0.900006747140851, 
    0.757466773035521, 0.608870125381678, 0.535445853549014, 
    0.439474391069128, 0.390223795900099, 0, 0, 0, 0, 0, 0, 0, 
    0.477305943961009, 0.971371926090808, 1.05448347171238, 1.0556006299815, 
    1.14916143785221, 1.33269621427838, 1.48058223847017, 1.57730251168569, 
    1.55522711333418, 1.2916876178816, 1.18192797061984, 1.2759089347588, 
    1.41689713780036, 1.40959777634976, 1.37342044113749, 1.1860866423331, 
    0.994090334112646, 0.834040167715935, 0.754285809542638, 
    0.761941446018092, 0.749629049687168, 0.728523673601625, 
    0.699772453611905, 0.741380954388073, 0.870387939603492, 
    1.00392727987836, 1.16637944313648, 1.42220740301034, 1.62294789706473, 
    1.80949274983556, 1.92007431178028, 1.93636501327636, 1.8749926228064, 
    1.77831355264225, 1.63685750822938, 1.43343691942197, 1.15450395070651, 
    0.741187958676936, 0.124702646313286, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.534074148002793, 1.14118157418539, 1.20444947075212, 1.2680323595913, 
    1.33239651130886, 1.42178905298673, 1.4614237644332, 1.48240529798749, 
    1.61337697200009, 1.35946850513832, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.214591056568182, 0, 0, 0, 0, 0, 0, 0.271587811212183, 
    0.766953046991305, 0.96656696202211, 1.05997327913198, 1.26902418436245, 
    1.4652038610865, 1.54231234577927, 1.63357861733217, 1.71483712130082, 
    1.77755813779826, 1.65797264973526, 1.1016082927873, 0.796346743389622, 
    0.765998291285014, 0.549939992441526, 0.365862952916386, 
    0.412600704840965, 0.338892203406426, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.489747976029651, 0.718127803849803, 1.11522814841706, 1.35480910132312, 
    1.21095543650678, 0.778631023759367, 0.576363447257983,
  0.609820610631325, 0.627679089741808, 0.681429722071324, 0.796154524917885, 
    0.908637924367538, 1.00226777262747, 1.00893733609615, 0.95375275805907, 
    0.969016441632925, 1.03258624915964, 1.14164976743001, 1.18336112006093, 
    1.22385241868742, 1.30021883260621, 1.31224410308236, 1.26200349088465, 
    1.25073284038885, 1.26121344310124, 1.29245356458163, 1.26548169977754, 
    1.19709648625323, 1.12007047389153, 0.934037069018341, 0.716870315604517, 
    0.701334352705873, 0.751453982542386, 0.609923025816182, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.961863818843486, 0.9214604223484, 0.926730644046553, 
    1.07609168096202, 1.22838280551923, 1.34760729310259, 1.39714663745179, 
    1.24615751201337, 1.06001249635466, 1.00709667244278, 1.00566483602987, 
    1.04051148658989, 1.03202659706959, 0.921556564281257, 0.927353092865144, 
    1.06644336601819, 1.1232741283855, 1.07044058688197, 0.882658896487016, 
    0.49394332005273, 0, 0, 0, 0, 0, 0.421296145512797, 0.887502778683533, 
    1.14133681752391, 1.33721158833481, 1.530287055493, 1.70674152819521, 
    1.75156189950896, 1.66121725011905, 1.48722596817958, 1.17080889348894, 
    0.760339325982371, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.02322572332152, 
    1.14674064577529, 1.25133292375656, 1.34541844046403, 1.43828237295176, 
    1.42017412936796, 1.50652204435427, 1.66619717463472, 0.990690549997113, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.489777970271494, 0.662684684400634, 
    0.655319495677584, 0.599663918146934, 0.600489392733989, 
    0.612203548385864, 0.503875395074426, 0, 0.168677610555348, 
    0.223421763198554, 0.529213645823894, 0.72415073815229, 
    0.861494761196925, 1.1176866868108, 1.39228952196303, 1.48023164013045, 
    1.50087190389732, 1.51843233175128, 1.45015465815734, 1.10777043106419, 
    0.889007824717179, 0.940364184992922, 0.834795435198674, 
    0.704519010429922, 0.600431161648702, 0.404592978622948, 
    0.212100857822567, 0.394105455204612, 0.378333155862696, 0, 0, 
    0.42140676742698, 0.567845088639671, 0.499606170878511, 
    0.465726740303772, 0.568184946288808, 0.721839643399851, 
    0.931453133928809, 0.753512299989355, 0, 0.123407098524054, 
    0.571356199965117,
  0.661934380216636, 0.658675091385388, 0.592330119469945, 0.644165239224228, 
    0.745718880628697, 0.826350587268179, 0.930491703737426, 
    1.00629799715391, 1.02388815147491, 0.985715132098206, 1.04990584228254, 
    1.14244814333475, 1.20648122214789, 1.21577228067989, 1.20496312508971, 
    1.1818422060662, 1.16662459237339, 1.18061622152984, 1.19139857280348, 
    1.17618644581754, 1.15748040029555, 1.10536734942297, 0.927214216577596, 
    0.776274390721057, 0.733791892575095, 0.358143666830924, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.730967096730274, 0.845036099161705, 0.84641511957036, 
    1.0510954986977, 1.17316387357879, 1.23776924284943, 1.25262433535146, 
    1.19154610327651, 1.08306060887997, 1.00830104531415, 0.99981739690826, 
    1.05796979875812, 1.10848756068422, 1.18499519044266, 1.26501378564944, 
    1.27990194616584, 1.19455765980481, 1.09884067656191, 0.909595658098978, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.647772425449136, 0.998904538035011, 
    1.24173389760351, 1.22148985461339, 0.992807990300201, 0.145000082241752, 
    0, 0, 0.119153122649546, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.01471441364957, 
    1.17563133284305, 1.34567170345007, 1.40379883057599, 1.43000044079736, 
    1.40533578742438, 1.57820874031523, 1.65301265523666, 0.856692017263285, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.405779087986114, 0.679031140588337, 
    0.830402711785158, 0.829329514397297, 0.757972311817614, 
    0.716723620365421, 0.679710969703999, 0.662186654814715, 
    0.639293039999224, 0.544710996531426, 0.482879134479637, 
    0.470467404677174, 0.584824025174505, 0.802631259480325, 
    0.851698730882001, 0.782159751836873, 0.885143921341093, 
    0.996372340987434, 1.09607129165848, 1.06509562541781, 1.05344535216178, 
    1.08378553916608, 1.18933657552695, 1.17116925698933, 1.07031220792767, 
    0.809974053790146, 0, 0, 0, 0, 0, 0, 0, 0, 0.518182892810826, 
    0.679638736061475, 0.677179224659747, 0.64525441747386, 
    0.738648798082785, 0.675170492117482, 0, 0.388366208899988, 
    0.604953783349244, 0.63440318716405,
  0.556202953078627, 0.632560605354306, 0.710648324099203, 0.582741398453335, 
    0.526525636046301, 0.644280777648557, 0.831843048704202, 
    0.885387675435747, 0.898129279603235, 0.948300213748375, 
    1.00225700182354, 1.08646769308585, 1.1751728849648, 1.22699321431288, 
    1.19764792708737, 1.18563979983122, 1.17107927771385, 1.16626302184316, 
    1.16603521079267, 1.10855756728732, 1.04611527408626, 0.970268727894282, 
    0.809154016077965, 0.601236352376873, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.605148209167171, 0.836700784866961, 0.813837429525158, 
    1.05958865100064, 1.22346961274601, 1.28478604984184, 1.26744690840783, 
    1.1746523076095, 1.00875943089115, 0.884321385904126, 0.943859023507582, 
    1.07430156615049, 1.19655640980634, 1.23532854030667, 1.19297504490851, 
    1.14020272354112, 1.02386356319359, 0.62888106647344, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.459402459578065, 0.795174172638895, 0.762846129974879, 
    0.594791672744952, 0, 0, 0.375429833212075, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.563179913977687, 1.0813924101632, 1.30531897227998, 1.45353982558798, 
    1.42807952931555, 1.3711402730029, 1.36757918003384, 1.58648914486649, 
    1.63993671068051, 0.759591525449083, 0, 0, 0, 0, 0, 0, 0, 
    0.363523183943184, 0.626504445413825, 0.815630675336887, 
    0.889957701381079, 0.917408497258031, 0.832818320628043, 
    0.757903549076695, 0.737920968777105, 0.684110555965468, 
    0.695427883359111, 0.721170331574567, 0.672148006808767, 
    0.668344313681153, 0.740555223955127, 0.883502538782567, 0, 0, 0, 
    1.00081643936579, 0.902940197576358, 0.889402397419613, 1.06527054808718, 
    1.19591475247704, 1.29412892891373, 1.15597087743811, 0.803603157805955, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.698426989214269, 0.797028146704449, 
    0.726829035424942, 0.772269786114019, 0.551393093651879, 
    0.420510391389326, 0.65642809453416, 0.800651786179542, 0.666559300657607,
  0, 0, 0.798856038988149, 0.87916408856468, 0.621338044833198, 
    0.564838856540935, 0.795873992471461, 0.782169477501185, 
    0.740322559349867, 0.87215814984807, 0.99769653086752, 1.09037003142591, 
    1.17781522954967, 1.23010644135386, 1.19923653585699, 1.15507631606468, 
    1.15155368952236, 1.13691526819275, 1.02318868353188, 0.994462661778231, 
    0.900092543084135, 0.802178438228576, 0.718500695500157, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.898324461970851, 0.935813902039072, 
    1.16189062280674, 1.2927024138988, 1.35919377932554, 1.30798687544292, 
    1.19419147191562, 1.02119321268595, 0.961268839243546, 1.02403825892998, 
    1.1299224130457, 1.16382223548892, 1.08010889808365, 1.02729661178998, 
    0.932662852078015, 0.495497754053933, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.449584181251153, 0.718513055527656, 0.783251949605989, 
    0.773480857616005, 0.661889098686264, 0, 0, 0, 0, 0, 0.478076465975015, 
    0.295453410765314, 0, 0, 0.606636373352084, 0.640506832979511, 
    0.434388085201015, 0.5621253390241, 0.76208244530525, 1.17134441397282, 
    1.40636044930254, 1.45166151532071, 1.37446621615165, 1.28401138051137, 
    1.31908414176876, 1.53104006184318, 1.58076243095371, 0.650972523613323, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.42106857638401, 0.736704635881679, 
    0.896416298312612, 0.946105961894292, 0.851823181057575, 
    0.72733763717536, 0.749482214704192, 0.770478062545783, 
    0.758574351473725, 0.752201655572259, 0.769408554235547, 
    0.795591709919002, 0.910322202321094, 0.922273019634204, 0, 0, 
    0.999445034491313, 1.1250770792291, 0.961806301189586, 0.673018648840772, 
    0.708900833705407, 1.15359678549562, 1.13892533377595, 0.907485423671501, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.583317155493272, 0.70982620674116, 
    0.790068928485625, 0.685373068403103, 0.729954853393841, 
    1.00981659629847, 0.690134788857705, 0,
  0, 0, 0, 1.08266773601988, 1.15020043820368, 0.774748973032181, 
    0.887111098217257, 0.844324169345062, 0.854616238161354, 
    0.96110938523304, 1.09469392829606, 1.17272544051149, 1.25905337866198, 
    1.25228183969988, 1.18444685471014, 1.16329939080776, 1.0987436904296, 
    1.01892155173838, 0.958643202764394, 0.756733224729466, 
    0.815205066382595, 0.819399305584576, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.688783448567357, 0.839146914780508, 0.994820429522103, 
    1.24709763127583, 1.35843743632002, 1.41552985767785, 1.40290530355325, 
    1.35359069408465, 1.2528527445356, 1.21038792420545, 1.20956293862785, 
    1.1917777613493, 1.11436655855398, 1.0722567234726, 0.87505786221631, 
    0.503825985909293, 0, 0, 0, 0, 0, 0, 0, 0, 0.416026988234988, 
    0.511542753135395, 0.470339605422617, 0.534996053463095, 
    0.797759269037802, 0.893652879811264, 0.900522571190638, 
    0.529375106101848, 0, 0, 0, 0, 0, 0, 0.715584555231635, 
    0.683314003409939, 0.616860442671525, 0.680815338414394, 
    0.734590479041259, 0.731409853740756, 0.617195194907722, 
    0.651655491939858, 0.736951556361066, 1.20512315116846, 1.42976682031329, 
    1.40513944849806, 1.32215712832253, 1.2199576581775, 1.20306138272154, 
    1.34394089244028, 1.38490064406133, 0.579648050219912, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.15403029849456, 0.674079949892518, 0.821019847296875, 
    0.829561972147615, 0.685019372320669, 0.712207266784899, 
    0.792775447592526, 0.766420936863659, 0.795936778459074, 
    0.853384373582538, 0.93226885187011, 1.05812414553786, 0.683243753618941, 
    0, 0, 0, 1.09998045414156, 1.02443999259941, 1.0700645945537, 
    1.16916535835193, 1.12433229466591, 1.18150109660216, 0.891607041343078, 
    0.322807035375841, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.58519990256415, 
    0.704810035264868, 0.812467247214275, 0.727084047032114, 
    0.907572427740325, 1.14960886153191, 0.723299776041673, 0,
  0, 0, 0, 0, 1.10377933934182, 1.15732218597776, 1.09689876150131, 
    1.05104679819906, 0.974418244865243, 1.0176172023033, 1.07963895136599, 
    1.20230417440215, 1.28667085372763, 1.27917481404916, 1.21856411249627, 
    1.10972000394786, 1.10273372468487, 0.993563728195503, 0.803015811646942, 
    0.860487163218843, 0.655200310387958, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.663444717271449, 0.84255811774214, 0.919148521500336, 
    0.873885639364376, 1.00556571844369, 1.34407816948096, 1.5120019226248, 
    1.5863448154166, 1.60433594862268, 1.54160811499489, 1.38705884955312, 
    1.34163499740931, 1.29679065702589, 1.17989151916112, 1.13737531435016, 
    0.959767965662684, 0.706648558155932, 0.6514967423953, 0.564808452137321, 
    0.570109461983138, 0.6900650886163, 0.650369164560137, 0.598108656237277, 
    0.540109613662672, 0.552195938842855, 0.661575850863141, 
    0.716427730370668, 0.74700786140722, 0.717090106037206, 
    0.699752398437212, 0.774003198392319, 0.701858928822968, 
    0.0844371420992248, 0, 0, 0, 0, 0, 0, 0.500018640757403, 
    0.751892400429716, 0.754332893719015, 0.749016153445245, 
    0.76689100064414, 0.728795896577477, 0.671819197341348, 
    0.567364000328642, 0.593429107627974, 0.723526694322294, 
    1.22831036071785, 1.3753367095321, 1.33394752418724, 1.26219228626844, 
    1.13985258239204, 1.04826321675275, 1.10633655263995, 1.14901899293072, 
    0.672886641725691, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.390249283672377, 
    0.59494430944306, 0.798261031033185, 0.781313675983757, 
    0.727248885169272, 0.811343268734989, 0.846194537503426, 
    0.917548784826097, 0.992622067833689, 1.07084834827067, 1.14181306623331, 
    1.1153989110575, 0, 0, 0, 0.776675148906408, 1.15432781709887, 
    1.07009515373762, 1.03275438331881, 1.14264597236898, 1.24877265737362, 
    1.02972871859858, 0.792457499425963, 0.597833728394104, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.649234922221727, 0.726966362810416, 0.731689381699192, 
    0.840453346854427, 1.06944460463473, 1.30699910147213, 1.02069128246362, 0,
  0.599845148968907, 0, 0, 0, 0.399276790073153, 1.32574205989475, 
    1.21695563093254, 1.21596714124327, 1.09687946309314, 1.05864403989888, 
    1.17280847736406, 1.30547985393263, 1.35298937429723, 1.2892203278178, 
    1.12085357901695, 1.0920062479753, 0.987296790865501, 0.886644850692082, 
    0.906978566222439, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.258616682927478, 
    0.515049536774102, 0.682344855315143, 0.872279926859806, 1.0193581056343, 
    1.0774774629161, 1.05359701780344, 1.02042357274867, 1.09141425635466, 
    1.42339350730882, 1.61165123641931, 1.69582807825681, 1.64392705650953, 
    1.41920890826855, 1.34264023746383, 1.35531244126988, 1.24333662698321, 
    1.18387521434578, 0.957220367506261, 0.638620418286423, 
    0.667954384037315, 0.750803943170405, 0.888815007126481, 
    0.89010078442849, 0.907758050367146, 0.859705554304005, 
    0.814065983939608, 0.801455353544824, 0.816950045964789, 
    0.784538541116845, 0.798827407407048, 0.870198522936929, 
    0.965795411326908, 0.869164451212791, 0.368505442371831, 0, 
    0.73654038054691, 0, 0, 0.409751506708269, 0, 0, 0.44218444820594, 
    0.697233753363826, 0.792138325310928, 0.759736257819094, 
    0.727133018616384, 0.67212139749151, 0.656549005182354, 
    0.664503787407202, 0.550235994050221, 0.544723566283683, 
    0.801187432641784, 1.27487027208646, 1.32547061460823, 1.27956477549727, 
    1.2248142033381, 1.10272710385746, 0.95799419064487, 0.910498211532964, 
    0.920175512534327, 0.83262383222002, 0, 0, 0, 0, 0, 0, 0, 
    0.394974113107818, 0.398020193877214, 0.330250672579192, 
    0.595391608526039, 0.688332657702768, 0.775867647680696, 
    0.808409444696147, 0.811684929003529, 0.87193946605151, 0.97500966073618, 
    1.0152684258294, 1.10309383501931, 1.13202714340376, 1.14216080631877, 
    1.13223833929956, 0, 0, 0, 1.09812879238364, 1.28640216305835, 
    1.09401347619898, 1.00046895937183, 1.19497301770375, 1.31598150621347, 
    1.17554093781735, 1.06202821825397, 1.04746327943713, 0.782854751258753, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.773682591877251, 0.808064711494451, 
    0.851307592689173, 1.11001266013457, 1.33181739218617, 1.51807436768923, 
    1.36257325839312, 1.0771632536606,
  0.79715231133863, 0, 0, 0, 0, 1.3152324567422, 1.29390814119649, 
    1.25424677275681, 1.13609449889982, 1.11659446525893, 1.25743832342211, 
    1.37077873448716, 1.38652467575268, 1.26208557598826, 1.16754089785428, 
    1.04055757336839, 1.06543357710785, 1.23290660465833, 0.545902274411093, 
    0, 0, 0, 0, 0, 0, 0, 0.348190562823743, 0.67603144325167, 
    0.898192756159517, 0.925166066544001, 0.856756847372132, 
    0.890951012532056, 1.03937205531696, 1.13274991157534, 1.20683499804674, 
    1.19620224426745, 1.18065886849807, 1.15223256014363, 1.21592210320773, 
    1.39198623348904, 1.50596523475018, 1.52811362807555, 1.35168592362007, 
    1.27665729519898, 1.32305092761024, 1.27649679949506, 1.23440059592776, 
    1.00800051812886, 0.573598635082735, 0.570626435205107, 
    0.778316898341645, 0.879963199643684, 0.964831683473441, 
    0.956955721044117, 0.93634496686311, 0.867112478228536, 
    0.798947560388362, 0.745490137393599, 0.550659845589776, 
    0.939670213398275, 1.10922954012891, 1.12852286009879, 0.942835233583684, 
    0, 0, 0, 0.674534608897601, 0.818376847625029, 0.908429904114836, 
    0.854231194733298, 0.702887868415318, 0.69237238132452, 
    0.722344845494643, 0.784259139762893, 0.779668352660505, 
    0.710636540974769, 0.677364190882844, 0.7055704584698, 0.73314097209172, 
    0.753884403872582, 0.742503746539318, 0.78738376898411, 1.02782254201451, 
    1.29557425595198, 1.29242364390206, 1.25396102188591, 1.22307349543947, 
    1.11195472628836, 0.91602845459571, 0.813306485532846, 0.796204597628515, 
    0.854433451045719, 0, 0, 0, 0, 0, 0, 0, 0.395408701961161, 
    0.675603599558803, 0.700397894311656, 0.584126878569739, 
    0.715133343544252, 0.728363428267617, 0.76715165499876, 
    0.826277104608487, 0.869442952519998, 0.97761035974677, 1.01369993050875, 
    1.0892755531233, 1.11713909139985, 1.12933341421744, 1.0839808503298, 
    0.692379035871887, 0, 0, 0, 1.47890587907762, 1.08719898965238, 
    0.844474594230263, 0.989705175679847, 1.28563720309687, 1.28882064385969, 
    1.18230381829157, 1.00705004661318, 0.654406650376423, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.566920684776061, 0.755422003863281, 0.970281389713595, 
    1.23185369861002, 1.43082552642078, 1.53229994710575, 1.44667113290827, 
    1.23183207355661,
  0.710787692849758, 0, 0, 0, 0.370976165784187, 1.27615722830915, 
    1.43517796286228, 1.34505985744309, 1.10729041798153, 1.21489210422058, 
    1.37043765932589, 1.45970604176189, 1.44785052820162, 1.34624436079231, 
    1.23126836642677, 1.28105582572852, 1.54750235468173, 1.03932775452548, 
    0, 0, 0, 0, 0, 0, 0.691741544853129, 0.782983854528866, 1.00551696470935, 
    1.02958808934808, 1.05686959782056, 0.998791717329152, 0.963132280189604, 
    1.00345021922224, 1.14609834420115, 1.19382419358882, 1.21535907880698, 
    1.21899086155748, 1.20745321086258, 1.19607680741219, 1.20676202556051, 
    1.22614722218091, 1.22191582576973, 1.22200264795326, 1.18006137894075, 
    1.28761436134251, 1.31456216119476, 1.32203703302379, 1.07398967753477, 
    0.717981965708136, 0.706177608574481, 0.879256918134871, 
    0.927091988283212, 0.940853976219296, 0.960162145766191, 
    0.821515929627328, 0.698474710697964, 0.714946050324226, 
    0.679181442960283, 0.752897170812395, 0.577543407692237, 
    1.14534197241308, 1.22443226750945, 1.07509992840502, 0, 0, 0, 0, 
    0.558231156309265, 0.72306726698442, 0.919234847066983, 1.0345514143075, 
    0.927520704448128, 0.782550610834738, 0.712207374447755, 
    0.720129170243103, 0.676273614212947, 0.634948399806513, 
    0.668608564508587, 0.751469285577752, 0.805807704888357, 
    0.843200446449335, 0.907283934332872, 1.0089527348198, 1.2058138722146, 
    1.29296249504939, 1.28333851852565, 1.28339988441819, 1.27500703382522, 
    1.12817795823009, 0.89663018806077, 0.829177182028605, 0.823955566212313, 
    0.91662231830957, 0.258250228088269, 0, 0, 0, 0, 0, 0, 0, 
    0.694692635987645, 0.797350197726058, 0.656753103194168, 
    0.886615699562698, 0.780599318825926, 0.831589857318146, 
    0.830070340030735, 0.85911963930029, 0.92051262971066, 0.975919697994135, 
    1.0527354497535, 1.10349976963882, 1.1118189078086, 1.05922069961286, 
    0.882418432205231, 0, 0, 0, 1.33014623214179, 1.27594963160969, 
    0.829313252059124, 0.470148351363704, 1.11482309081206, 1.4331908068942, 
    1.35146371172261, 1.09541120100617, 0.977573091595616, 0.586876621590415, 
    0, 0, 0, 0, 0, 0, 0.374142130453898, 0.577814323937503, 
    0.611114071236818, 0.783505578953291, 1.03008906575239, 1.24150478243112, 
    1.35705587094599, 1.39771055274045, 1.38811932391424, 1.09862843867493,
  0.768882961861186, 0, 0, 0, 1.12704486893821, 1.41631933546166, 
    1.47108527504213, 1.30067280502391, 1.12033607059631, 1.32147539709767, 
    1.42336901220196, 1.48619717274801, 1.48308057608943, 1.35947880331174, 
    1.36865307067006, 1.65440286621298, 1.34859636576192, 0, 0, 0, 0, 
    0.356322864554516, 0.671706654223169, 0.732846119609672, 
    0.778534294183854, 0.881595317161527, 1.01205051903799, 1.00158634075898, 
    0.938996879858032, 0.840032344207613, 0.928749821097888, 
    1.04048640989923, 1.16089165709615, 1.20898022073944, 1.17916935264967, 
    1.1770493443337, 1.20064688957253, 1.2051279383233, 1.17533830733588, 
    1.15341824134024, 1.1783903326049, 1.2290938730697, 1.28832034513148, 
    1.35966772151166, 1.39507984826666, 1.18635564814014, 0.876911505177225, 
    0.860283214260843, 0.942535170985998, 1.02116104713572, 
    0.924254762592484, 0.822933983272166, 0.710684478185993, 
    0.654566938245346, 0.710511086671095, 0.764554418679709, 
    0.677939942782836, 0.805676693693875, 1.15634046058701, 1.3489278907849, 
    1.14400505951986, 0.373454188874807, 0, 0, 0, 0.365961903281655, 
    0.650774279780438, 0.728840775006949, 0.880419492003335, 
    0.953738702913615, 1.0932945895655, 0.815426680179148, 0.728600661926844, 
    0.69566387437243, 0.684940879322373, 0.684865674384085, 
    0.734362074670544, 0.827689613428565, 0.905431259313763, 
    0.939969431098939, 1.04117842670788, 1.15885973170447, 1.27207221790105, 
    1.29180926287631, 1.3191569130403, 1.34365464466482, 1.30992901462336, 
    1.09168933460551, 0.930633667690941, 0.896624170282194, 
    0.903226708462331, 0.984261573062539, 0.296313707655669, 0, 0, 
    0.325756149198034, 0.320243488344739, 0, 0, 0, 0.245750316712631, 
    0.728658173530569, 0.767387932605061, 0.882203045043305, 
    0.886609116611252, 0.891574204273141, 0.899646059901192, 
    0.889458910748853, 0.912034274758237, 0.96920455295291, 1.05199528318131, 
    1.11289547002308, 1.11355624858239, 1.08996912466315, 0.479195701351515, 
    0, 0, 0, 0, 1.02294848183606, 0.833458066150193, 0.768541138263367, 
    1.17221208581329, 1.57859003090998, 1.43668212428768, 1.16869091847442, 
    0.984481612532209, 0.494765407467573, 0, 0, 0, 0, 0, 0.435179763071438, 
    0.66874649991872, 0.691098138145193, 0.620662140466286, 
    0.672211046006729, 0.87077216750139, 1.0293516470361, 1.11439085887717, 
    1.14966749842829, 1.09984734632029, 1.00567415389614,
  0, 0, 0.284315963820188, 1.14701681665654, 1.33868895248161, 
    1.40765890485539, 1.33112615868942, 1.09667739392522, 1.17874639198357, 
    1.42270174815506, 1.52226485919483, 1.54068360710456, 1.5016628716003, 
    1.38573398251534, 1.51020822612062, 1.43980678227089, 0.551479884618085, 
    0, 0, 0.616003444103694, 0.669676881153759, 0.755916881958864, 
    0.788224739664833, 0.772218662116458, 0.814320865423277, 
    0.923008375616279, 0.993941759216854, 0.97188837687658, 1.00955368516347, 
    1.00304130755365, 0.994353310403836, 1.03277806944605, 1.11138493039462, 
    1.14328025332827, 1.17777511056967, 1.18396470470384, 1.19305732699498, 
    1.19111671926127, 1.19566975266682, 1.20998871268446, 1.25563012585681, 
    1.31542697781628, 1.36920143860855, 1.42719168032744, 1.29704442958218, 
    1.06786534656003, 1.05708321955103, 1.05606525404985, 1.10891846740046, 
    0.958656570737559, 0.754825082152991, 0.714096788194342, 
    0.667264059181886, 0.721266124894825, 0.793380082305457, 
    0.726152145841635, 0.379965086521394, 0.752548505976448, 
    0.562726601150006, 0.664829546548751, 0.679621373542547, 0, 0, 0, 0, 
    0.567906100125978, 0.698983218980849, 0.752413655657435, 
    0.782862255230531, 0.852759659489558, 1.00717124231674, 
    0.944445544665851, 0.866366004260883, 0.831840614656543, 
    0.818121634958613, 0.81159696733722, 0.867076267976997, 
    0.923734052930484, 0.978868205540723, 1.01908726625626, 1.09772129299538, 
    1.18230116029834, 1.26426630785391, 1.32246811982791, 1.36984413035867, 
    1.37810424201045, 1.24777554864751, 1.10211688841286, 1.014324304229, 
    0.942028712210345, 0.946468412108634, 0.973056669348628, 0, 0, 0, 
    0.587226550748571, 0.665251292279882, 0.519814048772361, 
    0.396000358327309, 0.125078861055636, 0, 0, 0.714477832498133, 
    0.95313659067236, 0.979619473468105, 0.981243694077532, 
    0.996280438363504, 0.954777693839038, 0.943878773970028, 
    0.997729076778143, 1.0764954492803, 1.1165152127944, 1.12456632245213, 
    1.10084811920988, 0.759114279803918, 0, 0, 0, 0, 0, 0, 0.888646135966743, 
    1.23554706139528, 1.41518732896877, 1.15799127776349, 1.11281488946813, 
    1.01076650417485, 0, 0, 0, 0, 0, 0, 0, 0.444793304700916, 
    0.671992496174053, 0.672657882465636, 0.584757498312633, 
    0.778970808142191, 0.938634657894009, 1.05479159127456, 1.11617547230813, 
    1.13203921235661, 0.97864662363964,
  0, 0.417578430395718, 1.03404721994155, 1.23661838584574, 1.27240085055813, 
    1.1895354637783, 1.05093865786131, 0.875090210325934, 1.09260036164627, 
    1.38948041383128, 1.48284003224611, 1.51701394995372, 1.46634909383637, 
    1.44309411444298, 1.44728311464539, 0.797111756926709, 0, 0, 
    0.548584081764022, 0.626677647714173, 0.709466656996645, 
    0.826749967327596, 0.833806825791531, 0.77224057419022, 0.77853034528646, 
    0.885676607474367, 1.01136888316032, 1.09099375784835, 1.16294858988542, 
    1.19553294295806, 1.1526176277028, 1.13062323546396, 1.1450460472925, 
    1.17059837255554, 1.2141627657096, 1.22630380714387, 1.21819364718501, 
    1.20298693750145, 1.23625417417956, 1.28884204479739, 1.35717558826416, 
    1.42772876027517, 1.47223584379456, 1.25743014520046, 1.14781720453826, 
    1.18963040993234, 1.02316369190573, 1.04246188932522, 1.137500515314, 
    0.957318603176987, 0.856711649862275, 0.838102977143458, 
    0.816576996394508, 0.86534743507217, 0.574158462142975, 
    0.327961190557167, 0.967015536031167, 0.931996780912327, 
    0.826514329563756, 0, 0.839799868504118, 0, 0, 0.50906104557442, 
    0.715195333962191, 0.722795553337812, 0.753787428505577, 
    0.796163571205001, 0.880230450231724, 1.03555554039297, 
    0.960221878726229, 1.02121939273857, 0.942117896697966, 
    0.946253691517065, 0.939867898591617, 0.934998080301901, 
    0.978572352257022, 1.02588232706482, 1.08325067130481, 1.12167723327127, 
    1.18163947542439, 1.23762629053352, 1.30692904535669, 1.36708355883725, 
    1.37033964763611, 1.28352513531294, 1.17164373283913, 1.11360074629367, 
    1.02266591926446, 0.928815986296706, 0.933816250592503, 
    0.841515249959647, 0, 0, 0, 0.597917540042721, 0.751625193900327, 
    0.722306187854896, 0.611360382530958, 0.570225671797623, 
    0.295484500835898, 0, 0, 0.805108190747273, 1.13258264330393, 
    1.06455551497726, 1.11643631088388, 1.05436959097954, 1.04845874159726, 
    1.07935586774919, 1.12177031725735, 1.14682946905823, 1.16230482497995, 
    1.17636201766841, 1.32132709926736, 0, 0, 0, 0, 0, 0, 0, 
    0.920107807613405, 1.12562731677993, 1.25914969430615, 0.989525021852261, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.401549664012716, 0.615632336815167, 
    0.687106347151782, 0.772263839635149, 0.87761486965517, 
    0.952492297657767, 0.904972342674945, 0.669489722870075, 0,
  0.786651672703865, 0.947491780178889, 1.09342743301692, 1.0916444083799, 
    1.00139848192808, 0.968086319210347, 0.98872807799872, 0, 0, 0, 
    0.595252442125519, 1.43951937986901, 1.42365615497579, 1.42806021018336, 
    1.22115484210489, 0.438029860066621, 0, 0, 0.406564168153055, 
    0.727476203453254, 0.774708966937779, 0.85402157787703, 
    0.845259791982207, 0.823904362274051, 0.808844463518302, 
    0.886765835402586, 0.992938300390839, 1.13867897787146, 1.23675001872912, 
    1.27274896127883, 1.30919142058018, 1.30127178665076, 1.30250675306415, 
    1.29440941171938, 1.29729623369074, 1.29738974882253, 1.2999938394573, 
    1.29092396038389, 1.32412924466384, 1.3915854875912, 1.4857868030037, 
    1.47090870153051, 1.2459716946064, 1.07156638204168, 1.19551037347871, 
    1.24131955843016, 0.214519186042999, 0, 0, 0, 0.882602494341132, 
    0.990523008885391, 0.991775972303132, 0.865258462987482, 0, 
    0.808007330465359, 0.991190484494416, 1.0947882563527, 1.05929925666187, 
    0.408945602855141, 0.95481089547832, 0.610299916020556, 
    0.756412467668193, 0.896379098518187, 0.859342401171831, 
    0.901016262593373, 0.889186712161165, 0.85869773446386, 0.91463778739611, 
    0.991508409396903, 1.03566899072027, 1.02230275562108, 0.997311172580857, 
    0.991364558140051, 0.998211975206563, 1.01502990371189, 1.06015116478312, 
    1.10118729947566, 1.14390012436689, 1.17256541232475, 1.20460466685642, 
    1.22465970229927, 1.26169867549136, 1.27875235126241, 1.23993972776278, 
    1.17352190172109, 1.15686660849133, 1.12695692149725, 1.02839165529408, 
    0.933420589238639, 0.931230987604517, 0.661813929141138, 0, 0, 
    0.564165870297466, 0.814529747082454, 0.832557937877054, 
    0.812818046689064, 0.783690918981775, 0.744012812813108, 
    0.574632703430051, 0.316266503620507, 0.463193285019173, 
    0.299911619348041, 1.14343522797846, 1.14139949641476, 1.17366813466975, 
    1.15001631950606, 1.1410824460245, 1.1509451697267, 1.17841115397995, 
    1.19307034254952, 1.21549141468047, 1.2217678395649, 1.33300581248911, 0, 
    0, 0, 0, 0, 0, 0, 0.442924206423015, 1.20263994018618, 1.32197355905763, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.286720504464527, 0.38592536499992, 
    0.4726722214121, 0.504500347893059, 0.525544650518873, 0.478478351943175, 
    0.311428718529382, 0.358226524971471,
  0.882235522512224, 0.921054785474056, 0.87215660219468, 0.908435956417775, 
    0.995856348972098, 1.0574241410399, 0.995590300874523, 0, 0, 0, 0, 0, 
    1.44342655765583, 1.49307651435749, 0.959275925345844, 0.534565040944199, 
    0.490255264520785, 0.408329700876483, 0.591297061921707, 
    0.779314066258712, 0.863662015425181, 0.929865886878928, 
    0.940465408109012, 0.935420566441368, 0.924310415402232, 
    0.942217876644898, 1.00098958857767, 1.09089725706151, 1.16927438005234, 
    1.2380759189577, 1.34358827706894, 1.3992984501578, 1.42565242949739, 
    1.42274065488628, 1.431110732745, 1.44394695643037, 1.45879899411179, 
    1.47061821357173, 1.48657133126923, 1.49251106864657, 1.42458477694545, 
    1.22382489220071, 1.10401229362761, 1.1690859892253, 1.28749385604975, 
    1.22474334508345, 0, 0, 0, 0, 0, 0, 0, 0, 0.865496168274885, 
    1.11561317432721, 1.10343557628302, 1.27095079499343, 1.32506286721076, 
    0.981994826296994, 1.0294828311157, 0.797426588820485, 0.792480787277035, 
    0.921031663608387, 0.968033106389225, 0.958381480242553, 
    0.987281193855031, 0.93602781480892, 0.979390483472886, 1.03994289075091, 
    1.06261035712442, 1.07505943530221, 1.07784613495399, 1.06128322128642, 
    1.06582969388598, 1.08618632959401, 1.12520117554705, 1.14636194098497, 
    1.17596510003386, 1.19387032435011, 1.20270385641945, 1.20385742075485, 
    1.2067266544945, 1.1858493459981, 1.16383092740636, 1.16221895092062, 
    1.18114308170155, 1.12678553084661, 0.994604322648685, 0.951671013720887, 
    0.958386228385124, 0.580226311964542, 0, 0, 0.70924017288847, 
    0.921035927477501, 0.894673577261497, 0.775400515308713, 
    0.763646696532379, 0.809378258612711, 0.562376480400179, 
    0.49966790619046, 0.718393980096824, 0.698528626171272, 
    0.919895097108629, 1.28511948461381, 1.19962097607869, 1.22634929458637, 
    1.20336829867153, 1.20240513728589, 1.23942969364155, 1.26588896571507, 
    1.2713668696859, 1.23100523749993, 1.22328417786559, 0, 0, 0, 0, 0, 0, 0, 
    0.369500558835071, 0.693989930309871, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.157851523593197, 0, 0.218138652064915, 0.270458929700819, 
    0.377807761991452, 0.365555614510791, 0.416131744185162, 
    0.443413962300706, 0.499884853408543, 0.529521516088345, 
    0.585984539766913, 0.764427060051008,
  0.771753246005309, 0.914131289170451, 1.00954684960995, 1.07212128627986, 
    1.13230386287028, 1.09408525132341, 0.536108225533821, 0, 0, 0, 0, 0, 
    1.00787732215329, 1.18005293010004, 0.66259394282186, 0.737302854232302, 
    0.830706540624363, 0.78556203544962, 0.78841703843081, 0.83178588281782, 
    0.943486981075326, 0.991472029051695, 1.04894986334803, 1.04775330017285, 
    1.05628312093175, 1.04034097992886, 1.02662619728489, 1.06750172767691, 
    1.11940556283904, 1.18793368366357, 1.28142048898993, 1.35776219721102, 
    1.40525271606194, 1.43989130555111, 1.46472349507133, 1.49017485339454, 
    1.51011818659655, 1.50497739314908, 1.44136510328466, 1.34039669847001, 
    1.21013212944424, 1.12147679212242, 1.14555911746909, 1.20593167026635, 
    1.30262647522846, 1.1906595706956, 0, 0, 0, 0, 0, 0, 0, 
    0.223006534590551, 1.01521789304008, 1.06268923048427, 1.05973461589318, 
    1.26237861464221, 1.19755955043473, 0.696739417633218, 0.956617357455266, 
    0.978822943615308, 0.643014960010286, 0.635482057916827, 
    0.814613928190934, 0.871785623936944, 0.989630445042978, 1.0012605773587, 
    1.02164640696507, 1.08426552915525, 1.09279829403276, 1.1024826355941, 
    1.13812034988918, 1.15040872799657, 1.15810102855719, 1.19903041989577, 
    1.22595953808298, 1.21628378217591, 1.22561162723708, 1.25473778367294, 
    1.24501506641834, 1.23915950169402, 1.24102394853328, 1.23573729018849, 
    1.19489618425522, 1.15696595503272, 1.13118934164408, 1.06798741699648, 
    1.04761020984639, 1.03396734201566, 0.841741722690991, 0.585650702514391, 
    0.442227905017624, 0.343895639313084, 0.853829538597459, 
    0.907292481272845, 0.8862100438088, 0.74727412267492, 0.862948506626522, 
    0.816490567651538, 0.611994604129199, 0.59652641283516, 
    0.795729661133961, 0.807056482004455, 0.687865305405654, 
    1.19878899985725, 1.2553729764875, 1.28269208557628, 1.26537006506557, 
    1.26845259044293, 1.28107803031479, 1.27552042907726, 1.28369731322239, 
    1.23866219417072, 1.15575760742907, 0.404667197467371, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.335240251779841, 0.410987140586479, 
    0.435748995738256, 0.355504743839985, 0.479853802031695, 
    0.466281377822424, 0.506355119199839, 0.535698446227036, 
    0.547361519102614, 0.598221731340351, 0.624792148019148, 
    0.695664241746443, 0.667535219314709, 0.71650885955593,
  1.05079881585618, 1.09466966296289, 1.15794565485146, 1.18055968305231, 
    1.16668260625823, 0.924929939533347, 0, 0, 0, 0, 0, 0, 0, 
    0.391658057781943, 0.707527102270337, 0.78589894088437, 
    0.798322390439548, 0.832870782636713, 0.894598776033709, 
    0.933755806455069, 0.968195798676968, 1.07017473547287, 1.11209845209663, 
    1.1369050350657, 1.14735834707281, 1.1340686686083, 1.12329609457221, 
    1.1382873955862, 1.16736232910561, 1.19741567181458, 1.2474503972552, 
    1.29974440465984, 1.33225050096037, 1.3595273285538, 1.37064279945711, 
    1.37304179976508, 1.36238435817788, 1.32863248818447, 1.26511921696808, 
    1.18320256927296, 1.11359362177517, 1.09208390800935, 1.12585759195267, 
    1.18457389188484, 1.19262596995972, 0.779005286002479, 0, 0, 0, 0, 0, 0, 
    0.278495112803098, 1.07704262668136, 1.16635659462033, 1.0446909752963, 
    1.31797241992635, 1.28205981891582, 0.941314344671502, 1.02161694600386, 
    1.0706985183703, 0.905230386042507, 0.511548935426374, 0.43983409972763, 
    0.596599668081306, 0.745315717932212, 0.896127133384152, 
    0.98414358217038, 1.02127045518412, 1.08165547907281, 1.11863817571789, 
    1.09546375159145, 1.13475263503567, 1.1939949595273, 1.22846570218306, 
    1.27365509916581, 1.33490667637267, 1.32140855404692, 1.34995774933833, 
    1.37404438476818, 1.37927197585032, 1.38346081048794, 1.37402351119272, 
    1.32106216509515, 1.25222260628955, 1.16314549890798, 1.09803234248697, 
    1.08571909373251, 1.06655590322874, 0.866022092735833, 0.801770922559553, 
    0.835159865737283, 0.605715485795988, 0.712183558030207, 
    0.935996659771507, 0.900053157396223, 0.830971671806961, 
    0.742995389885778, 0.96552264408024, 0.763191678042171, 0.64131715535055, 
    0.713745998317776, 0.894206095324012, 0.744915177636932, 
    0.618314481353827, 0.937623981348994, 1.23651305011574, 1.26165828991194, 
    1.29313654953338, 1.30867839588342, 1.33486896912707, 1.32083340765051, 
    1.32048123728993, 1.27874158382686, 1.22550035346689, 0.773195008030811, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.426720378006943, 0.387418292111491, 
    0.343052961357969, 0.570896389091419, 0.58108933514407, 0.56332333864315, 
    0.558905380625333, 0.637839552476798, 0.697114628499423, 
    0.712882665212263, 0.635552936373162, 0.778374883642571, 
    0.855693421404894, 0.859070889423281, 0.852769481504805, 
    0.943283678327979, 0.929634561734707, 0.994043982334296,
  1.12168363336229, 1.18884426299644, 1.21399501902282, 1.22962166842378, 
    1.10580467308782, 0.784860621527524, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.803374888688585, 0.735736000823989, 0.768285308135815, 
    0.764700390267851, 0, 1.03498124921903, 1.02230703971793, 
    1.0413221601572, 1.09934484538623, 1.13716831762498, 1.18252423211844, 
    1.18896800330976, 1.18421860302199, 1.21353579872443, 1.23593525159116, 
    1.24349481020763, 1.28798926168911, 1.32035989466019, 1.31792036851712, 
    1.32670797646165, 1.32513682354095, 1.298534135595, 1.24695022422443, 
    1.20688741985084, 1.18032620989332, 1.14346072282207, 1.09537200251464, 
    1.08414343360578, 1.11810992098479, 1.11494136957258, 1.07553189297555, 
    0.614245659949368, 0, 0, 0, 0, 0, 0, 0.712534714700462, 1.05748776906504, 
    1.02161828797124, 1.30611275007351, 1.45142399395696, 1.33421404814019, 
    1.41878243714654, 1.38969346069011, 1.17884917434651, 0.724513933836868, 
    0.528764281546019, 0.435459967017849, 0.494279833996642, 
    0.713321674341068, 0.865057785830005, 0.936110951213462, 
    0.967218542590502, 1.02006922646475, 1.09196057541274, 1.12313760794445, 
    1.15962899576838, 1.23343464814241, 1.21677008786787, 1.22138483901121, 
    1.31800700781618, 1.38181790457487, 1.40660892264796, 1.42549704639928, 
    1.40813981340914, 1.4019775629745, 1.40276895066391, 1.40361708834688, 
    1.32360186155705, 1.23933662555994, 1.12886802960502, 1.02335160330612, 
    0.869444415706055, 0.759568204318211, 0.713553528394389, 
    0.767879858666898, 0.579906931601289, 0.784756777199742, 
    0.928939496573876, 0.97237465617317, 0.938117147996656, 
    0.927144568863722, 0.870201162128658, 0.677412032860191, 
    0.635381521866366, 0.764382461483807, 0.774534088433028, 
    0.694534160316423, 0.734085044443409, 0.828814036611795, 
    1.03849070087405, 1.17995449994963, 1.27755128438455, 1.31575126344152, 
    1.29916100039181, 1.29943395731479, 1.29812218444938, 1.29551559704047, 
    1.16947066928463, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.625686201187914, 
    0.660442308244098, 0.729870006403329, 0.707517882999776, 
    0.716520105934754, 0.725380870387318, 0.757707744895189, 
    0.796369517887788, 0.872300901338535, 0.902356159363978, 
    0.945588382470773, 0.95341726938545, 1.0224824874478, 1.01976367659538, 
    1.03111624112228, 1.07191995784512, 1.11314615546228,
  1.1680599653287, 1.23162532408229, 1.27183998235886, 1.29071861465855, 
    0.822134324790031, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.783379262974569, 
    0.800030147942056, 0.832462542002385, 0, 0, 1.05725108993157, 
    1.03872094038612, 1.03920846951889, 1.13305947811711, 1.13474864082933, 
    1.14446238249699, 1.16848601098763, 1.25467047601372, 1.26626136622468, 
    1.28775129085154, 1.32048114463968, 1.33116700631182, 1.34453845286628, 
    1.32151125167312, 1.32094196606615, 1.32934091519788, 1.31180277567673, 
    1.24896592379445, 1.2085945247174, 1.20563154003461, 1.18373652680655, 
    1.15236002403173, 1.13420365929859, 1.12708741771277, 1.0961779191427, 
    1.09919918515872, 0.611298288614923, 0, 0, 0, 0, 0, 0, 1.11832192086119, 
    1.14476467392518, 1.21735779008415, 1.38968925065729, 1.44182603227744, 
    1.45568252066767, 1.51752673651209, 1.47868536896854, 0.999874139785622, 
    0.599387645843738, 0.562674233374767, 0.452206239682401, 
    0.414327373559395, 0.627821820650005, 0.801119611440427, 
    0.92226805521738, 0.923425682546902, 1.00013889332689, 1.16091799116496, 
    1.21158046727508, 1.30815445067301, 1.38430233683618, 1.36350085751171, 
    1.36922714251558, 1.42584466663187, 1.44047500112269, 1.44598832710904, 
    1.48252938943678, 1.48799871926476, 1.52517963413986, 1.53381612833181, 
    1.42688543823643, 1.32264473261318, 1.16500461241471, 0.990948702415101, 
    0.782785708790316, 0.863865812038683, 0.821952773334874, 
    0.644992029604621, 0.548433565807172, 0.677287024111795, 
    0.749094495410187, 0.823811013373043, 0.881687526761599, 
    0.879257979095307, 0.81607576276349, 0.710288685739037, 
    0.617936864911971, 0.577596358517337, 0.638268565244773, 
    0.693192150917898, 0.797228530808575, 0.833009166929217, 
    0.833359039492558, 0.928969468104703, 1.03466488754124, 1.1338790242625, 
    1.19581713691273, 1.24276215935957, 1.31313478496149, 1.29292880159466, 
    1.27289245453832, 1.01803371329947, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.650041603907795, 0.770948551643367, 0.817729763985945, 
    0.776900601706191, 0.777456018600015, 0.80757724091957, 
    0.838052001593052, 0.865887292099853, 0.906771795214722, 
    0.954204439334511, 0.999623197007066, 1.01698092101085, 1.04228634459334, 
    1.05440571512076, 1.06171382407385, 1.11307447752135, 1.1435393473429,
  1.16297560681221, 1.17649484701615, 1.19736680201167, 1.13158212103164, 
    0.660994508021366, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.809266136561494, 
    0.881992077921312, 0.896337404646336, 0, 0, 1.0656335251768, 
    0.917577421603121, 0.910636439496974, 1.05578799666388, 1.11393209972037, 
    1.13249941905287, 1.17343018158244, 1.30399644725339, 1.31754164042896, 
    1.3281935936726, 1.3840125037689, 1.37811966873776, 1.3779976501402, 
    1.3506378472487, 1.33769038908087, 1.33364930986445, 1.32222257098765, 
    1.2758853220453, 1.23028740398706, 1.21992339628748, 1.21500645717867, 
    1.19186474808556, 1.16081678596328, 1.14115099337362, 1.13417040479503, 
    1.16579393028339, 1.1781087470756, 0, 0, 0, 0, 0, 0, 0.943678519198467, 
    1.2172840010509, 1.32849839954322, 1.37032988445407, 1.4431121276233, 
    1.46178182646086, 1.55253410603313, 1.2945725141524, 0.60787893014149, 
    0.635691757713402, 0.62358259826922, 0.600885036378642, 
    0.575501091666707, 0.56071732666915, 0.929155649691017, 0.86982131967918, 
    0.957955223229645, 1.01959015582365, 1.09855943142843, 1.20243096609222, 
    1.23685842897145, 1.26655531026292, 1.24497209142395, 1.26755184416191, 
    1.30882951357737, 1.35117976105684, 1.39377397481743, 1.38293670591382, 
    1.32468229568095, 1.19073334121661, 0.98770271315902, 0.799265099880007, 
    0.787354071833196, 0.873271351826513, 0.887139470725912, 
    0.806380969787252, 0.722763774044418, 0.534256093729869, 
    0.570349054759046, 0.663057737214179, 0.719734611508057, 
    0.78490866113459, 0.831438925057773, 0.874108238167119, 
    0.867704415209221, 0.828706899199157, 0.675855771417787, 
    0.573866511125533, 0.604631960046676, 0.683830688284562, 
    0.757262758429335, 0.823600220309296, 0.854226888503117, 
    0.805637020671892, 0.862486165700676, 0.880634540795573, 
    0.929239684803492, 1.02060650224602, 1.09354911516863, 1.11813133520753, 
    1.06324380965753, 1.05262371506532, 0.786651766309034, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.791220411276268, 0.846410317721621, 
    0.844962621345979, 0.854111784068555, 0.881338725111985, 
    0.906444380954871, 0.915285126203222, 0.929793492332309, 
    0.96719763524483, 1.02485318774547, 1.0596405790528, 1.07148476159201, 
    1.10662275968605, 1.11108203230884, 1.14140580150837, 1.1387894967313,
  1.07447784306325, 1.12515058447167, 1.08109997585446, 0.835844062884168, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.413168800912631, 0.976392137433606, 
    0.947544903406554, 0.230199581536995, 0, 0.531650996625195, 
    0.876211339300464, 0.869478849079937, 0.880394641511189, 
    0.969091928786054, 1.03536587835154, 1.16170126430416, 1.28265559295253, 
    1.28653269364889, 1.3123423975822, 1.37039029935419, 1.36458028981886, 
    1.34621158173057, 1.32330265098513, 1.30701937506768, 1.28507907846896, 
    1.26315696134058, 1.23758725776065, 1.20871351097341, 1.21595454687309, 
    1.21934774532662, 1.22566795290895, 1.21339427462352, 1.20668064235603, 
    1.20043580256159, 1.18554137416988, 1.09675004366561, 0.950735387392032, 
    0.732328726981869, 0.593745463564478, 0, 0, 0.697576238911152, 
    1.06380790995154, 1.21207616794255, 1.3202672380111, 1.36279687458094, 
    1.43219538107923, 1.46956793560917, 0.705739181964586, 0.695107117129375, 
    0.694183681180133, 0.726302043794721, 0.757033644887723, 
    0.788077085513282, 0.783974412932201, 0.687473849611269, 
    0.628307721174471, 0.73416932159226, 0.784274436425157, 
    0.751172346710197, 0.758300179206926, 0.772928635790689, 
    0.767041861940129, 0.817148587654234, 0.874109361242159, 
    0.922180399967573, 0.955398596226125, 0.97398060560764, 
    0.862096633463093, 0.698057823356086, 0.568705021787142, 
    0.617098721916179, 0.658930508926011, 0.674465673130396, 
    0.592693949402357, 0.615916117627965, 0.656465640297371, 
    0.660142309663982, 0.634045677604237, 0.657956034570745, 
    0.669134947830524, 0.714093850014309, 0.788289480981718, 
    0.838141584045943, 0.864019371594827, 0.899946252467743, 
    0.888931335232653, 0.830614565187177, 0.743033577145808, 
    0.688591386535416, 0.724651250599223, 0.772271729064041, 
    0.795007948666514, 0.82833282906957, 0.857107630018992, 
    0.864126445716998, 0.864667066164627, 0.902279857908369, 
    0.906297708395732, 0.96378551700724, 1.0142597452544, 1.03538770863103, 
    0.984399440798415, 0.953087129762603, 0.804669376033025, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.782100658554142, 0.876052911889228, 
    0.910992652204369, 0.900057514518431, 0.923258594480575, 
    0.941306950348653, 0.969959905801421, 0.989976775652194, 
    0.985211430517091, 1.01836494967597, 1.08259090843234, 1.07666138075632, 
    1.08405901940249, 1.11628000031836, 1.11417285487093, 1.09551580114449,
  1.0933910555539, 1.11503006162709, 1.03700653123041, 0.757920054974199, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.442020141311613, 1.03298795933046, 
    0.563912077526701, 0, 0, 0.901532896008858, 0.874951171463175, 
    0.874254756456557, 0.911849777875243, 1.00816630035162, 1.11302921988145, 
    1.20597034081487, 1.21866491996439, 1.24217176661916, 1.27642809716545, 
    1.29117389206178, 1.27252639983228, 1.26703943779487, 1.25836214365516, 
    1.25247556547685, 1.26232279129841, 1.26231744430472, 1.24267647090771, 
    1.22343285576703, 1.19805987077214, 1.16095134740563, 1.16808190702344, 
    1.155610720919, 1.1352697854701, 1.04816446937138, 0.948451511765802, 
    0.898465119510588, 0.836327046326267, 0.678306790171008, 0, 0, 0, 
    0.987321969078742, 1.13127408092578, 1.21281723690264, 1.17828419730922, 
    1.36552653873547, 1.48031504854247, 0.889343993496044, 0.702744271076424, 
    0.757290842082291, 0.788431039404946, 0.850748536902195, 
    0.883122515250286, 0.876518091045567, 0.788598748395817, 
    0.785637478000018, 0.726806622992958, 0.725114825872197, 
    0.737728491406643, 0.843372087566008, 0.928787399080025, 
    0.587036223809685, 0.572314109090313, 0.568440920425925, 
    0.519731378548139, 0.48267099352774, 0.55697169127832, 0.626510008727502, 
    0.674506709692327, 0.806006518832825, 0.734503005961289, 
    0.612941058118925, 0.6539909769233, 0.701475131651694, 0.737132397192988, 
    0.742566453922725, 0.7260505794855, 0.687410845087263, 0.663726683112249, 
    0.691733315787912, 0.732405612187902, 0.794919553491046, 
    0.874832318646696, 0.893047533159773, 0.881281896173638, 
    0.845288438625419, 0.782007276745376, 0.7645378483287, 0.781353663453707, 
    0.768883349166236, 0.799634935855055, 0.819267693092679, 
    0.834443416859139, 0.808736090447658, 0.918018567166086, 
    0.925907509184071, 0.911156261408962, 0.986923159397611, 
    0.96735001742026, 0.9876010643478, 0.991281661217392, 0.833879299855061, 
    0.432323500654284, 1.08833431056253, 0.232015041556273, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.435375390116051, 0.920512115631921, 
    0.934342441596028, 0.956796785876242, 0.978565594939544, 
    0.998975714680503, 1.01388157008184, 1.00962790205607, 1.01317693527591, 
    1.03009783389124, 1.07776180922061, 1.0756379523993, 1.05302392501835, 
    1.05709097906212, 1.03945831726203, 1.05947296290114,
  1.1450640767135, 1.16618289652137, 1.10209054080534, 0.754010488966642, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.06620679363781, 0.897982191629913, 
    0.961866894344418, 0, 0.905029198176578, 0.840275146294356, 
    0.859819124268293, 0.919148198584054, 1.01039145015839, 1.10372532790188, 
    1.17680336335016, 1.18503564308172, 1.19121595917219, 1.19791255922164, 
    1.18540328051572, 1.18967831122085, 1.2194378994464, 1.24513842467033, 
    1.24721150616759, 1.23686855382666, 1.23026085476522, 1.25120058308322, 
    1.21577580416192, 1.18206833426039, 1.11860438237384, 1.07429159913583, 
    1.01770710300364, 0.955707545908466, 0.921028501680377, 
    0.932522535611358, 0.926764931818794, 0.850421515803206, 
    0.744442916799809, 0.506141595801005, 0, 0.660232578047331, 
    1.17448526365427, 1.18497805810817, 0.98213738532133, 0.694577820477147, 
    0.897957465235141, 1.48985707001679, 0.833602776440657, 
    0.838550537962211, 0.839816484266125, 0.871558095086972, 
    0.928526103230193, 0.913979686234128, 0.806351834282733, 
    0.770631961675005, 0.774676346503659, 0.774397688076661, 
    0.788054553973564, 0.856403926691818, 0.878809729613235, 
    0.774935990730578, 0.685616330736615, 0.657831335722963, 
    0.579110401824665, 0.476715584222675, 0.522872410536443, 
    0.548703444090091, 0.566320093746022, 0.593477632730618, 
    0.637271776477712, 0.670588750098297, 0.714624200788907, 
    0.738119594961697, 0.7470820171718, 0.75536951364619, 0.75484528358198, 
    0.717972341299061, 0.682587257794408, 0.713624609448641, 
    0.749145469274454, 0.772809183714704, 0.804580672065611, 
    0.840828397226507, 0.832212627678074, 0.824421154705844, 
    0.792870657792695, 0.780525076389619, 0.823705598855549, 
    0.834901011623734, 0.851813776377569, 0.839084404925403, 
    0.872408872805178, 0.873372718934915, 0.881807538881013, 
    0.915162909553661, 0.919935232352477, 0.999772564515238, 
    1.00827272946973, 1.01430793503642, 0.891560850590651, 0.888881862764104, 
    0.727314035564355, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.416058220105727, 0.927231777797199, 0.938640202425952, 
    0.989357272759895, 1.02126685685207, 1.02241778319364, 1.01934117080893, 
    1.0503657927703, 1.09088452503616, 1.04826777936984, 1.07540709374043, 
    1.07400660351825, 1.05034367269179, 1.08243113152447, 1.06985674728069, 
    1.06440876793609,
  1.20400619412966, 1.19257793948231, 1.09167209929673, 0.889904042885556, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.07133763741875, 0.957224602256657, 
    0.997680863111355, 0.645826248019151, 0.853675391022184, 
    0.812066735142978, 0.848983421973269, 0.904466219560585, 
    0.996989554915664, 1.07539201709296, 1.10951308352653, 1.14138790267398, 
    1.14923161848979, 1.15893110711968, 1.14472498419593, 1.14102786329623, 
    1.16794202046307, 1.15859893714646, 1.16163935482201, 1.16011295271148, 
    1.12870085481297, 1.10128206385384, 1.06797516611992, 1.00454625269217, 
    0.944932399399757, 0.918796977364619, 0.902415649133672, 
    0.890592512414077, 0.896024947793222, 0.88364733849414, 
    0.930584248722065, 0.875360063222761, 0.819232197744003, 
    0.736449204533553, 0.694987664470136, 0.799583375195359, 
    1.23501818454655, 1.23962415086575, 1.18219531591719, 0.867767241258438, 
    0.997711353420399, 1.41119689308816, 0.859780956705951, 
    0.904800968173097, 0.927277903589886, 0.950390388074791, 
    0.959483868277461, 0.926297470912672, 0.826994715279269, 
    0.843831043880512, 0.815818932912034, 0.889326519697322, 
    0.891698769539203, 0.870669353518588, 0.781234080719323, 
    0.723190406794213, 0.70430142847086, 0.611092662967507, 
    0.570343820434344, 0.576246985205769, 0.614267988412004, 
    0.620663882510278, 0.653625703699802, 0.667921514710029, 
    0.68908350250118, 0.718264574856368, 0.746456836885385, 
    0.749745769458259, 0.747001175010553, 0.76356722301124, 
    0.754943154051563, 0.724148022897137, 0.730551811201782, 
    0.758306142676532, 0.775668051661666, 0.820312193986562, 
    0.827539451951007, 0.8340225323108, 0.804914802227289, 0.814508976972545, 
    0.834256245808011, 0.8432304994073, 0.865269157871563, 0.899875239194207, 
    0.856591592225306, 0.860147104102907, 0.878615683773866, 
    0.894093161074428, 0.89486896341692, 0.906664328826713, 
    0.926886592477158, 1.00523397824897, 0.939256199996258, 
    0.909760052857703, 0.844971005421391, 0.782165935088951, 
    0.896767401017891, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.927593205752864, 0.954907481657712, 0.997927773726382, 
    1.01069005140709, 1.0232728531925, 1.03237248063775, 1.06678508294511, 
    1.09031387372735, 1.09933211628545, 1.14580766945781, 1.1430522957211, 
    1.12650195046641, 1.1017120147902, 1.12836986390527, 1.13326768071815,
  1.09248162106829, 1.08059576552481, 1.02647831842823, 0.923643082928806, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.05338818629476, 0.999410428518864, 
    0.932583882601561, 0.928862422827389, 0.811072019034716, 
    0.800792734874814, 0.842641482303982, 0.911607822158768, 
    0.993486915572752, 1.02343396942664, 1.03941791953272, 1.08830380712454, 
    1.10598732158606, 1.11514338200016, 1.0727675364473, 1.05111644593133, 
    1.0275144751177, 1.06625250613889, 1.10254845524063, 1.06675661589956, 
    1.00826171663108, 0.958216189966809, 0.8942725076022, 0.85130375251388, 
    0.869551823181729, 0.884260840345904, 0.912563836616197, 
    0.933934766416685, 0.924498482145256, 0.918337060424383, 
    0.936916659542386, 0.882300034990164, 0.893481862322523, 
    0.924718751155224, 0.908062216836188, 0.910540042352883, 
    1.10804030573188, 1.07711787720294, 0.972333448600769, 0.922814903536757, 
    1.08919013273679, 1.07823838052731, 0.882344510117889, 0.894464035063421, 
    1.03148359390201, 0.965359031134274, 0.979219076419121, 
    0.934166729255344, 0.865987702077992, 0.862671481747123, 
    0.828984561948929, 0.857817908353114, 0.825945432161666, 
    0.769168095768875, 0.740829355313012, 0.714642541363092, 
    0.605595867741812, 0.610646003576427, 0.663964184923684, 
    0.67627127155153, 0.666976713049929, 0.652736034778387, 
    0.661204130669948, 0.663561123348352, 0.694488797417045, 
    0.747426018337102, 0.758431157283259, 0.764323591657977, 
    0.763250173407635, 0.76090197681089, 0.744981697605984, 
    0.737193768673164, 0.749651547821219, 0.790725085757682, 
    0.782528200529825, 0.796143164391805, 0.802491307292044, 
    0.830246476114313, 0.842250710892578, 0.87422790689474, 
    0.898489842439731, 0.873485340400002, 0.868222036589315, 
    0.868331433280723, 0.852087099246675, 0.85708088192754, 
    0.877816053560673, 0.891478787436762, 0.887264729580402, 
    0.894410525783683, 0.904448109389959, 0.955318163125776, 
    0.920594816860234, 0.930672450719688, 0.748115263877776, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.613692977700417, 
    0.944972352285483, 0.995963122150908, 0.999303753726738, 
    1.04401990512108, 1.06427213345993, 1.08617540095807, 1.10802384151655, 
    1.11595670113105, 1.16911596277276, 1.19084319003331, 1.16192748685291, 
    1.12346460431341, 1.14732233634083, 1.13322112138996,
  1.08043329200176, 0.999565928235428, 0.879523055539488, 0.764991240269003, 
    0.59939047261182, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.02504222095974, 
    0.994670808067972, 0.931288074892839, 0.867174799706914, 
    0.810754371845536, 0.817929756401601, 0.824060356536169, 
    0.89550212077506, 0.960998376471638, 1.00754688936653, 1.01882552493964, 
    1.04537816805044, 1.06703547023419, 1.06646028809487, 1.02130506174627, 
    1.00763881753269, 0.991445843719129, 1.00786696131059, 1.03534618719657, 
    1.02434046584504, 0.945948917589527, 0.885438236739546, 
    0.837997366130431, 0.82605223205133, 0.869539553258234, 0.90104522090752, 
    0.981576682167979, 1.00216883402331, 0.957124342688182, 
    0.941720152850595, 0.896201327494187, 0.941609330507411, 
    0.910559222508976, 0.957703528077123, 0.993334005522098, 
    0.958377502651066, 0.981175289567451, 0.954858734971432, 
    0.894880109240051, 0.839424418511623, 1.4178094700632, 1.07729222729271, 
    1.12700669956594, 1.17746020365717, 1.00945099468593, 1.02168684083557, 
    0.971295945405281, 0.836004755463219, 0.773591415307386, 
    0.770721016360344, 0.756077053633404, 0.744498051717332, 
    0.735634743627805, 0.711992756672752, 0.63856204661519, 
    0.570128094065794, 0.635787834183117, 0.717278873917261, 
    0.688616560685929, 0.641923465554961, 0.631235456353154, 
    0.649434604041192, 0.665798802481473, 0.700634112549496, 
    0.755135834532061, 0.777107225429695, 0.776119906529187, 
    0.775827034205368, 0.765504556839035, 0.758849827658425, 
    0.750990090276502, 0.76033582918661, 0.776945198889876, 
    0.795741910694512, 0.792159102167437, 0.816322303099159, 
    0.81664081291799, 0.810986043216335, 0.816521293576932, 
    0.872735766743151, 0.924347883491836, 0.906161843009348, 
    0.87003027248074, 0.882852815841872, 0.869905473035692, 
    0.839552491312233, 0.855391549566601, 0.852749549743932, 
    0.821910558496152, 0.836406711024852, 0.920260395552836, 
    0.931141429980691, 0.848136663406236, 0.806151780027976, 
    0.455939910149498, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.918896503511648, 0.963931888863691, 0.992558926877633, 
    1.01305959449932, 1.06037119702952, 1.08415319766468, 1.10015961314828, 
    1.12671145413016, 1.14033525852801, 1.14488890931907, 1.09949785086146, 
    1.08838328882779, 1.06040500270465, 1.12287953982618,
  0.967727154590201, 0.958017922590135, 0.899120473826741, 0.796120300971582, 
    0.636421929999063, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.0173707531876, 
    1.00411060534568, 0.96405738765483, 0.929269841659453, 0.889046344391546, 
    0.850224786755512, 0.80482611031096, 0.864908460467946, 
    0.928091835863439, 0.996187267280057, 1.04924830963206, 1.08328660017084, 
    1.10287589140426, 1.08856270298692, 1.06551033393915, 1.02549377735023, 
    1.04001380040074, 1.01530772114569, 1.00834648596428, 0.978612508336083, 
    0.930253995833217, 0.878122559981952, 0.852741572144151, 
    0.845092190543985, 0.853528324280981, 0.779421129056579, 0, 0, 
    0.517442369243551, 0.775630645675976, 0.97689237735321, 
    0.969026204349398, 0.930789777513533, 0.978837969338722, 
    0.99252558701443, 0.920110228884078, 1.00699172837324, 0.830816824316816, 
    0.846620142440927, 0.505018400320175, 0.709929708592391, 
    0.799245676254491, 1.59341606261282, 1.20892286683611, 1.02524479459838, 
    0.94680350344665, 0.847645185415552, 0.647712110545798, 
    0.600317122662474, 0.566505211979887, 0.580373920053211, 
    0.615703470235972, 0.597635915296145, 0.571042428248597, 
    0.597638420399673, 0.699803729493266, 0.737904430724284, 
    0.678177821998436, 0.640426202616229, 0.629190325237751, 
    0.667088043432967, 0.70127427120337, 0.720469797311225, 
    0.741639068286655, 0.757318210261534, 0.760772389149533, 
    0.762015054160594, 0.757900712043746, 0.747377587871832, 
    0.758587456472334, 0.755813980387443, 0.769307713124779, 
    0.78249793465785, 0.79925480909963, 0.812467983443696, 0.815735405721024, 
    0.806909469224472, 0.774701138747566, 0.792090864249987, 
    0.80337986057411, 0.835389827395866, 0.828685743465386, 
    0.829753135339557, 0.850323439563841, 0.859960454473327, 
    0.882618230870701, 0.822636035445237, 0.763335143059194, 0.8338665827031, 
    0.859134631305668, 0.84730799749694, 0.799106538566652, 
    0.723997321529972, 0.704490579542035, 0.515042944640038, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.888619095364, 
    0.946153004774006, 0.956430007543801, 0.965681950966855, 
    0.969810253316856, 0.984680905866256, 1.03950729745258, 1.04194759048608, 
    1.0154824755761, 1.05697260349312, 1.05611088111289, 1.01037561646898, 
    1.02161788796319, 1.04722462645177,
  0.867313682927354, 0.833705611635863, 0.800313854594844, 0.735907942951332, 
    0.573262411294192, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.014749480184, 
    1.01050494215409, 0.995357013698765, 0.986675450142493, 
    0.947129802145806, 0.903093632894761, 0.834710609422448, 
    0.851784714844517, 0.899115330729883, 0.962939062642835, 
    1.05314830655819, 1.09418495564871, 1.10938722755703, 1.09720006162782, 
    1.0811370472667, 1.04172694166286, 1.04350928418212, 1.01972045097771, 
    0.966502142231431, 0.935171538112667, 0.910174983722475, 
    0.887480916813081, 0.860398417146775, 0.836358300724568, 
    0.893430324775985, 0, 0.221317720549022, 0.892182130547847, 
    0.907862644192297, 0.891681264986338, 0.934984739173713, 
    0.831583435995941, 0.90667581866982, 1.03686519275877, 0.9103555905205, 
    0.867078117137255, 0.850010102659789, 0.989967905149124, 
    1.15376925794529, 0.83483789339988, 0.778614208997522, 1.16679186413352, 
    1.06753007452589, 0.990475620266186, 1.06002851480153, 0.745798088701659, 
    0.640104096138816, 0.603140172063082, 0.646479593987985, 
    0.622840968438569, 0.619277512237756, 0.641036572116026, 
    0.665379637745699, 0.694426852674956, 0.70594084149235, 0.70176362315229, 
    0.697115862943025, 0.674474160425324, 0.673266518104258, 
    0.694670947773995, 0.718271292412701, 0.720624302192304, 
    0.72760771363087, 0.741763472307327, 0.745938804970965, 
    0.743802921439996, 0.740047194312144, 0.757731971191724, 
    0.754491152216012, 0.776816562107347, 0.783296285890562, 
    0.791509465071763, 0.807519236585934, 0.810146993777718, 
    0.81984694709739, 0.820203388384547, 0.810425750793013, 
    0.801072474097309, 0.788478945483725, 0.773054330760904, 
    0.769700532510486, 0.777017956793879, 0.750238372528789, 
    0.77847398993632, 0.809117370018737, 0.82326144663642, 0.797839990996213, 
    0.764837841944849, 0.779677014981226, 0.73091182686636, 
    0.722503363391701, 0.656648402357319, 0.532268393575231, 
    0.595176317721477, 0.40752361701875, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.893840556010294, 0.898202062847297, 
    0.92302371151176, 0.914415300928158, 0.915901916890028, 0.92077609421088, 
    0.93455266017534, 0.96398257043729, 0.94284689742806, 0.923580489034436, 
    0.892833427016958, 0.867535924050293, 0.879044997132899, 0.893336869091718,
  0.731627625688029, 0.74256115765656, 0.735621026932167, 0.757717304144847, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.998560266610332, 1.0261941342995, 
    1.0023101540105, 1.00572858725641, 1.00230384786101, 0.940361788994217, 
    0.877177218372792, 0.908238488865075, 0.917361738097743, 
    0.953852612612547, 1.01788746904367, 1.01826552572731, 0.96621345194174, 
    0.975114328842057, 1.0286040056918, 0.990637556012358, 0.920977015899151, 
    0.873304073443878, 0.863741066950852, 0.86054428024124, 
    0.857747895124649, 0.850580024839486, 0.864466182215223, 
    0.865493187190038, 0.756947295611925, 0, 0, 0.864339472567798, 
    0.575888089268586, 0.291797197811376, 0.928296875798455, 
    0.939925344641087, 0.848353435557921, 0.949960015541119, 
    0.978496570649783, 1.04947234839762, 0.920827584241604, 1.23611764257774, 
    0.607464814476138, 0.748722908798968, 1.19811787106976, 
    0.989255092804737, 0.73154429953823, 0.758291004215747, 
    0.782926430506543, 0.723364022419936, 0.665737127142743, 
    0.680199706833105, 0.68576445227996, 0.656807493627247, 
    0.659590403497845, 0.684304083708877, 0.678642807144962, 
    0.694438589538636, 0.709657074003222, 0.722692155375049, 
    0.733501554146487, 0.717482985543773, 0.712521665886684, 
    0.720612568304769, 0.732009259007574, 0.734326997916192, 
    0.733333790561912, 0.756058033860673, 0.753370654336963, 
    0.747726626706738, 0.760008674554076, 0.793073091946468, 
    0.795312963295127, 0.807185721992057, 0.808460578310444, 
    0.816641012075731, 0.821537981674769, 0.809203219762753, 
    0.820437894035514, 0.801910109451096, 0.79193445861708, 
    0.786854515150106, 0.781143163062225, 0.768721829803391, 
    0.759074683638849, 0.747392650401389, 0.72142468661406, 0.73597309518884, 
    0.740177498139333, 0.73168628695205, 0.718959813002901, 
    0.698889203874522, 0.676886262661722, 0.660435275217995, 
    0.590227984319618, 0.553895070906417, 0.539114967797599, 
    0.517784205364194, 0.655040835224112, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.423009642207568, 0.883763845067047, 0.877517163884677, 
    0.846926488312776, 0.854781936539617, 0.842632571195243, 
    0.824009524750175, 0.802601814630928, 0.763481169191775, 
    0.770149833508004, 0.774852728125931, 0.723776301426377, 
    0.677912749314136, 0.664585372604094, 0.691050727368451, 0.679230396685102,
  0.699317390011081, 0.74067857625843, 0.778803854699118, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.983180546501021, 1.00397114816628, 
    1.00990948751573, 1.02577693683343, 0.971914870518322, 0.944048210803259, 
    0.947189195743519, 0.944181135509748, 0.941913730282814, 
    0.96710197069931, 0.98319150625573, 1.01026201717658, 1.02671354305969, 
    0.934242476947747, 0.806313971311271, 0.738991590227538, 
    0.725073453534084, 0.733806129441323, 0.737683077495814, 
    0.771845377042719, 0.807897827337574, 0.840468616505043, 
    0.895043889995397, 0, 0, 0.86284421238235, 0.791489803180931, 0, 0, 
    0.867926319467572, 1.03316202814691, 1.08683180673866, 1.07729085848222, 
    0.965557500377051, 0.914152038412426, 0.828296114647865, 
    0.83219538902202, 0.690737747169142, 0.670435922867839, 
    0.636391373380017, 0.701711806921733, 0.732889329798377, 
    0.750738547555976, 0.744947894397916, 0.714986182330286, 
    0.723111167975732, 0.740694289289531, 0.731402494141181, 
    0.71412572752123, 0.711929098657857, 0.729318957338656, 
    0.731628178066487, 0.73378485532847, 0.720640245067953, 
    0.716930728091073, 0.744536940180809, 0.74454654996625, 
    0.735522086737566, 0.743425628275491, 0.761531271443327, 
    0.760137805987092, 0.767509045906797, 0.794363803853044, 
    0.771162690961861, 0.757156667641432, 0.770415910252982, 
    0.786067496446617, 0.797998064301949, 0.804584211598189, 
    0.803421459931082, 0.803840478300906, 0.793819907330726, 
    0.768065771235053, 0.755738668602238, 0.749112674126707, 
    0.741769319863555, 0.735427768040352, 0.749840778540597, 
    0.73955001327369, 0.712850920022309, 0.686419430726398, 
    0.660928072853604, 0.663020693713587, 0.659614455577578, 
    0.635019123324922, 0.611193075423936, 0.577158355556767, 
    0.553460109719458, 0.559000957052754, 0.500093236888575, 
    0.49952801169655, 0.588007318614035, 0.633145839042865, 
    0.810266284669025, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.73813147640742, 0.844096492431349, 0.840465155836054, 
    0.893634031766752, 0.857656478092064, 0.851249882540619, 
    0.813535186151004, 0.8089414092036, 0.776961552993683, 0.760646842090993, 
    0.679200526921408, 0.623028700635467, 0.652911433775154, 
    0.605426162055172, 0.586324438721446, 0.613129588055017, 
    0.675962205424701, 0.731474191322569,
  0.807217581249958, 0.785188334152542, 0.791281609018404, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.963445811743534, 0.989561171187236, 
    1.0007285939164, 0.956674217896481, 0.965148985305443, 0.989064075809255, 
    0.962759812770619, 0.931688935371436, 0.888029130235078, 
    0.906761053347902, 0.977239891346831, 0.962782508732051, 
    0.74132553185375, 0.669683403675761, 0.634792603271105, 
    0.645260829402139, 0.67814835422419, 0.71977594640976, 0.733046084499533, 
    0.764718638138537, 0.855105482083702, 0.347781180781638, 0, 
    0.791587389302364, 0.933887627971184, 0.679887627196718, 0, 0, 
    0.874488200537249, 1.11469360991086, 1.02079382450476, 1.07762662836972, 
    1.03330743168382, 0.825233853364547, 0.895174239937438, 
    0.786085845816861, 0.68018930279953, 0.662424300367827, 
    0.694342602061094, 0.717104505402735, 0.726715052427519, 
    0.739150890128999, 0.74332398222517, 0.737017094216554, 
    0.746677753418606, 0.751941466785985, 0.726049498549336, 
    0.719103517269187, 0.725752347459537, 0.744217194536087, 
    0.748914872954583, 0.728733456606089, 0.706674209598313, 
    0.696276629782307, 0.745183958770502, 0.771854457315378, 
    0.777025965974019, 0.801500733545223, 0.792432959638907, 
    0.785926317186943, 0.797110383539104, 0.816843885931006, 
    0.791908866972888, 0.779589930572204, 0.781321176182969, 
    0.789900127463939, 0.80354628882654, 0.799322299234184, 
    0.817157393389799, 0.827597576074193, 0.793394541331932, 
    0.773272782464657, 0.781651054943832, 0.791673988729326, 
    0.775638574602109, 0.76529428562843, 0.781626912611228, 0.77579847969198, 
    0.778135003996827, 0.772379246795072, 0.759077888629238, 
    0.763410201782116, 0.7507111838637, 0.743443114904733, 0.721151714833153, 
    0.713975131706369, 0.685787154669918, 0.683586692802018, 
    0.678902516991994, 0.696271483715382, 0.719817461275523, 
    0.75332340676454, 0.865752549900783, 0.830869579836757, 0.42577709345157, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.83546066306869, 0.801034096368676, 
    0.846016890576355, 0.873431724279466, 0.878980054799898, 
    0.885021508796447, 0.872433864624478, 0.887902601172935, 
    0.87286847177521, 0.883632572632495, 0.851696179989544, 
    0.839747037685713, 0.799895806058517, 0.770648908424165, 
    0.726295303589764, 0.726949421232556, 0.75060499446934, 
    0.821357318362417, 0.885140003882159, 0.878369301918897,
  0.80485820998, 0.808882264552425, 0.76481639860625, 0.700527430942809, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.277165605931447, 
    0.924984672444747, 0.939515036575807, 0.943648639771952, 
    0.977774374031942, 0.983686331058887, 0.987645864460608, 
    0.945639222389454, 0.864450573645423, 0.835309494622665, 
    0.867979668152369, 0.839784030214951, 0.697376618907492, 
    0.627291143180068, 0.636122156564019, 0.678975455683886, 
    0.726505976087454, 0.752173140874028, 0.785392825330049, 
    0.803387074733116, 0.906115130513306, 0, 0.574257314124508, 
    0.69324146678804, 0.91412209263728, 0.97825831519947, 1.04593395211657, 
    0.652256780934299, 0.668946551824437, 1.14342380650752, 1.04974910783035, 
    0.97542808121962, 0.944829862224955, 0.963305003527453, 
    0.860554761084433, 0.768980163625647, 0.678047383991845, 
    0.652363280116815, 0.695645052073909, 0.731041933202817, 
    0.747397669329649, 0.733173889527864, 0.72584547703406, 
    0.718258358450318, 0.731776152548751, 0.734797238447401, 
    0.70970587502408, 0.694114208961974, 0.717301462755339, 0.73369184719218, 
    0.737330319148205, 0.706180929576829, 0.659851145011953, 
    0.601092701741827, 0.684364060895369, 0.770713403519754, 
    0.821354090567105, 0.826606548175916, 0.799317292137618, 
    0.787055829164157, 0.804071879794166, 0.827769404448949, 
    0.801087554981322, 0.778885026235142, 0.785682648902766, 
    0.79772233852546, 0.815491773580885, 0.785601187768332, 
    0.803319194440564, 0.844189663518667, 0.830662259092252, 
    0.840777706323684, 0.852022474267789, 0.875887513622419, 
    0.884677358437009, 0.866131047370574, 0.84914806095155, 
    0.832975639175753, 0.862854995630216, 0.879722030051509, 
    0.864092679078293, 0.875203495214004, 0.878221243189278, 
    0.870465901354224, 0.858599583435052, 0.852495966522256, 
    0.812691007137976, 0.805798588293091, 0.829370562172881, 
    0.831910848185243, 0.81198401832519, 0.786035940906474, 
    0.811788061908834, 0.687074750589659, 0.692078580445794, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.805662496096376, 0.794671810367734, 0.8291516513144, 
    0.855652855980272, 0.855758770625929, 0.8782886942774, 0.88959602014795, 
    0.899946501836566, 0.920121195550751, 0.972449250547943, 
    0.975046572732024, 0.984852501010482, 0.963482835559447, 
    0.940526311782288, 0.919340474863018, 0.932841627989533, 
    0.949195672021692, 0.93177581415206, 0.947388167408495, 0.902520031616202,
  0.627189584768978, 0.745925622597947, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.600864602959656, 0.881983862370416, 0.961956936488129, 
    1.05100496226806, 1.0512944944129, 0.944404059805739, 0.938085388369358, 
    0.896223025034908, 0.845606813605845, 0.79731343320768, 0.75910773700709, 
    0.69012761395022, 0.636767481404927, 0.648446328859344, 
    0.721293779658921, 0.788177141560916, 0.799923176306327, 
    0.817047148626796, 0.852749155816569, 0.733464213461508, 
    0.962233030116627, 0.598325266970243, 0.890056070718765, 
    0.830440547597472, 0.862459204866557, 0.923971700823115, 
    0.950675858512652, 0.520201350404648, 1.01011360330533, 0.9333760345924, 
    0.922963599806551, 0.935829253051638, 0.999731541704338, 
    0.908407601826932, 0.829987241138856, 0.755102384790155, 
    0.723701717867842, 0.689004682272765, 0.682904764791812, 
    0.685343771365358, 0.688956845958683, 0.697054717199869, 
    0.685858062050579, 0.694174476303153, 0.705510742994556, 
    0.663231922491406, 0.652179803926394, 0.676394463107273, 
    0.697419550588996, 0.712130886107122, 0.662149417359427, 
    0.595898914425681, 0.527848105498842, 0.581382443712338, 
    0.638019195918472, 0.672005754661952, 0.675183766349061, 
    0.640765682512392, 0.60937614705037, 0.621944849598283, 
    0.679874384697956, 0.723951345119967, 0.705856859542584, 
    0.716145542404568, 0.761713307418208, 0.780042005818608, 
    0.729578094853559, 0.727929981068242, 0.756978091593789, 
    0.770508643015732, 0.783533336884952, 0.765425961123041, 
    0.773623149721182, 0.814808838371162, 0.831883640084554, 
    0.811860247136376, 0.785598848995592, 0.814694405720538, 
    0.836658687684705, 0.834593250718548, 0.84424907753339, 0.86614043368002, 
    0.852870092467595, 0.823737803818396, 0.806373278193846, 
    0.780549635232982, 0.758104403405566, 0.74231300234229, 0.71955047799778, 
    0.677938474910008, 0.623363593542954, 0.513964926898093, 
    0.33915244347183, 0.655711915694447, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.713881445125121, 0.717884836198947, 0.733471252508904, 
    0.788932537872664, 0.788408470481269, 0.779706283778994, 
    0.795122416737227, 0.801146346784765, 0.784316916669357, 
    0.792638239482685, 0.852648675748185, 0.889515569960657, 
    0.906976511195017, 0.912177339410361, 0.929706352276647, 
    0.940587861793805, 0.925543624009187, 0.290935992971554, 
    0.253043153242649, 0.400991598532842, 0.392127373768181,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.630231673716345, 
    0.738023841354857, 0.896374347298054, 1.07449630962366, 1.08668412224682, 
    0.966713415132845, 0.866948218540841, 0.849906481347077, 
    0.841066672975489, 0.809993015720385, 0.758121987188796, 
    0.683728990642794, 0.628486688889545, 0, 0.940318749386394, 
    0.844761728437625, 0.856463742513454, 0.852924382602038, 
    0.877333373214231, 0.910053949505033, 0.698391882001522, 
    0.615891914610644, 0.822616176732373, 0.756301006054745, 
    0.778802975246013, 0.741828268747557, 0.744601319144599, 
    0.721334002222013, 0.874620850617044, 0.925167311952825, 
    0.774675524078845, 0.882856681957372, 1.0747571413652, 0.943326659556202, 
    0.859482020748149, 0.798345040176353, 0.759285898057266, 
    0.721303285445116, 0.670399958457632, 0.661505133214002, 
    0.70117164002851, 0.638473307281736, 0.634326677299179, 
    0.646588545071745, 0.655063451549265, 0.609587808394915, 
    0.616100590775505, 0.659755843149968, 0.679457034950573, 
    0.663280515055919, 0.606577625581233, 0.543203089236638, 
    0.563289945811351, 0.548340665025203, 0.566650851093074, 
    0.588053488436914, 0.589667769640224, 0.598299146311093, 
    0.622079657754816, 0.619790813519287, 0.641887838962748, 
    0.637064463953078, 0.63422403993723, 0.6643958353389, 0.705576520105149, 
    0.723254907233194, 0.73004933676672, 0.723695170126013, 
    0.716263777698948, 0.724324661167648, 0.737259015771088, 
    0.703797518108479, 0.692207792569524, 0.717886254206008, 
    0.732609059290417, 0.715482797458506, 0.693058826298095, 
    0.712103952009136, 0.733635453702127, 0.723553325190962, 
    0.721239096903156, 0.738176839829598, 0.763800639049822, 
    0.728537930727962, 0.713406535027618, 0.715058786188523, 
    0.696223636883032, 0.649960913480281, 0.630394208697608, 
    0.607716721000264, 0.54606213293073, 0.570618193504167, 
    0.473664554856396, 0.466548799929655, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.562065380243592, 0.630281327327005, 0.671873365064219, 
    0.682626387788455, 0.677052799059499, 0.677840034035763, 
    0.661334004321657, 0.643370485335207, 0.666009639036014, 
    0.669534350428842, 0.643793433443471, 0.648228714802746, 
    0.673135608457568, 0.702525068474281, 0.740241654664882, 
    0.740480806951477, 0.773658139923959, 0.822051114469144, 
    0.485968471465814, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.279535209137033, 0, 0, 0, 0, 0, 
    0, 0.769566995806602, 1.04643262661354, 1.07662688980759, 
    1.01246313847369, 0.893526972834823, 0.82032232516771, 0.815589186762308, 
    0.826848614784614, 0.769661889416775, 0, 0, 0.868462660459915, 
    0.954498183364018, 0.865158587676053, 0.868773971612312, 
    0.855594520856961, 0.852826166154923, 0.869256017495871, 0, 
    0.971804294595544, 0.893097279284315, 0.524097729609788, 
    0.772757550587822, 0.932313295321016, 0.924008449232831, 
    0.839599951159297, 0.77914922073953, 0.96043248980475, 0.751505004385333, 
    1.10382646219009, 1.079530565772, 0.970940354332734, 0.875683681286533, 
    0.81306127142398, 0.775733974852148, 0.75991529061804, 0.702376540912518, 
    0.644248714476801, 0.667268808499598, 0.653257799337141, 
    0.622586685432686, 0.627223470176366, 0.650361864706728, 
    0.630455018802009, 0.632135533170656, 0.639669511314687, 
    0.603754262365588, 0.610854133878459, 0.544832501263895, 
    0.556333633186982, 0.557430482692901, 0.5935768818645, 0.632320281274472, 
    0.66182740337958, 0.645098545027369, 0.646594368994214, 
    0.672298533785488, 0.661206232651942, 0.683957915006798, 
    0.673369441770891, 0.69686351742761, 0.711236788506094, 
    0.709632460122895, 0.733516788661008, 0.716258098953325, 
    0.691709005425368, 0.647429916866276, 0.630437271248278, 
    0.646101036053367, 0.662077594437445, 0.651501996012639, 
    0.644333261698315, 0.641135116364246, 0.62739345841746, 
    0.634739389697144, 0.66728155761487, 0.669263919570888, 
    0.664600011660489, 0.686851162129043, 0.71541812308436, 
    0.714217760372848, 0.67238661332052, 0.650882810292784, 
    0.685727536416615, 0.685445805079689, 0.637400835552836, 0.6615364840437, 
    0.666749620239247, 0.574138595957902, 0.246577961194154, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.643543592436617, 0.636339642748043, 0.629889742562953, 
    0.63928236095723, 0.647046113399749, 0.646545261696275, 
    0.620401613034154, 0.59707634391869, 0.54817571825507, 0.532700444508883, 
    0.525209020035275, 0.511166102703858, 0.498838327869504, 
    0.506900384888303, 0.5663781322153, 0.647892689879595, 0.705551686639837, 
    0.740440928632286, 0.538471222252527, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.857931692937253, 1.05819165590058, 1.0770482731006, 1.0005248532709, 
    0.94259700408071, 0.853436130333345, 0.831323078095385, 
    0.808548026401664, 0.781413756087147, 0.536325165531595, 0, 
    0.807940252563564, 0.774249516491365, 0.755821993010763, 
    0.735303679044204, 0.702931361757759, 0.743323380200918, 
    0.829738806577529, 0, 0.989130314080642, 0, 0, 0.716842484012181, 
    1.05046496352514, 1.03628190418188, 0.915925264730777, 0.816739321371866, 
    0.826171269008353, 0, 1.10035672908898, 1.04545683455841, 
    0.945323590641065, 0.851136094138582, 0.786308897482214, 
    0.752723786385028, 0.721465875503271, 0.722459221393462, 
    0.684947295416228, 0.690064475853506, 0.685933108501976, 
    0.632963803093322, 0.591333785383797, 0.643395440752401, 
    0.679875962043748, 0.641365202086165, 0.617985490190383, 
    0.629604775187439, 0.536517080366994, 0.559277239260484, 
    0.579503693129264, 0.599528104053644, 0.638394988916605, 
    0.670413730448366, 0.660959213285518, 0.627151662682285, 
    0.615755569817797, 0.660316377698596, 0.659005616446176, 
    0.682521513653326, 0.669128588643149, 0.701004647774437, 
    0.715814908012448, 0.68496145379074, 0.686466280390228, 
    0.678983363177171, 0.686398412746767, 0.640884686893568, 
    0.573403164597877, 0.524068575193027, 0.558773764697705, 
    0.593745646755307, 0.599792894509506, 0.578660311388667, 
    0.528327977228877, 0.567856106259116, 0.627950856231978, 
    0.619675907103887, 0.615028554601209, 0.66541559765324, 0.68496050966541, 
    0.68231928340745, 0.661682286479368, 0.651307627600193, 
    0.720245692512427, 0.732501294637064, 0.660468131313694, 
    0.692880935739861, 0.820043243369228, 0.560208417325183, 0, 
    0.735772156420413, 0.693147091691836, 0.546997487038619, 0, 0, 0, 
    0.187124145866759, 0.249530995477371, 0.450604085386181, 
    0.658635945231394, 0.667850805155756, 0.660064651322601, 
    0.643879954374159, 0.630314955206094, 0.611546450923569, 
    0.591243060851966, 0.589113615171008, 0.547982290821684, 
    0.524006202064292, 0.491680102562194, 0.441926918670172, 
    0.413822382635491, 0.424079602190422, 0.459681912670675, 
    0.586743519376028, 0.68428389294378, 0.725359504261019, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.746466254261383, 0.993977230284778, 1.06103569554148, 1.012529377103, 
    0.949207108795401, 0.898216165885979, 0.882255018374878, 
    0.857666017986957, 0.867919031644751, 0, 0, 0.770042700533265, 
    0.794888795386523, 0.734485806290812, 0.670297523883256, 
    0.588193547255024, 0.653158585798455, 0.810849521965456, 0, 0, 0, 0, 
    0.64737538258708, 0.799191648341024, 0.7744983739304, 0.882486140471614, 
    0.813231685498436, 0.676199643522259, 0.864222270942286, 
    1.10902109556436, 1.04413565592485, 0.971460793257102, 0.874379338264805, 
    0.794543222141375, 0.747084749322299, 0.685520458636044, 
    0.640249250239807, 0.681210557842371, 0.692252885604586, 
    0.655597317861827, 0.566378783777619, 0.513658616102338, 
    0.513585862859113, 0.659184360412369, 0.638032148013605, 
    0.619996011553205, 0.51275989994268, 0.534460699690071, 
    0.550064036751562, 0.598048657064984, 0.608264075014949, 0.6510350508855, 
    0.662486717622765, 0.677204751695409, 0.665658376660208, 
    0.667898871809144, 0.668305232350757, 0.673374518933634, 
    0.692236848989847, 0.685583667567941, 0.702490161036991, 
    0.703219480664059, 0.657421226099033, 0.640791599352315, 
    0.679693661459136, 0.698199994052706, 0.670597403263736, 
    0.586000389466813, 0.458322493379505, 0.521024148257601, 
    0.62119262336394, 0.643488152632117, 0.649529232654213, 
    0.607630717385068, 0.612734307014849, 0.626900351163716, 
    0.591561363936235, 0.58947369826085, 0.640507043036165, 
    0.631759658309574, 0.607353540683198, 0.617524841491778, 
    0.666057322389339, 0.773944425875923, 0.799345836617252, 
    0.712281944082974, 0.717895666922344, 0.720995943070463, 0, 0, 
    0.803515500270605, 0.736643832844252, 0.704197714062362, 
    0.758900285049367, 0.761417866532183, 0.742978308097091, 
    0.687414932033304, 0.701195250324436, 0.74136470423848, 
    0.731042840497814, 0.747252131120736, 0.739250479147054, 
    0.727214059832023, 0.69884581490681, 0.665689673315839, 
    0.672358943944851, 0.707987838500949, 0.703981337349685, 
    0.682266396649261, 0.625393923873046, 0.608263338835001, 
    0.585999221712127, 0.550505027832059, 0.527124597711169, 
    0.612575040489653, 0.754116591527717, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.905972999320394, 0.928135311233687, 0.969373957212002, 
    0.988637328359328, 0.931816371872331, 0.875786864595832, 
    0.90667242406738, 0.926064001406657, 0.558991456641443, 0, 0, 
    0.836958296649482, 0.862229468382385, 0.765481009561014, 
    0.66548590162579, 0.535622314837846, 0.565964017770478, 
    0.796204912701971, 0, 0, 0, 0, 0.847444218819066, 0.659366206108913, 
    0.710389869153794, 0.808521850116841, 0.850260871523473, 0, 
    1.14279725978266, 1.13990638502013, 1.08326827431196, 0.987604777756425, 
    0.876685545283352, 0.788160776328076, 0.749590271032659, 
    0.674575951996941, 0.599880123418197, 0.639240810581498, 
    0.633454929352816, 0.53902315097971, 0.486007708601928, 0.46860334775372, 
    0.411607685447753, 0.515012029254573, 0.614290171794028, 
    0.503453022680545, 0.461246152561588, 0.475491228179727, 
    0.594932943515547, 0.604918333539881, 0.622013271707256, 
    0.630109446411164, 0.62475067690938, 0.642190469297414, 
    0.657807663461358, 0.689719123424295, 0.687836744957431, 
    0.692799763299633, 0.721863602335004, 0.75464668079732, 0.76262549292048, 
    0.782530297471993, 0.757009878959695, 0.748705598375902, 
    0.76520812934482, 0.775168635045214, 0.762414079273938, 
    0.673777860984469, 0.64899363935119, 0.701608498390732, 
    0.774706517329708, 0.782013391391671, 0.773183943368998, 
    0.744703816720561, 0.708197232880858, 0.674569941936733, 
    0.661389511323544, 0.683346623668015, 0.669765745973967, 
    0.606685745824798, 0.540648383476913, 0.554188555253409, 
    0.605272972436298, 0.940859232117272, 0.920892390617579, 
    0.859599819440245, 0.458567148654909, 0, 0.3189933362477, 0, 
    0.805414675627821, 0.718322989812719, 0.658727574459033, 
    0.69194300549391, 0.740199231619271, 0.786951800192714, 
    0.769548525506988, 0.811064197241106, 0.836699630601024, 
    0.804817920793471, 0.794010523197333, 0.78085512158972, 0.7575398996588, 
    0.732011469062899, 0.696433528360172, 0.714377961024872, 
    0.767071746960913, 0.766599936662346, 0.749105196342311, 
    0.695961389586024, 0.695036874667081, 0.678258387592105, 
    0.636004208877299, 0.579790223323418, 0.605625094425638, 
    0.672829410907932, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.491168784252801, 0.690769711542215, 0.926523240372621, 
    0.926619857887355, 0.886072772196927, 0.898440550148678, 
    0.933772368693058, 0, 0, 0, 0, 0.81486262288444, 0.676733712170518, 
    0.618759133688609, 0.564122706177423, 0.480581231953738, 
    0.366981655251751, 0, 0, 0, 0.821975126248012, 0.736498730615869, 
    0.797104983698449, 0.802508689227823, 0.829690729868261, 
    0.754556358392467, 0.597577710194524, 0.903878366592419, 
    0.818093830643376, 1.00925054217891, 0.956111067935596, 
    0.856665651888405, 0.784894085169244, 0.731681108324054, 
    0.642158647435843, 0.568883752290991, 0.577414063254852, 
    0.587086689112498, 0.4649287555069, 0.499536152745925, 0.545785091024105, 
    0.45601265208508, 0.462455526914184, 0.57001320895754, 0.497326617925501, 
    0.459942537117981, 0.508611685176706, 0.579798512720803, 
    0.618610780474016, 0.650354977631002, 0.61232535528504, 
    0.588777745500179, 0.621466977697211, 0.648756338209119, 
    0.716604643165365, 0.681296697089751, 0.669807267439192, 
    0.731443557931013, 0.791404991520159, 0.780932087140754, 
    0.790371097905697, 0.795674244089221, 0.762211923307838, 
    0.75073090453071, 0.73399699870916, 0.740802642642558, 0.721265797514754, 
    0.748916739017765, 0.811188923713266, 0.842089771057396, 
    0.783334493231568, 0.752659012883889, 0.710251369701517, 
    0.672425261373034, 0.637251428461787, 0.579625218043693, 
    0.597668801358812, 0.554705729656495, 0.50835331332317, 
    0.515383121147033, 0.638766404915675, 0.610588060419607, 
    0.765850095306566, 0.690923702950444, 0.658089399235856, 
    0.350122123388873, 0, 1.07605692238408, 0.772674358042329, 
    0.757495066019729, 0.745385109218366, 0.719296929818905, 
    0.672779763682765, 0.582898347232003, 0.812708672791267, 
    0.78536668275141, 0.899033802995986, 0.893193285979598, 
    0.869952860636721, 0.856661766518972, 0.829313811939144, 
    0.79235294020032, 0.756410853987971, 0.734139465048937, 
    0.747332029347929, 0.758297486800292, 0.785202358858571, 
    0.732325266612707, 0.689374876103249, 0.704271876383283, 
    0.70046042810784, 0.689457731409372, 0.684427791622319, 
    0.680601757791382, 0.676379847983648, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.434315754894572, 0.791388533570178, 0.881780375997132, 
    0.849328935333381, 0.813831985382564, 0.824833154945827, 0, 0, 0, 0, 0, 
    0.386185352150859, 0.531854291252616, 0.63019088593847, 
    0.611585491926011, 0, 0, 0, 0.74288610223247, 0.498088584715925, 
    0.697804628798641, 0.803223757144612, 0.841187537050232, 
    0.814795950540992, 0.749868855298364, 0.959848875977977, 
    0.965622302288573, 0.530833460097355, 0.741398539721085, 
    0.722874904295647, 0.783812152271482, 0.762904297362944, 
    0.709204213345533, 0.583688690230024, 0.550083218453035, 
    0.54877617531015, 0.528131865287952, 0.522313833229917, 0.57477161513297, 
    0.55820065126009, 0.526937414813142, 0.521681498382125, 
    0.574241583333243, 0.523373189878583, 0.547496086581504, 
    0.56061212864904, 0.61500027342952, 0.662361805935883, 0.654118461054492, 
    0.598347391152666, 0.595814947925189, 0.635776467363023, 
    0.61733180508637, 0.674194490980876, 0.646231642194454, 0.60528696201118, 
    0.674818942257099, 0.782915146689241, 1.03578144122083, 
    0.795596641410276, 0.878147649645144, 0.897260805735911, 
    0.850779751393182, 0.828478147968422, 0.821739982157516, 
    0.834395619272873, 0.822424630697042, 0.799433575802017, 
    0.782505485012729, 0.731419125672687, 0.71320030754521, 
    0.706986700755491, 0.656856493818049, 0.541475011567078, 
    0.51433984672054, 0.527464548547817, 0.493267094684078, 
    0.498092514107837, 0.558928877100727, 0.778591367495671, 
    0.373996106424285, 1.13541329610299, 0.96524611925126, 0.721280407079565, 
    0.475094208289865, 0, 0.834180396812128, 0.672061095770986, 
    0.500343410260277, 0.411560952788786, 0.388555207559803, 
    0.525996311671656, 0, 0.719997009809236, 0.746775053794502, 
    0.871516475662967, 0.855150085597537, 0.86143078059184, 
    0.866181510728398, 0.872283639852543, 0.861641298863653, 
    0.81571625884637, 0.775580283353865, 0.776901326470907, 0.81120667548304, 
    0.850761111795837, 0.80824175339438, 0.778983645257545, 
    0.775784859784655, 0.778231173213795, 0.802502158991794, 
    0.785114784269651, 0.715947923937295, 0.630529380310779, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.813755038460173, 0.88146008952185, 0.856575785850072, 
    0.614832745384833, 0, 0, 0, 0, 0, 0, 0, 0.49090496686588, 
    0.745391205079741, 0, 0, 0, 0, 0, 0.620033023676049, 0.488799800784976, 
    0.409744595406334, 0.772578400255117, 0.793625171513916, 
    0.87447340776143, 1.05780519450387, 1.02613957522033, 0.778109797902216, 
    0.470907920633157, 0.491141648780638, 0.628707784080484, 
    0.647359611911781, 0.499765848349517, 0, 0.311613196663686, 
    0.430961748188752, 0.504242301975115, 0.532218668296534, 
    0.572921094280516, 0.596445867280186, 0.56797296786059, 
    0.527629798331112, 0.591518902431182, 0.602850134140439, 
    0.617437153024957, 0.64837010150554, 0.643803059754241, 
    0.695975851538912, 0.749134841398148, 0.811582092371134, 
    0.835806423911184, 0.773356414832848, 0.566107992465644, 
    0.624862102640605, 0.626568597766586, 0.584001593630028, 0.6011031537466, 
    0.75363371663063, 0.854235344319205, 0.787597453908505, 
    0.885422143727547, 0.909440067490844, 0.815501042549255, 
    0.83244509395596, 0.881255573698808, 0.925945508572359, 
    0.968456394940871, 0.928045642617313, 0.884031132542767, 
    0.846803986068593, 0.774858791466577, 0.770740939108774, 
    0.730444587734584, 0.557643019517853, 0.509317223881155, 
    0.548495909561517, 0.421177946718429, 0.537182767232387, 
    0.719603538798501, 0.798280398649319, 1.32011287207115, 1.07565561082453, 
    1.14165692391404, 0.80237988157067, 0.65101965897264, 0.410232230332956, 
    0.603347975730684, 0.487426595934361, 0, 0.69843442235727, 
    0.715104316347055, 0.935680436884737, 0.928246866917078, 
    0.860956955279724, 0.823542328438264, 0.832365700841599, 
    0.819714656758368, 0.816130479008331, 0.83410073051432, 
    0.845775492227275, 0.845944383025797, 0.833828450882898, 
    0.831456053269247, 0.831631566476141, 0.811401265610328, 
    0.823898744605816, 0.817046488385182, 0.817022408986866, 
    0.823924277594444, 0.847932404071443, 0.81163523444661, 
    0.824331745801898, 0.77677237603175, 0.600119813541654, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.793832086684669, 0.840609397554274, 0.819154799546565, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.284569286514944, 0, 0.343572386805524, 
    0.534996993023742, 0.676608125049249, 0, 0, 0, 0.904898425898097, 
    0.990725732574449, 1.55735410344269, 1.09596611245097, 0.946714824335352, 
    0.821842156793573, 0.511434526270119, 0, 0, 0, 0, 0, 0.380056369742972, 
    0.562956688761054, 0.663553807093839, 0.644931136627553, 
    0.671907138613028, 0.734493199667007, 0.80058559380841, 
    0.898418057119396, 0.966482008673847, 0.985297157346092, 
    0.949963962371265, 0.872675310315975, 0.876095073594701, 
    0.899240607884016, 0.941746761520684, 0.923951753458293, 
    0.848001490316481, 0.6751953441707, 0.612990958832438, 0.573688711500097, 
    0.554205101549418, 0.591500919612381, 0.66479090983377, 
    0.744013305416372, 0.806356623651805, 0.82598198194212, 0.86443143987891, 
    0.876386450266467, 0.929069721425918, 0.970174634606413, 
    0.98840790061706, 1.01237102937906, 1.02697857520744, 1.01429899417441, 
    0.89461696843291, 0.81951617437458, 0.676004243633917, 0.58074509138568, 
    0.545737440887962, 0.498338298963554, 0.490394402191567, 
    0.748197852154657, 0.525573942929693, 1.46830876953501, 1.6471645100687, 
    1.32857481384555, 1.24892902890939, 0.90855629711949, 0.823425011981679, 
    0.749706711957173, 0.659362662326064, 0.542221935399909, 
    0.476243616973138, 0.723526484490674, 0.82977139249062, 
    0.835437898892133, 0.812455578707762, 0.837172391241141, 
    0.818893014077279, 0.802110673446958, 0.800511005834987, 
    0.80632374870849, 0.81594833258356, 0.814086091741081, 0.827616325991704, 
    0.831063417056264, 0.823411522257978, 0.83791439403676, 
    0.837698870435933, 0.805537921234822, 0.79844204916242, 
    0.812034258083747, 0.789403096242106, 0.828584702858119, 
    0.895212190364346, 0.88361401785573, 0.87787868459639, 0.906620800489615, 
    0.759292244952488, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.242757090969082, 0.445199631367539, 0.502625787960072, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.291745453214532, 0, 0.566631152921997, 
    0.610795545848176, 0.52123548774854, 0, 0.294018606914636, 
    0.941854193385651, 1.07306587214404, 1.21287811937423, 1.24056057114053, 
    1.09546949288547, 0.814469663190946, 0.55051915296641, 0, 0, 0, 0, 0, 
    0.413690206103176, 0.863971275200271, 0.946989409374653, 
    0.931820359107595, 0.877929905162422, 0.933598394028801, 
    1.05011512895295, 1.0480391680874, 1.08275941682066, 1.13159272690563, 
    1.09206071950259, 0.993555898485924, 0.772252654553805, 
    0.736207494219488, 0.72842764025612, 0.665708382676518, 
    0.676995845893499, 0.627313727285787, 0.586426393376277, 
    0.522765624209405, 0.477839551392436, 0.550833291568673, 
    0.63700178192484, 0.669892783320481, 0.718182437660371, 
    0.730983915414049, 0.812173686248354, 0.952765933514881, 
    1.04132722049283, 1.03175059546636, 1.01993546120673, 1.03996991475684, 
    1.04030782536975, 1.02248963138982, 0.974720791755453, 0.923192656101487, 
    0.749558384866687, 0.599772109638302, 0.493210728872467, 
    0.475002341853848, 0.331151636630598, 1.02780474841436, 
    0.991417181737198, 2.18326363146712, 1.97284916852003, 1.86709116039931, 
    1.52234839328484, 0.855061266575576, 0.824749109780438, 
    0.777536724858427, 0.79834395161298, 0.760720302574833, 
    0.630007995467999, 0.724419101409276, 0.817471155581394, 
    0.751388506096137, 0.741469718425474, 0.745869841402892, 
    0.739167594092916, 0.75830647429853, 0.760859970209898, 
    0.763410650057807, 0.769044137766077, 0.772810290480052, 
    0.785053364640852, 0.804658557226985, 0.817551458588247, 
    0.835824456479704, 0.829763107598476, 0.798074878079483, 
    0.779717853871172, 0.797209438519486, 0.831730658058015, 
    0.889802478910591, 0.896872390272051, 0.899910248013724, 
    0.855736902550574, 0.874633515010959, 0.855390969798301, 
    0.71362424099472, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.340384567219187, 0.313015797509433, 
    0.468799741427495, 0.157012477175666, 0.556545629100005, 
    0.691068959986922, 0.482750125166356, 0.295843666786589, 
    0.72350148730524, 0.957155576989339, 1.09935442246329, 1.18254899942631, 
    1.08170960235084, 1.21120653587313, 0.697075148635974, 0.090224347711877, 
    0, 0, 0, 0, 0, 0.64064615966433, 0.806345299164406, 0.893290884926108, 
    0.901727210675719, 0.780492622055583, 0.825555162061465, 
    0.913052405794189, 0.961820048219201, 0.978969944947194, 
    0.992353285444933, 0.964863309769842, 0.903397203642639, 
    0.867871848409445, 0.838779735800315, 0.775788647788455, 
    0.746804198254223, 0.735597253584225, 0.671176249249545, 
    0.626793156135875, 0.529469091400543, 0.424401329228497, 
    0.457775777440929, 0.581531332994405, 0.649983994265554, 0.6125359492011, 
    0.681838883120006, 0.778543484543288, 0.948956091749432, 
    1.06241892327272, 1.01892317667377, 1.01416123631349, 0.999433454947297, 
    0.998117696552819, 0.930571787960507, 0.883042796794058, 
    0.931003178377858, 0.90653016921786, 0.727051251841368, 
    0.513136510411512, 0.37390271955772, 1.19269508122103, 0.804982710111928, 
    1.93374139826436, 1.90584917138406, 2.00062156097584, 2.03193763917366, 
    1.92930871456915, 0.966615102237338, 0.851351124592094, 0.81845440690964, 
    0.754785632309726, 0.594542579198071, 0.441943619274294, 
    1.11632740790382, 0.82935636487375, 0.732609765138546, 0.686393874188426, 
    0.688576609127527, 0.689236926492076, 0.6964803148983, 0.708510090295556, 
    0.685577227292893, 0.702301342410189, 0.686102042221391, 
    0.670371427594203, 0.692325411968216, 0.697489319105607, 
    0.743902336084372, 0.779942455868336, 0.774334043475188, 
    0.735825500429442, 0.781586381574206, 0.840476745682246, 
    0.877456906912224, 0.894314179688642, 0.894686687349091, 
    0.870938319564022, 0.851641037621456, 0.901103262780792, 
    0.780417236829306, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.40629782363478, 0, 0.3394839679596, 
    0.404498195884411, 0.35784140347043, 0.476318026660609, 
    0.801289472962994, 0.50163656748401, 0, 0.757451197892093, 
    0.856475919725111, 0.674982520396469, 0.968159083449094, 
    0.836266774922643, 1.18119643682584, 1.08537348204156, 0.642313606091803, 
    0, 0, 0, 0, 0.333457891234804, 0, 0.423131708288202, 0.601852180283696, 
    0.630352978660812, 0.554980768155992, 0.712304339273336, 
    0.86250503423534, 0.940847018070348, 0.934595043524682, 
    0.973376838733001, 0.958085310209402, 0.915029758154876, 
    0.848875587731007, 0.819716094424778, 0.800442206995287, 
    0.807351210511365, 0.792710209859225, 0.732914711450219, 
    0.664649561589996, 0.548120150908528, 0.415839785094233, 
    0.343143587872145, 0.391619840453277, 0.560130813474153, 
    0.594317292665967, 0.628344653952061, 0.755446828401403, 
    0.887358063240511, 0.981131225566805, 0.954748480190086, 
    0.969655961290115, 0.928359166245687, 0.891067734928319, 
    0.841409113489119, 0.815917087328855, 0.893184117396006, 
    0.855647191523644, 0.695048151458054, 0.529954449984569, 
    0.647869260762624, 1.91484192231505, 2.10088983008018, 2.22971926888116, 
    0.990182281049287, 1.91936049123835, 2.01957078523754, 1.95555371948684, 
    1.62445585458937, 1.49077044628062, 1.24804794210859, 0.887632257859356, 
    0.58148721088671, 0.651541530312, 0.883838483222987, 0.610677206951662, 
    0.704345597263369, 0.676352669192847, 0.699507174704277, 
    0.729090243799261, 0.781572601639461, 0.808864403786841, 
    0.783213685383725, 0.764356515607614, 0.74568170204647, 
    0.713724535183221, 0.67870416009451, 0.652791021695322, 
    0.624283716614517, 0.617587149170302, 0.64187548126778, 0.6648195206078, 
    0.672541863336348, 0.771672619580662, 0.837647111636204, 
    0.845171418272861, 0.815209627540475, 0.865663149810934, 
    0.858112339997543, 0.861773359376279, 0.656668637258242, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.208916619051685, 0, 0, 0, 
    0.359931538176504, 0.59492826838812, 0.930196019124156, 
    0.824368209968663, 0.877652385534106, 0.858317131027003, 
    0.751424390060614, 0.95785156468538, 0.889768978025704, 0, 
    0.89815906335688, 1.27199986913815, 1.08546715560737, 0.96773948555895, 
    0.688186790912065, 0.421387339402377, 0, 0, 0, 0, 0.472075568390784, 
    0.326494203496157, 0.362139104545779, 0.647658133523384, 
    0.897855238819086, 0.962919299176562, 0.937448001972265, 
    0.932273938830177, 0.924169390945572, 0.88544745375204, 
    0.838001008550002, 0.864987761435166, 0.881512091710038, 
    0.876798087537239, 0.861791246609721, 0.789676749372544, 
    0.697034815224819, 0.626385886610557, 0.504844268287453, 
    0.524746444068598, 0, 0.344129860392884, 0.560701672366581, 
    0.629796329532061, 0.649658611662017, 0.855024453187264, 
    0.920895465865313, 0.914258251205781, 0.81568288057903, 0.79109671639576, 
    0.760583425967697, 0.716742864721313, 0.732349282932342, 
    0.759685068435296, 0.777035917828113, 0.596889555177898, 
    0.650529234691716, 1.7430003639875, 2.12208422104965, 2.11573887827011, 
    2.13125856161755, 1.56049470626607, 1.97308874303991, 2.02852508310691, 
    1.95320447845053, 1.89100068525637, 1.79129523079092, 0.862572788929231, 
    0.347913547923936, 0.664155938072508, 1.12969261000788, 
    0.734071374575864, 0.434472476905052, 0.399709528240592, 
    0.415472339250587, 0.428440637794814, 0.567168268401927, 
    0.686608681262336, 0.727350858209634, 0.678123760353774, 
    0.634841952507673, 0.652388759576251, 0.641442695904298, 
    0.543357690133145, 0.524717388107029, 0.52742716969867, 0.55175381303445, 
    0.603371989362199, 0.57176383852018, 0.523855688304499, 
    0.637486430847304, 0.771022688882192, 0.803790168999615, 
    0.835551666866076, 0.864587868563251, 0.941321701530855, 
    0.887200145328847, 0.56232945455521, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0.475063183006242, 0.481231624526117, 0, 
    0.306124667436074, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.478992412716188, 0, 
    1.09330712610398, 1.1800852688262, 1.30616873314181, 1.41069285066407, 
    0.762102329386101, 0, 0, 0.658560043195563, 0, 0, 0.803696745057605, 
    0.588657627309461, 0.495607698448238, 0.341178714119344, 0, 
    0.497797606966999, 0.659381850795448, 0.248484053312316, 0, 
    0.504242731266022, 0.786650710628632, 0.862941535804496, 
    0.862122285159864, 0.84515323224145, 0.85034624807251, 0.817367648537382, 
    0.831768563500386, 0.876001923128406, 0.880873388986771, 0.8518232897974, 
    0.860910372569106, 0.834931326761668, 0.730878508402374, 
    0.642077174815046, 0.535954674375527, 0.460605993938585, 0, 0, 
    0.399556746289916, 0.487049069280769, 0.601519259092471, 
    0.839674758694643, 0.862608490089693, 0.797976673363066, 
    0.759998025472836, 0.761543504481508, 0.728950941122985, 
    0.681707181328689, 0.586825001600681, 0.67284270775736, 0.60506847800847, 
    0, 1.16363780766022, 2.14767192926819, 2.14426962677168, 
    2.14209767661754, 2.15236863447488, 1.93315549949477, 1.64710428447701, 
    1.98104955809288, 1.93529315524039, 1.85685800262087, 1.26190595692144, 
    0.668670564548701, 0.353685768937919, 0, 0, 1.29638688228373, 
    0.35818847296134, 0.378630579097404, 0.391367261655669, 0, 0, 
    0.342223450887241, 0.527888182053695, 0.488851165109113, 
    0.317683446105892, 0.423860576123488, 0.491989039278379, 
    0.409279860602341, 0.414252168507009, 0.439719115263257, 
    0.453730074094046, 0.394729294073266, 0.463659980695984, 
    0.506853556319771, 0.538541448827207, 0.63792878919269, 
    0.709702414486014, 0.762780125399875, 0.874561709996681, 
    0.962646404627411, 0.874141831521944, 0.80540140861715, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0.377515174848656, 0.364445708389554, 0.472743250475834, 
    0.417163520262447, 0.351079999964872, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.206050038601655, 0, 0, 0, 
    0.408933675027859, 0, 0, 0, 0, 0.889835991312848, 1.22429744371427, 
    1.33808459642673, 1.33149137970481, 0.210982098515044, 0, 
    0.985759988321688, 0.930542870064705, 0.587973190517379, 
    0.944678454733382, 0.809023381389697, 1.19005075218064, 
    0.803253033546461, 0.429470936366502, 0, 0, 0.710430255531044, 
    0.645727614419753, 0.44265562738381, 0.441853173996532, 
    0.627713424285186, 0.733956595231321, 0.744739908875796, 
    0.752907781238306, 0.741365782392092, 0.70972873571821, 
    0.745396758907601, 0.813990689403119, 0.802637916661387, 
    0.762203141616509, 0.738805590359998, 0.761703715635452, 
    0.755329022348298, 0.688442378934345, 0.580201895864355, 
    0.340661527251058, 0, 0, 0, 0.269189539158446, 0.600353575965674, 
    0.759416909866241, 0.739765419691655, 0.764950954778877, 
    0.742563481048563, 0.735013697729786, 0.704629864367841, 
    0.677525336849638, 0.569757470746817, 0.711975290337774, 
    0.464733404114093, 1.32785893292901, 2.34004980294758, 2.28309737512484, 
    2.20072825864738, 2.20001823800518, 2.26250381634843, 2.18654367997186, 
    1.46483932689259, 1.77971856193853, 1.41817612978799, 0.558548658939258, 
    0, 0.399844586264614, 0, 0, 0, 0.860883009589428, 0, 0.344068617345628, 
    0.929452378494558, 0.881789829009102, 0.658418892220673, 
    0.416516454019923, 0, 0, 0, 0, 0, 0, 0.415181795957479, 
    0.476539185805461, 0.410330279645415, 0.312605758021483, 0, 0, 0, 
    0.487174140397166, 0.585609264253109, 0.622992484093697, 
    0.739306068514371, 0.830639105017189, 0.877514121702318, 
    0.88212081527006, 0.638787583317201, 0, 0, 0, 0, 0.422496378394821,
  0.808857921312309, 0.508974389977537, 0.638941861716778, 0.530308782988123, 
    0.200433255684458, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.794761186977073, 1.41219844052656, 1.27947316436684, 0, 0, 
    1.3854753158857, 0.811384006450157, 0, 0, 0.738790618300339, 
    0.873616700179617, 1.06647712769808, 0.532822319836491, 0, 0, 
    0.615658778808681, 0.696235356198346, 0.573009448246069, 
    0.532902743746475, 0.572388601751445, 0.579904856308574, 
    0.662909536243405, 0.674937668846386, 0.645250404221645, 
    0.646890812595515, 0.685233202676356, 0.724181289624284, 
    0.688247642821901, 0.622186417654744, 0.573716214662113, 
    0.626923291999184, 0.672277932591648, 0.685969937756444, 
    0.647208958564505, 0.473371890069749, 0, 0, 0, 0, 0.528933061798221, 
    0.646693447893175, 0.702553193719837, 0.678990817095415, 
    0.685552002160277, 0.72838624231534, 0.675563350030686, 
    0.623063705661353, 0.580633754615814, 0.462172264619684, 0, 
    2.08664500761333, 2.36393894351356, 2.30849117361557, 2.23690413208823, 
    2.27594154290945, 2.234846019497, 2.22650830558514, 1.59405354121772, 
    1.24247104407457, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.504215866081263, 
    1.04034646879086, 1.242686617664, 1.26615537839447, 1.02547521794419, 
    0.130675426591011, 0, 0, 0, 0, 0.345412120820541, 0.377493999360797, 
    0.388250363667587, 0.362963578169777, 0, 0, 0, 0, 0.39050041450866, 
    0.547836134407514, 0.622528098054061, 0.694550415080564, 
    0.777542125458795, 0.775685193709362, 0.647246107478764, 0, 0, 0, 0, 
    0.286442353332305,
  0.727737671351554, 0.743041327693401, 0.719360966250557, 0.520540199505984, 
    0.565060423105441, 0.383032479966937, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.800686453080257, 1.07303802583154, 0.878394324945334, 
    0.480852752519259, 0.480531432188867, 0.808148997894816, 
    0.991552578720049, 0, 0, 0, 0, 0.179461461000289, 0, 0, 0, 0, 
    0.393565970830572, 0.442332458503142, 0.426623250054116, 
    0.42575758177609, 0.400388641896016, 0.509616790409677, 
    0.582628794009534, 0.567186033056656, 0.546166526785732, 
    0.576228234357071, 0.588371641872348, 0.590419437277851, 
    0.523186292013068, 0.453037561007217, 0.457774711528388, 
    0.536965198987684, 0.616960088995317, 0.605713624000549, 
    0.443554686748857, 0, 0, 0, 0, 0.453838491499867, 0.599646779552813, 
    0.629493693661409, 0.606774503456427, 0.65431510048964, 
    0.635821397083749, 0.602682762151845, 0.581187719089356, 
    0.571006978350652, 0, 1.62564818595292, 2.35004794660666, 
    2.35818388661094, 2.3221083988381, 2.25238759031845, 2.27449039648466, 
    2.2841916561305, 2.08134211270636, 0, 0, 0, 0, 0, 0.634214832439681, 
    0.506894913444816, 0, 0, 0, 0, 0, 0, 0, 0.97871389567374, 
    1.24673206036062, 1.37653971389908, 1.25228158807997, 0, 0, 0, 0, 0, 
    0.429678420922318, 0.443832950127346, 0.382950587777583, 
    0.306573619601423, 0, 0, 0, 0, 0.391376776117896, 0.474927256431083, 
    0.530522134600055, 0.598815593170245, 0.629320380279151, 
    0.730165499269998, 0.53737851196665, 0, 0, 0, 0,
  0, 0.209273906149892, 0.386472857332915, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.353276687917658, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.05323078763281, 0.895736319814274, 
    0.32221818800239, 0, 1.15414581491114, 0.701964197536939, 
    0.734006103752661, 0.183713095728753, 1.11400319157109, 0.88917055624895, 
    0.768983504478775, 0.190464840088719, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.260497136929882, 0.350189063668023, 0.361281831705734, 
    0.375316255776129, 0.384710316433313, 0.454866877079887, 
    0.419697448295945, 0.472612570127021, 0.516115689277909, 
    0.541830851604621, 0.546972044629326, 0.40051518466645, 
    0.308472923047164, 0.383370430355844, 0.35278942139203, 
    0.429491714344108, 0.399047721508272, 0, 0, 0, 0, 0.571398927520516, 
    0.576381976889856, 0.545524022807211, 0.541573993564283, 
    0.58436243119267, 0.619365871264221, 0.590299260001547, 
    0.555700453696507, 0.547665807322224, 0, 1.90649904500527, 
    2.53247474604074, 2.07341221109574, 1.98183410957383, 2.30906769036989, 
    1.50510174180924, 1.15808324089172, 0.835125532683549, 0, 0, 
    0.598163537894439, 0, 0.609706736756547, 0.663622426175335, 0, 0, 
    0.350701160409277, 0.399845783575979, 0, 0, 0, 0, 0, 0, 
    0.861527593083548, 0.998317398445672, 0.741265159603177, 0, 0, 0, 0, 
    0.743921465655538, 0.699017587038197, 0.484689164074929, 
    0.329774671758864, 0, 0, 0, 0, 0, 0.281751303023251, 0.354242940907249, 
    0.413433733880154, 0.500913712029291, 0.586200259355925, 
    0.480147445816727, 0, 0, 0, 0,
  0, 0, 0, 0.129411228555596, 0, 0, 0.352805127034772, 0, 0, 0, 0, 0, 
    0.282784177866278, 0.245518598075898, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.08289340173369, 
    0.731381791977472, 0.299246171724598, 0, 0.180275030737542, 
    0.928334404181646, 0.642350232024838, 0.883734840406911, 
    1.05638862788331, 1.22346704439161, 0.86091899767485, 0.835968286199209, 
    0.786246828664195, 0, 0, 0.397787188686794, 0.672048177329608, 0, 0, 0, 
    0, 0.247252518311671, 0.241551100975018, 0.173107434880391, 
    0.225276836620797, 0.277922625504683, 0.338770491874782, 
    0.404267170939965, 0.432697770170657, 0.46024154652712, 
    0.466108651960854, 0.502879007843992, 0.489156803248638, 
    0.456813895775083, 0.263440683257121, 0, 0, 0, 0, 0, 0, 0, 
    0.194170679353888, 0.416600317527482, 0.423258832180593, 
    0.401512160356882, 0.476069703537377, 0.546243984777409, 
    0.59094946326099, 0.62113672603347, 0.595026009967987, 0.565123710281366, 
    0.472149833663828, 1.84060149813668, 2.35806033197402, 1.73497984806357, 
    1.81306555748547, 1.76139737706669, 1.87602488662153, 1.49318306049567, 
    1.18977827973295, 0.879213740242837, 0.900955515662361, 
    0.967112630490361, 0.935727080016095, 1.06229959286822, 0, 0, 0, 
    0.344875490286618, 0.733510318764518, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.750878933232747, 0.809759848801816, 0.777846518188476, 
    0.469562677426803, 0, 0, 0, 0, 0, 0, 0, 0.172028660604198, 
    0.158995742654819, 0.354898953825987, 0.358138210487672, 
    0.270831117266148, 0.30277760446416, 0.467206752119211, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.02917615827575, 
    0.807410771085054, 0, 0, 0, 0, 0.830401583351746, 0.60885958365018, 
    0.916207796902541, 1.28285574728874, 1.21303673191127, 0.700568621299711, 
    0.761647970076489, 0.69975460970557, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.207653590964885, 0.278284758165304, 0.324629487533863, 
    0.390515242120562, 0.433540749461913, 0.431477261378763, 
    0.363924127071451, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.199978083447782, 
    0.284176540783847, 0.356198626112582, 0.442310217970728, 
    0.52450219454863, 0.600434488444862, 0.592745782810264, 
    0.639137703612061, 0.647283568531075, 1.52439604850157, 1.4399058062969, 
    1.54161787374149, 1.79392236292137, 1.58445747036149, 1.50535613577067, 
    1.40124257486919, 1.3937221023396, 1.19538769225224, 1.12658819781201, 
    1.05182767192257, 0.767226756513029, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.67650114910134, 0.838605530232929, 
    0.805427204011987, 0.642095618612763, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.209554640910489, 0.391298725558531, 0.559805221170811, 0.442416683878938,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.606931074872642, 
    1.02036177190014, 0.862842290205674, 0, 0, 0, 0.43123571009909, 0, 
    0.977987540842204, 1.32938085337247, 1.10860272847751, 1.01954619696564, 
    0.785953030294517, 0.47039531979879, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.306547934029772, 0.376046548998852, 0.311609616694099, 
    0.294334925829223, 0.133745822528021, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.233240526194208, 0.348535932689952, 0.423101901516316, 
    0.544666069311222, 0.564933019982108, 0.609922617781462, 
    0.463171503956276, 1.45403855153618, 1.64376479706158, 1.50700707285532, 
    1.45683682022436, 1.49536390682277, 0.867357563620988, 1.15530470319991, 
    1.31721695830656, 1.36333418598836, 0.939977016579679, 0.515257067274866, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.613969094948458, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.527623418203711, 0.773397260984106, 0.833679387344595, 
    0.607165982112973, 0.302499693703191, 0, 0, 0, 0, 0, 0, 0, 
    0.0471686187998361, 0.33211981917308, 0.132704377180659, 
    0.329725565300129, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.864636047812148, 
    0.973117925781167, 0.362845041108324, 0.853588098201764, 
    0.752321148877674, 0, 0, 0.276461012262908, 0, 0.835556963697866, 
    0.952038533396189, 0.862244016255062, 0.807699827445394, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.228748621424788, 
    0.403937523804386, 0.453432390352234, 0.294903101721068, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.383548544747889, 0.522707840526261, 
    0.526307845935976, 0.765077464439675, 1.71666250407778, 1.65527732211244, 
    1.35587697900036, 1.51380610042054, 1.40069963797763, 1.10250549483412, 
    0.823258141286468, 1.15712970308496, 1.2304886608872, 0.762266330449571, 
    0.493093493538001, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.715647172318758, 0.633437127670383, 0.497144878949338, 0, 0, 0, 0, 
    0.39850496403927, 0.464251590454802, 0.676262665846065, 
    0.449702580839683, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0986786952170912, 
    0.257201365508933, 0.30828860996233, 0.462114525508758, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.410449662907932, 0, 0, 0, 0, 0, 
    1.06476354922666, 1.2154208362294, 0.904568017523874, 0.633456990819506, 
    0, 0.541118849779526, 0, 0, 0.649480688966909, 0.683268288474428, 
    0.856934556295022, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.174024522100245, 0.4942132003171, 0.453725664229245, 
    0.30363424417723, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.396305465731762, 
    0.506920168851774, 0.616451617944297, 1.15637673892763, 1.56885671182689, 
    1.28129592101444, 1.39082649395465, 0.812034391960959, 0.439356545051629, 
    0.750747826538489, 1.00564302741803, 0.954742195979852, 1.00877462872077, 
    1.10078863479596, 0.980003053909557, 0.74122101121449, 0, 0, 0, 0, 
    0.55198531651636, 0.567005443999427, 0.62121247418291, 0, 
    0.505620051907383, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.483852292400771, 
    0.269105906736878, 0.390922651379795, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.305885705007347, 0.343260501523528, 0.266590775710774, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.180515473409564, 0.411341773976054, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.646894126513745, 0.458156655167334, 0, 0, 0, 0, 0, 0, 0.73287081701812, 
    0, 0, 0, 0.644567476845983, 0.8637194716798, 1.13632359774697, 
    1.20956120687815, 1.24033489520648, 1.14820388416532, 1.15038584915231, 
    0.773820344566106, 0.854224065614795, 0, 0.526333154109202, 0, 
    1.22469187274628, 0, 0, 0, 0, 0, 0, 0, 0.570984223095539, 
    0.798015192490218, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.522350038587425, 
    0.806315441056339, 0.403239272682041, 0.76069531983342, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.271576401627218, 0.483033974718349, 0.453197445072223, 
    1.06832215339625, 1.98834935179822, 1.32935729872136, 1.3509362949763, 
    1.41361645448791, 1.5176121843882, 1.4102333603769, 1.19067510130922, 
    1.07406922473001, 1.05759270841437, 0.847819801723542, 1.81350520598685, 
    1.15086461753049, 1.69574611389922, 1.14615675537675, 0.764586470009472, 
    0, 0, 1.15907014413449, 1.33823817632697, 0, 0.661836891974984, 0, 0, 0, 
    0, 0, 0.680832269291561, 0, 0.413756674032635, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.430841659102671, 0.409706993554218, 
    0.231862995384511, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.783003837275633, 0.73006622974775, 0, 0, 0, 0, 0, 
    0.72015539350348, 0.67496801070607, 0.375820517228677, 0.616135987389328, 
    0.862723741258861, 0.16352039529592, 0.576498227615313, 0, 
    1.09252321933124, 1.49870375369756, 1.34857118594647, 1.31046968140271, 
    0.847128407334532, 0, 0, 0.387862915370859, 1.10904004694039, 0, 0, 0, 0, 
    0, 0, 0, 0.587640849000488, 0.982140695278635, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.492768518440369, 0.50349435041748, 0.805430336063184, 
    0.842957468505571, 0.605146159451575, 0, 0, 0, 0, 0, 0, 0, 
    0.454263870160613, 0.485528844558065, 0.987409500724152, 
    0.899629054245325, 1.20551139350574, 1.42480648316539, 1.35613746386078, 
    1.3038939544822, 1.29663940776679, 1.15045569868226, 1.02314532480607, 
    0.601738944294606, 0.7465506345477, 2.05512458494098, 1.97825828125206, 
    1.98449211818044, 1.45440419522199, 0.813244022377763, 0, 
    0.794921500987495, 0.530598514483292, 0.895773459057859, 0, 0, 0, 0, 
    0.833279232241648, 0, 0, 0.90832873673453, 0.579643425736743, 
    0.0330678534726228, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.210274734669208, 0.331770411928348, 0.401211131083983, 
    0.147259517415412, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.823544806853553, 0.985075878545547, 
    0.622970766623854, 0.758238429408754, 0.627230107018409, 
    1.00386344888727, 0.539428399555812, 0.991670400958024, 1.08059023550279, 
    1.18923439477754, 1.03910144212073, 0.423001752314344, 0.442060723159844, 
    0.201246271203921, 0.347825889322398, 1.13155303156074, 1.46625204491705, 
    1.55689702123059, 1.4935060728954, 0.817119510860392, 0, 
    0.663316305271452, 1.81960721834515, 1.89147837599349, 0, 0, 0, 0, 0, 0, 
    0, 0.573255696227964, 0.879606512064103, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.435693526097547, 0.731573864280402, 1.51117802755681, 
    1.39400469379895, 0.551110012022924, 0, 0, 0.295294433176925, 
    0.441444442105993, 0.532529269450467, 0, 1.01536085815006, 
    0.846453936750412, 0.80325103100942, 1.5192191520509, 1.61291264832304, 
    1.79308341693499, 1.51084682476949, 1.52089517763439, 1.23305853479365, 
    0.668244482805888, 1.77799177260845, 1.66998777367918, 1.54710238783779, 
    1.64143278372294, 1.85933403899109, 1.08846541039676, 1.20182417042165, 
    0, 0, 0, 0, 0, 0, 0.748785939103275, 0.496658922820853, 
    0.436775203235454, 0, 0, 0.76101246621342, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.116649426902692, 0, 0, 0, 0, 0.444213464059909, 
    0.574209004930512, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.992124478951638, 0.571894278384552, 
    0.680923354596536, 0, 0, 0.640882533368811, 0.951021855079683, 
    0.778599799235813, 0.969070310117053, 0.974895288818441, 
    0.740490441490161, 0.948506373849508, 0.932016645209942, 0, 
    1.00771390255782, 1.30492595455433, 1.37443011677932, 1.37005781210673, 
    1.11182898201669, 0, 0, 0.86720034882421, 1.22816590485422, 
    0.679431141771518, 0.73001339698843, 0.742938908379866, 
    0.591860739955784, 0.266860829779501, 0, 0, 0, 0.683848069818877, 
    0.505976169755278, 0, 0.398196106594058, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.929739443652492, 1.47938614158537, 1.60143535879478, 1.57984691397149, 
    1.4893225046677, 0.991644693400504, 0.312462465128433, 0.94991529526606, 
    0.518077395039241, 0.601602913344635, 0, 0.817501273906397, 
    0.832326546960178, 0.629968024118155, 0.821016995084694, 
    0.841995490139953, 1.16412107701241, 2.1774089911578, 1.53485763588035, 
    2.11792311225201, 2.07557115058761, 2.07396981170859, 1.38384297010336, 
    1.33871022235293, 1.44079942344893, 0.961477073509679, 0.83239022555548, 
    1.2006835958932, 0.421404149992984, 0, 0, 0, 0, 0, 0, 0.753722147755645, 
    0, 0.847616671195422, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.129905917347402, 0.569843795108482, 0.550335945060939, 
    0.555211947069508, 0.494545647350979, 0.436436112812523, 0.480883057506564,
  0.418115813014633, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.96630429307536, 0.684892373001109, 
    0.886148400098633, 0, 0, 0, 0, 0, 0.348538363656214, 0, 0, 0, 0, 0, 
    1.01984082586837, 0.979328221014745, 1.18362698816251, 1.36969890496747, 
    1.52569615236312, 1.44743888802424, 1.1750659087291, 0.793288030726268, 
    0.887643463031128, 0.601529660515969, 0.677422384352821, 
    0.495999588004283, 0, 0.155362603477054, 0.486341761268927, 
    0.32759202141266, 0.223830570084074, 0.373810959193897, 
    0.144196420160337, 0, 1.44824867730791, 1.66249976793306, 
    1.87086289550199, 2.01082385020388, 2.15745772409085, 1.24377407197064, 
    0.807698896146926, 0.941930684930098, 0, 0, 0, 0, 0, 0, 1.29597589900224, 
    1.64534202097608, 1.69077231763906, 1.57179903399501, 1.95155587774746, 
    2.04368499897312, 2.01158439422387, 2.14656672082012, 2.17750422636652, 
    2.3647586337362, 2.37509814973006, 1.27287715769283, 1.33700361595024, 
    1.25860893716637, 1.01202402766579, 1.01720473879588, 1.604926702461, 
    1.92011276283106, 1.94041323560522, 2.1628107418597, 1.34158822038269, 
    2.08246773262755, 0.466149494658989, 0, 0.469939992295519, 
    1.57268635599537, 0.809287814212711, 1.39233033481725, 0.747622468481815, 
    0, 0, 0, 0, 0, 0, 0, 0.531752113644399, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.313329149932227, 0, 0.489816999064566, 
    0.617508318220538, 0.695625597071877, 0.639551859058294, 
    0.425249444169908, 0.474525816843076, 0.441767201002785,
  0.32282508803849, 0, 0.352385299660397, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.828768843421481, 0, 
    0.176426575232831, 0.865888316009155, 0, 0, 0, 0, 0.578652398014771, 0, 
    0, 0, 0, 0.778900880098397, 0.779888400121338, 0, 0, 0.393583385933839, 
    0.581448595588134, 0.637446420288259, 0.493362655873655, 0, 0, 
    0.889210915691181, 0.627779052113957, 0.734546807327458, 
    0.766968270170257, 0.798302222091877, 0.725443946618294, 
    1.27114116624166, 1.87706502381659, 2.07189244787606, 2.19342072847061, 
    2.16790977230995, 2.23392776435398, 2.2532219355607, 2.34970763225107, 
    2.37601283834135, 2.35927085950485, 2.39385154628818, 2.3896487693584, 
    1.8144354042631, 0, 0, 0, 1.03721016840962, 0, 0, 0.895462822735781, 
    1.34403685624233, 1.42007311164056, 1.47883346732355, 1.41268255127718, 
    1.64101621135865, 1.65104375791258, 1.68063424643746, 1.88257385050174, 
    1.80912315838891, 1.96705082422858, 1.56451434503912, 1.48414908387384, 
    1.37763175153214, 1.5620009994284, 1.25197243022342, 2.0065577668909, 
    1.52895517572646, 1.55253396174874, 2.15693069912539, 2.10694071760913, 
    1.34303587580857, 1.04984516778419, 0.781478409530096, 1.06717189545264, 
    1.51529942678795, 1.41897277691856, 1.40709209834011, 1.04273655235022, 
    0.959256765524774, 0.479938123000697, 1.05915023922294, 
    0.878413235446985, 0, 0, 0, 0, 0, 0.491203418412783, 0.80912229559359, 
    0.479739961964054, 0, 0.160614487887996, 0, 0, 0, 0, 0, 0, 
    0.365814361559546, 0, 0, 0, 0, 0, 0, 0, 0.197516103900903, 
    0.202965998221929, 0.388268260471462, 0.436781177955587, 
    0.73648131717751, 0.793850043757902, 0.799451954057269, 
    0.631046424889281, 0.619783460169391,
  0.798629864916664, 0.189551982554303, 0.328393428207466, 0, 
    0.25194134962244, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.792036729254814, 0, 0, 0, 0.865018035200041, 0, 
    0.649150033096037, 0.830561514787585, 0.901524961139088, 
    0.537517340499382, 0.894575174629027, 1.07230724061426, 1.0491845837409, 
    1.09656877073565, 1.20171626284088, 1.18828596356306, 0.50187992128919, 
    0, 0.618572727719451, 0.855077464878052, 1.33676738400695, 
    1.50726875022983, 1.0859444769563, 0.624583152982515, 0, 0, 
    1.90598338481354, 1.98346659995463, 2.07252346552873, 2.22198686002982, 
    2.12180849988847, 2.19867416698108, 2.31555817423439, 2.39310048943231, 
    2.39162535179887, 2.21329298750839, 1.98324770242615, 1.81743070644817, 
    1.64992284641066, 1.7046296017986, 1.86535650707028, 1.86325734539693, 
    1.29433316001517, 2.14250961997961, 2.16713631359958, 1.85989458067048, 
    0, 0, 1.00392941486083, 1.53706584145712, 1.46563472639859, 
    1.44435795778561, 1.30312588602021, 1.59824037245823, 1.74167991091066, 
    1.58137634050474, 1.68019426259125, 1.61518204689703, 1.81451150763972, 
    1.98080396327685, 1.9812260211038, 2.01405461480322, 0.715042460681278, 
    1.58448707802505, 1.65887086571472, 1.49220110625901, 1.31846949102239, 
    2.02983232762252, 1.9803016729373, 1.91477484565765, 1.69759595002897, 
    1.21288177741761, 1.29840889760767, 1.64313866796112, 1.60112490262672, 
    1.48011792093723, 1.0790935282129, 1.1910970951911, 1.02553433800616, 
    0.882040885240588, 0.763946127706448, 0, 0, 0, 0.339669872394087, 
    0.838427619827704, 1.23576481854806, 1.32432960073087, 1.17719318673113, 
    0, 0.509003414742785, 0.547858915569477, 0, 0.69382730559253, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.362645990363906, 0.621519586651759, 
    0.775488354281188, 0.863586933124369, 0.943544231148197,
  0.884057874868765, 0.806510305171356, 0.453014689933656, 0.246304822772519, 
    0.206906917568012, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.423161353182703, 0, 0.375220886440416, 0.663341838870819, 
    0.616521928286821, 0.546463859608579, 0.675143548050848, 
    0.468221846749257, 0, 0, 0.680703287045871, 0.78891006099135, 
    0.702494182854326, 1.04895291833473, 1.09146182054622, 1.05793941242631, 
    0.989707403517689, 1.04426522577567, 1.80551370142226, 0.973516779816798, 
    1.0567071392214, 1.12321132807055, 1.09015260729193, 1.19887069118675, 
    1.19579799272591, 0.820073853172606, 1.62895938842225, 1.81215434265152, 
    1.81483544176377, 1.70967566826896, 1.96775545153324, 1.90475590306264, 
    2.10637188057188, 2.11829767679954, 2.21859963960881, 2.13085410115426, 
    2.14215641028123, 2.16521268987342, 2.17438674992072, 1.99456668618785, 
    1.38145640509351, 1.21041018808359, 0.941175174537133, 0.982360235570439, 
    0.917872896074701, 0.911168618760393, 0.928228714497991, 
    1.21238046162501, 1.18187857217337, 1.38518869792583, 0.721443011522476, 
    0, 0, 0, 1.32336468469869, 1.41049486102805, 1.48350003641235, 
    1.34178850563546, 1.17841465893897, 1.27977939780003, 1.47095703655348, 
    1.57562881199924, 1.57233381617741, 1.89259908690922, 2.08971177617084, 
    1.94775984924141, 1.40629913854743, 1.32833979794485, 0.860548305840854, 
    0.46696855327118, 1.1425370084782, 1.296748081198, 1.37137823801043, 
    1.46923141498009, 1.60255332241842, 1.45018243608205, 1.43151062458787, 
    0.864403384876465, 1.32606014953272, 1.60595035692605, 1.84497571099236, 
    1.26363310914788, 1.21644752910299, 1.30506801855905, 1.16719334567088, 
    1.09436192614067, 1.33776209289867, 0.566012558268365, 0, 
    0.295732276192871, 0, 1.0144457628335, 1.37038690042534, 0, 
    0.770665688106074, 0, 0.372278358035854, 0.545464244517327, 
    0.447013448494961, 0.804034231722806, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.356392357116828, 0.264227483757681, 0, 0, 0.442063815310363, 
    0.691590593523407, 0.834267485480339, 0.893415173043181,
  0.84843509347782, 0.824592565191417, 0.750527640062474, 0.661919990060255, 
    0.55205634754146, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.274627145787236, 0.25254146537008, 0, 0, 0.615491191172187, 
    0.417094532072034, 0, 0.309922616847417, 0.638555969699837, 
    0.736605184792509, 0.932136979137486, 1.05279156499436, 1.15030620718528, 
    0, 0.545529915135715, 0.932884653081175, 0.728134918051786, 
    0.770698386125257, 1.00641757488477, 1.17602612407716, 1.06460857612169, 
    1.05545287194103, 1.06847768580364, 1.09095525006132, 0.875058428823372, 
    1.10023919533748, 1.15137669406313, 1.2032313594137, 1.21093214957482, 
    1.14536897950443, 1.76158581027784, 1.70442391828883, 1.69866068711571, 
    1.8478644933161, 1.81765658948267, 1.88153020418745, 2.07047176090617, 
    1.96473850348842, 2.1074252680019, 2.12119164108535, 2.05979275705926, 
    2.02473355331702, 1.69802912144135, 1.4005430397118, 1.00937736834568, 
    0.966440970608919, 0.971974255422632, 0.48381190571837, 
    0.706023116965373, 0.761330103080397, 0.861446064328877, 
    0.592929018488435, 0, 0, 0, 0, 0, 0.355956409446735, 0.512318531352599, 
    1.04391686634407, 1.16514196171462, 1.22450679896314, 1.51969481781845, 
    1.26425845376604, 1.40727115572094, 0.946972531979871, 1.45877119341196, 
    1.01946279052591, 1.23728281367092, 1.02306485942942, 1.01447569725291, 
    1.02759157234004, 0.934998576283456, 1.13249409297274, 1.05240389925385, 
    1.04393967749565, 0.578604869900531, 0.83173660908735, 1.2514349943487, 
    0, 0, 0.731020696939055, 1.28595862741323, 1.62672859097816, 
    1.71224042734027, 1.73235301957615, 1.38994299186006, 0.953800248086644, 
    0, 0, 1.54978452425799, 0.831507812514336, 0.526883092093257, 
    1.19446724044593, 1.4767449239109, 1.33925571034502, 1.05335931793111, 0, 
    0, 0, 0, 0, 0.694898622534892, 1.02385578277887, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.359982024617506, 0.632318635714687, 
    0.721177933318381, 0.776470143890816, 0.832158933137705,
  0.734026885263166, 0.779167506742211, 0.800797591646964, 0.914798946510683, 
    0.986439849316817, 1.05723317661581, 0.98462105574485, 0.906361288999611, 
    0.86606332620302, 0.77515446530631, 0.627308099642264, 0.648950833914014, 
    0.722848722511619, 0.528232095331631, 0.443480798062677, 
    0.376085364208517, 0.36768573606686, 0.162255569008149, 
    0.233687054236495, 0.353399456901776, 0.410693995594001, 
    0.58994484106241, 0, 0, 0, 0, 0.0353314793947282, 0.715899631388578, 
    0.613474596304396, 0, 0.304242178128745, 1.18771413335934, 
    1.2606033448744, 1.25703359208151, 1.02719630561787, 0.778862055247647, 
    0.922429633564582, 1.16395131590112, 1.21656233108672, 1.1710730748358, 
    0.984329867468383, 0.966773846960242, 1.02810447999506, 1.08808202660526, 
    1.0348010792719, 1.11527937484332, 1.57315106166965, 1.51611651517078, 
    1.71596682638935, 1.65719111619306, 1.62259353428676, 1.62605923643886, 
    0, 0, 0.448141022452889, 1.10680550300841, 1.37355074944709, 
    1.56327140961689, 1.72764946215215, 1.83097854819972, 1.13672278114929, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.617332989870159, 0, 0, 0, 0, 0, 0, 0, 
    0.312852524693037, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.816004405490157, 0.856169662162374, 0, 1.16755834817497, 
    0.864154679158579, 1.14804964536135, 1.72659504166002, 1.906703323688, 0, 
    0, 0, 1.43348996076786, 1.48174080634551, 0, 1.17267015956658, 
    1.50810146264232, 1.56426963962572, 1.53935548342885, 1.53553038759183, 
    1.49406480804051, 0.680193264139884, 0, 0, 0, 0, 0, 0, 0, 
    1.06051623609426, 0, 0, 0, 0, 0, 0, 0.382076195617944, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.352464647468272, 0.493806239941587, 0.55057943038431, 
    0.655851805639522, 0.730658014905998,
  0.678653399164859, 0.716044606875118, 0.723796068038415, 0.811277167510858, 
    0.851900984036124, 0.844335067496154, 0.756929312981454, 
    0.652690916061164, 0.540532972065487, 0.439942200714593, 
    0.428022531123965, 0.501066612219028, 0.482369415239858, 
    0.379075634638297, 0.243366417772918, 0.182348997757657, 
    0.358284055316841, 0.339766281265469, 0, 0.35683208905566, 
    0.249489277312108, 0.708781889649716, 0.555957959872279, 
    0.473619381312065, 0, 0, 0, 0.376506255547894, 0.471954783551427, 0, 0, 
    0, 0.992185725934206, 0.764893285988446, 0.658377245229414, 
    1.20345120401751, 1.14497249987611, 1.00427942349803, 0.995743344369722, 
    1.05953180499379, 0.920504638670494, 0.829295732393265, 1.10420686805902, 
    1.35073475789375, 1.51435238528149, 1.38538759788128, 1.40746152885404, 
    1.11343980555912, 0, 0.729678096504767, 1.10079625739784, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.756289962847804, 0, 0, 1.19981927512767, 1.13251072284307, 
    1.28106218741943, 0, 0, 0.787007919477107, 0.943383461535107, 
    1.12821249465979, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.661886911179939, 0.71243590725595, 0.296126287324277, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.493390172784373, 0.61665436964833,
  0.381368899761528, 0.591978991479905, 0.752028823109091, 0.904098772969815, 
    0.893837312239348, 0.613345931432977, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.326277734002365, 0, 0, 0.397225758522128, 0, 0.43484793361461, 0, 0, 
    0.156513034936976, 0, 0, 0, 0, 0, 0, 0, 0.64167330815193, 
    0.555895592503428, 0.809107721452746, 0.739014331449301, 
    0.698941675561843, 0.809787152268747, 1.18947800669674, 1.05340358276454, 
    1.05651144482533, 1.09868573033512, 0.970717950819677, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.557669732691767, 0, 0.433087685588831, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.575291427959538, 0.966104097304706, 
    0.806933704143338, 0, 0, 1.2559390956026, 0, 0, 0.900702204804406, 
    1.29641727411563, 1.21732519523591, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0.476426870076039, 0.678326037292369, 0.654980421722516, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.209324748862118, 0.244008975656911, 0, 
    0.164926714507309, 0.275189074449533, 0, 0, 0.419662898766773, 
    0.349509587043506, 0.332944816429118, 0.350596610318466, 
    0.311231999343016, 0.376799968303961, 0.328697474916696, 
    0.200480163218905, 0.133747295237724, 0.272397704612141, 
    0.464959970657147, 0.510984136394559, 0.500471964320565, 
    0.442803062444463, 0.348294720658541, 0.285097494815857, 
    0.326787718669924, 0.389024358737457, 0.568271614577876, 
    0.748428557676542, 0.673039602589092, 0.702270226528953, 
    0.492109595785327, 0.223787592093243, 0.329205148546915, 
    0.185447956970204, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.170520779257755, 
    0.424952507653855, 0, 1.27581777629185, 1.25745678023744, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.292758057279431, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0.429083083644087, 0.339344945390364, 0.279093453256093, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.392991104409144, 0.509242062064937, 0, 
    0.22447009103248, 0.327959835164993, 0.297835815340399, 0, 
    0.21444874650977, 0.245564512945317, 0.265065412651017, 
    0.283425049160897, 0.282042841931823, 0.272889074043279, 
    0.26301489568171, 0.288852646057119, 0.336921904905559, 
    0.374938166402334, 0.430354578578879, 0.408234545824115, 
    0.345506279547895, 0.229301928058508, 0, 0.818929060434795, 
    0.632955568924026, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.11508567022919, 1.23829440983105, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0.216017746192771, 0.226431946872288, 
    0.195312813900553, 0.208915826340865, 0.258159322024089, 
    0.329889808630425, 0.376411789054799, 0.407353140332676, 
    0.42507368330844, 0.420484932029818, 0.405006425101104, 
    0.384508933765842, 0.370002604887456, 0.344144967422818, 
    0.288732850100452, 0.20339237445048, 0.136718336887777, 
    0.134314370596649, 0.0438642655270794, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.331254511369297, 
    0.390657387257462, 0.412020719092056, 0.375412351310281, 
    0.291519925499765, 0.244155284551186, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.128449526686503, 
    0.251564905129232, 0.184444767724695, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.139393015640656, 0.297685731945459, 0.285501866678608, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;
}
