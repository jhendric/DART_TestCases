netcdf Prior_Diag {
dimensions:
	metadatalength = 64 ;
	locationrank = 1 ;
	copy = 24 ;
	time = UNLIMITED ; // (200 currently)
	NMLlinelen = 129 ;
	NMLnlines = 200 ;
	StateVariable = 1 ;
variables:
	int copy(copy) ;
		copy:long_name = "ensemble member or copy" ;
		copy:units = "nondimensional" ;
		copy:valid_range = 1, 24 ;
	char CopyMetaData(copy, metadatalength) ;
		CopyMetaData:long_name = "Metadata for each copy/member" ;
	char inputnml(NMLnlines, NMLlinelen) ;
		inputnml:long_name = "input.nml contents" ;
	double time(time) ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:cartesian_axis = "T" ;
		time:calendar = "no calendar" ;
		time:units = "days since 0000-00-00 00:00:00" ;
	double loc1d(StateVariable) ;
		loc1d:long_name = "location on unit circle" ;
		loc1d:dimension = 1 ;
		loc1d:units = "nondimensional" ;
		loc1d:valid_range = 0., 1. ;
	int StateVariable(StateVariable) ;
		StateVariable:long_name = "State Variable ID" ;
		StateVariable:units = "indexical" ;
		StateVariable:valid_range = 1, 1 ;
	double state(time, copy, StateVariable) ;
		state:long_name = "model state or fcopy" ;

// global attributes:
		:title = "prior ensemble state" ;
		:assim_model_source = "$URL: https://proxy.subversion.ucar.edu/DAReS/DART/releases/Kodiak/assim_model/assim_model_mod.f90 $" ;
		:assim_model_revision = "$Revision: 4933 $" ;
		:assim_model_revdate = "$Date: 2011-06-01 11:55:44 -0600 (Wed, 01 Jun 2011) $" ;
		:creation_date = "YYYY MM DD HH MM SS = 2012 06 03 13 24 51" ;
		:model_source = "$URL: https://proxy.subversion.ucar.edu/DAReS/DART/releases/Kodiak/models/lorenz_63/model_mod.f90 $" ;
		:model_revision = "$Revision: 4933 $" ;
		:model_revdate = "$Date: 2011-06-01 11:55:44 -0600 (Wed, 01 Jun 2011) $" ;
		:model = "Lorenz_63" ;
		:model_r = 28. ;
		:model_b = 2.6666666666667 ;
		:model_sigma = 10. ;
		:model_deltat = 0.01 ;
data:

 copy = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24 ;

 CopyMetaData =
  "ensemble mean                                                   ",
  "ensemble spread                                                 ",
  "ensemble member      1                                          ",
  "ensemble member      2                                          ",
  "ensemble member      3                                          ",
  "ensemble member      4                                          ",
  "ensemble member      5                                          ",
  "ensemble member      6                                          ",
  "ensemble member      7                                          ",
  "ensemble member      8                                          ",
  "ensemble member      9                                          ",
  "ensemble member     10                                          ",
  "ensemble member     11                                          ",
  "ensemble member     12                                          ",
  "ensemble member     13                                          ",
  "ensemble member     14                                          ",
  "ensemble member     15                                          ",
  "ensemble member     16                                          ",
  "ensemble member     17                                          ",
  "ensemble member     18                                          ",
  "ensemble member     19                                          ",
  "ensemble member     20                                          ",
  "inflation mean                                                  ",
  "inflation sd                                                    " ;

 inputnml =
  "&perfect_model_obs_nml                                                                                                           ",
  "   start_from_restart    = .false.,                                                                                              ",
  "   output_restart        = .true.,                                                                                               ",
  "   async                 = 2,                                                                                                    ",
  "   init_time_days        = 0,                                                                                                    ",
  "   init_time_seconds     = 0,                                                                                                    ",
  "   first_obs_days        = -1,                                                                                                   ",
  "   first_obs_seconds     = -1,                                                                                                   ",
  "   last_obs_days         = -1,                                                                                                   ",
  "   last_obs_seconds      = -1,                                                                                                   ",
  "   output_interval       = 1,                                                                                                    ",
  "   restart_in_file_name  = \"perfect_ics\",                                                                                        ",
  "   restart_out_file_name = \"perfect_restart\",                                                                                    ",
  "   obs_seq_in_file_name  = \"obs_seq.in\",                                                                                         ",
  "   obs_seq_out_file_name = \"obs_seq.out\",                                                                                        ",
  "   adv_ens_command       = \"./advance_model.ksh\",                                                                                ",
  "   output_timestamps     = .false.,                                                                                              ",
  "   trace_execution       = .false.,                                                                                              ",
  "   output_forward_op_errors = .false.,                                                                                           ",
  "   print_every_nth_obs   = -1,                                                                                                   ",
  "   silence               = .false.,                                                                                              ",
  "  /                                                                                                                              ",
  "                                                                                                                                 ",
  "&filter_nml                                                                                                                      ",
  "   async                    = 2,                                                                                                 ",
  "   adv_ens_command          = \"./advance_model.ksh\",                                                                             ",
  "   ens_size                 = 20,                                                                                                ",
  "   start_from_restart       = .false.,                                                                                           ",
  "   output_restart           = .true.,                                                                                            ",
  "   obs_sequence_in_name     = \"obs_seq.out\",                                                                                     ",
  "   obs_sequence_out_name    = \"obs_seq.final\",                                                                                   ",
  "   restart_in_file_name     = \"perfect_ics\",                                                                                     ",
  "   restart_out_file_name    = \"filter_restart\",                                                                                  ",
  "   init_time_days           = 0,                                                                                                 ",
  "   init_time_seconds        = 0,                                                                                                 ",
  "   first_obs_days           = -1,                                                                                                ",
  "   first_obs_seconds        = -1,                                                                                                ",
  "   last_obs_days            = -1,                                                                                                ",
  "   last_obs_seconds         = -1,                                                                                                ",
  "   num_output_state_members = 20,                                                                                                ",
  "   num_output_obs_members   = 0,                                                                                                 ",
  "   output_interval          = 1,                                                                                                 ",
  "   num_groups               = 1,                                                                                                 ",
  "   input_qc_threshold       =  3.0,                                                                                              ",
  "   outlier_threshold        = -1.0,                                                                                              ",
  "   output_forward_op_errors = .false.,                                                                                           ",
  "   output_timestamps        = .false.,                                                                                           ",
  "   output_inflation         = .true.,                                                                                            ",
  "   trace_execution          = .false.,                                                                                           ",
  "   silence                  = .false.,                                                                                           ",
  "                                                                                                                                 ",
  "   inf_flavor                  = 0,                       0,                                                                     ",
  "   inf_initial_from_restart    = .false.,                 .false.,                                                               ",
  "   inf_sd_initial_from_restart = .false.,                 .false.,                                                               ",
  "   inf_output_restart          = .true.,                  .true.,                                                                ",
  "   inf_deterministic           = .true.,                  .true.,                                                                ",
  "   inf_in_file_name            = \'prior_inflate_ics\',     \'post_inflate_ics\',                                                    ",
  "   inf_out_file_name           = \'prior_inflate_restart\', \'post_inflate_restart\',                                                ",
  "   inf_diag_file_name          = \'prior_inflate_diag\',    \'post_inflate_diag\',                                                   ",
  "   inf_initial                 = 1.0,                     1.0,                                                                   ",
  "   inf_sd_initial              = 0.0,                     0.0,                                                                   ",
  "   inf_damping                 = 1.0,                     1.0,                                                                   ",
  "   inf_lower_bound             = 1.0,                     1.0,                                                                   ",
  "   inf_upper_bound             = 1000000.0,               1000000.0,                                                             ",
  "   inf_sd_lower_bound          = 0.0,                     0.0                                                                    ",
  "/                                                                                                                                ",
  "                                                                                                                                 ",
  "&smoother_nml                                                                                                                    ",
  "   num_lags              = 0,                                                                                                    ",
  "   start_from_restart    = .false.,                                                                                              ",
  "   output_restart        = .false.,                                                                                              ",
  "   restart_in_file_name  = \'smoother_ics\',                                                                                       ",
  "   restart_out_file_name = \'smoother_restart\'  /                                                                                 ",
  "                                                                                                                                 ",
  "&ensemble_manager_nml                                                                                                            ",
  "   single_restart_file_in  = .true.,                                                                                             ",
  "   single_restart_file_out = .true.,                                                                                             ",
  "   perturbation_amplitude  = 0.5  /                                                                                              ",
  "                                                                                                                                 ",
  "&assim_tools_nml                                                                                                                 ",
  "   filter_kind                     = 1,                                                                                          ",
  "   cutoff                          = 0.00001,                                                                                    ",
  "   sort_obs_inc                    = .true.,                                                                                     ",
  "   spread_restoration              = .false.,                                                                                    ",
  "   sampling_error_correction       = .false.,                                                                                    ",
  "   adaptive_localization_threshold = -1,                                                                                         ",
  "   output_localization_diagnostics = .false.,                                                                                    ",
  "   localization_diagnostics_file   = \'localization_diagnostics\',                                                                 ",
  "   print_every_nth_obs             = 0  /                                                                                        ",
  "                                                                                                                                 ",
  "&cov_cutoff_nml                                                                                                                  ",
  "   select_localization = 1  /                                                                                                    ",
  "                                                                                                                                 ",
  "&reg_factor_nml                                                                                                                  ",
  "   select_regression    = 1,                                                                                                     ",
  "   input_reg_file       = \"time_mean_reg\",                                                                                       ",
  "   save_reg_diagnostics = .false.,                                                                                               ",
  "   reg_diagnostics_file = \"reg_diagnostics\"  /                                                                                   ",
  "                                                                                                                                 ",
  "&obs_sequence_nml                                                                                                                ",
  "   write_binary_obs_sequence = .false.  /                                                                                        ",
  "                                                                                                                                 ",
  "&obs_kind_nml                                                                                                                    ",
  "   assimilate_these_obs_types = \'RAW_STATE_VARIABLE\'  /                                                                          ",
  "                                                                                                                                 ",
  "&assim_model_nml                                                                                                                 ",
  "   write_binary_restart_files = .false.,                                                                                         ",
  "   netCDF_large_file_support  = .false.                                                                                          ",
  "  /                                                                                                                              ",
  "                                                                                                                                 ",
  "&model_nml                                                                                                                       ",
  "   sigma  = 10.0,                                                                                                                ",
  "   r      = 28.0,                                                                                                                ",
  "   b      = 2.6666666666667,                                                                                                     ",
  "   deltat = 0.01,                                                                                                                ",
  "   time_step_days = 1,                                                                                                           ",
  "   time_step_seconds = 0  /                                                                                                      ",
  "                                                                                                                                 ",
  "&utilities_nml                                                                                                                   ",
  "   TERMLEVEL = 1,                                                                                                                ",
  "   module_details = .false.,                                                                                                     ",
  "   logfilename = \'dart_log.out\',                                                                                                 ",
  "   nmlfilename = \'dart_log.nml\',                                                                                                 ",
  "   write_nml   = \'terminal\'  /                                                                                                   ",
  "                                                                                                                                 ",
  "&preprocess_nml                                                                                                                  ",
  "    input_obs_def_mod_file = \'../../../obs_def/DEFAULT_obs_def_mod.F90\',                                                         ",
  "   output_obs_def_mod_file = \'../../../obs_def/obs_def_mod.f90\',                                                                 ",
  "   input_obs_kind_mod_file = \'../../../obs_kind/DEFAULT_obs_kind_mod.F90\',                                                       ",
  "  output_obs_kind_mod_file = \'../../../obs_kind/obs_kind_mod.f90\',                                                               ",
  "               input_files = \'../../../obs_def/obs_def_1d_state_mod.f90\'  /                                                      ",
  "                                                                                                                                 ",
  "                                                                                                                                 ",
  "&obs_sequence_tool_nml                                                                                                           ",
  "   num_input_files   = 2,                                                                                                        ",
  "   filename_seq      = \'obs_seq.one\', \'obs_seq.two\',                                                                             ",
  "   filename_out      = \'obs_seq.processed\',                                                                                      ",
  "   first_obs_days    = -1,                                                                                                       ",
  "   first_obs_seconds = -1,                                                                                                       ",
  "   last_obs_days     = -1,                                                                                                       ",
  "   last_obs_seconds  = -1,                                                                                                       ",
  "   print_only        = .false.,                                                                                                  ",
  "   gregorian_cal     = .false.                                                                                                   ",
  "   /                                                                                                                             ",
  "                                                                                                                                 ",
  "# other possible obs tool namelist items:                                                                                        ",
  "#                                                                                                                                ",
  "# keep only the U and V radiosonde winds:                                                                                        ",
  "#   obs_types          = \'RADIOSONDE_U_WIND_COMPONENT\',                                                                          ",
  "#                        \'RADIOSONDE_V_WIND_COMPONENT\',                                                                          ",
  "#   keep_types         = .true.,                                                                                                 ",
  "#                                                                                                                                ",
  "# remove the U and V radiosonde winds:                                                                                           ",
  "#   obs_types          = \'RADIOSONDE_U_WIND_COMPONENT\',                                                                          ",
  "#                        \'RADIOSONDE_V_WIND_COMPONENT\',                                                                          ",
  "#   keep_types         = .false.,                                                                                                ",
  "#                                                                                                                                ",
  "# keep only observations with a DART QC of 0:                                                                                    ",
  "#   qc_metadata        = \'Dart quality control\',                                                                                 ",
  "#   min_qc             = 0,                                                                                                      ",
  "#   max_qc             = 0,                                                                                                      ",
  "#                                                                                                                                ",
  "# keep only radiosonde temp obs between 250 and 300 K:                                                                           ",
  "#   copy_metadata      = \'NCEP BUFR observation\',                                                                                ",
  "#   copy_type          = \'RADIOSONDE_TEMPERATURE\',                                                                               ",
  "#   min_copy           = 250.0,                                                                                                  ",
  "#   max_copy           = 300.0,                                                                                                  ",
  "#                                                                                                                                ",
  "                                                                                                                                 ",
  "                                                                                                                                 ",
  "&restart_file_tool_nml                                                                                                           ",
  "   input_file_name              = \"filter_restart\",                                                                              ",
  "   output_file_name             = \"filter_updated_restart\",                                                                      ",
  "   ens_size                     = 1,                                                                                             ",
  "   single_restart_file_in       = .true.,                                                                                        ",
  "   single_restart_file_out      = .true.,                                                                                        ",
  "   write_binary_restart_files   = .true.,                                                                                        ",
  "   overwrite_data_time          = .false.,                                                                                       ",
  "   new_data_days                = -1,                                                                                            ",
  "   new_data_secs                = -1,                                                                                            ",
  "   input_is_model_advance_file  = .false.,                                                                                       ",
  "   output_is_model_advance_file = .false.,                                                                                       ",
  "   overwrite_advance_time       = .false.,                                                                                       ",
  "   new_advance_days             = -1,                                                                                            ",
  "   new_advance_secs             = -1,                                                                                            ",
  "   gregorian_cal                = .false.                                                                                        ",
  "/                                                                                                                                ",
  "                                                                                                                                 ",
  "&obs_diag_nml                                                                                                                    ",
  "   obs_sequence_name  = \'obs_seq.final\',                                                                                         ",
  "   iskip_days         = 0,                                                                                                       ",
  "   obs_select         = 1,                                                                                                       ",
  "   rat_cri            = 4.0,                                                                                                     ",
  "   input_qc_threshold = 3.0,                                                                                                     ",
  "   bin_width_seconds = 0,                                                                                                        ",
  "   lonlim1   = 0.0, 0.0, 0.5, -1.0,                                                                                              ",
  "   lonlim2   = 1.0, 0.5, 1.5, -1.0,                                                                                              ",
  "   reg_names = \'whole\', \'yin\', \'yang\', \'bogus\',                                                                                  ",
  "   verbose   = .false.  /                                                                                                        ",
  "                                                                                                                                 " ;

 time = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 107, 
    108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 121, 
    122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 
    136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 149, 
    150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 
    164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 177, 
    178, 179, 180, 181, 182, 183, 184, 185, 186, 187, 188, 189, 190, 191, 
    192, 193, 194, 195, 196, 197, 198, 199, 200 ;

 loc1d = 0 ;

 StateVariable = 1 ;

 state =
  -77.6189152312488,
  0.666047915162125,
  -77.4585064213575,
  -76.7576060387359,
  -77.4880621233776,
  -76.7505481814382,
  -77.7316000257459,
  -78.9969022200512,
  -77.2351712352554,
  -78.3484475797791,
  -78.2958662859241,
  -78.735890591093,
  -77.230686978927,
  -78.5094263122399,
  -77.2104149260008,
  -77.138096722939,
  -77.8821150492247,
  -76.7551824973405,
  -77.7707522457994,
  -77.7356831820767,
  -77.1361249340919,
  -77.2112210735788,
  1,
  0,
  -77.3992408266583,
  0.506194907598424,
  -76.3189409995828,
  -77.5165131342934,
  -77.4268059478982,
  -77.1757862777486,
  -77.4960213185389,
  -78.1968947500926,
  -76.4641334921074,
  -77.7079172617253,
  -77.8447743967774,
  -77.3551282136969,
  -76.7080739464373,
  -77.4008299026983,
  -76.953759405301,
  -77.8439787261039,
  -77.9564498968702,
  -77.3309203206906,
  -77.5484860071628,
  -78.0472703966525,
  -77.0425960950891,
  -77.649536043699,
  1,
  0,
  -77.2703781388403,
  0.433258248258373,
  -76.4534890294724,
  -77.1229213785662,
  -77.3832335877069,
  -76.8108970329186,
  -76.8180172739769,
  -77.8105263985068,
  -77.5898406545314,
  -77.6457135798066,
  -77.6133120743764,
  -77.2986249451487,
  -77.1468111291291,
  -76.6515737865644,
  -76.6778925912132,
  -77.168045246843,
  -77.7420855098606,
  -76.9648928802149,
  -77.8169138719305,
  -77.6429779060899,
  -77.2480518036697,
  -77.80174209628,
  1,
  0,
  -77.3841881844721,
  0.36092913950603,
  -77.2271184438795,
  -77.5878756648131,
  -77.3815628385976,
  -76.5170074474666,
  -77.5063929197261,
  -77.302926460238,
  -77.3964270992056,
  -77.4899408275444,
  -77.5890626193765,
  -77.3606048440699,
  -77.1853893871713,
  -77.4898393544794,
  -76.7650947616963,
  -77.3747895552252,
  -77.5542084639818,
  -77.0967379663306,
  -78.2823637705463,
  -77.2425826999987,
  -77.8239697995244,
  -77.5098687655708,
  1,
  0,
  -77.4443274250274,
  0.463819390483465,
  -77.9722363785519,
  -77.3764127081813,
  -77.5394554751889,
  -76.8966816631522,
  -77.3191123652557,
  -77.1718670196304,
  -77.7699270682322,
  -77.7128490634769,
  -77.3650606319282,
  -77.7784817290994,
  -76.42827003158,
  -77.970068837569,
  -76.5572291241804,
  -77.5259772070678,
  -77.7544615750702,
  -77.5571435579052,
  -77.4578272005339,
  -76.9217194865089,
  -78.2209493374863,
  -77.5908180399486,
  1,
  0,
  -77.9777104988079,
  0.573914697763237,
  -78.3980569986509,
  -77.4772890847471,
  -78.758778718306,
  -77.631584696803,
  -77.0172879116042,
  -77.6791931801825,
  -78.7403864433618,
  -77.9118273278435,
  -77.851975206939,
  -78.0717965197659,
  -77.2038532511733,
  -79.1056832011045,
  -77.4447983396387,
  -77.6303121004516,
  -78.4832342903285,
  -77.9315042905477,
  -78.2487913496777,
  -77.4023952193278,
  -78.7039814690137,
  -77.8614803766914,
  1,
  0,
  -78.8002374466779,
  0.499667906776583,
  -78.6068810671351,
  -78.2800427172867,
  -79.4574201615932,
  -77.7635052419697,
  -78.5069358691743,
  -78.6823834476535,
  -79.2582431424471,
  -79.0695522552677,
  -79.2593976545235,
  -79.2428671659604,
  -78.3013781384662,
  -78.8918170101442,
  -78.0203138091022,
  -78.6886079698281,
  -79.784116739782,
  -78.5504427978893,
  -79.2695409480325,
  -78.7051101873743,
  -78.8424879768872,
  -78.8237046330408,
  1,
  0,
  -79.5640429023263,
  0.501724916913907,
  -79.1631059683339,
  -79.1350694943588,
  -79.2366776124558,
  -78.592923490037,
  -79.7961987430433,
  -78.9891306394673,
  -80.4087888578143,
  -79.984728422821,
  -79.8495129172091,
  -79.4180970433825,
  -79.3801601415357,
  -80.2959773503184,
  -79.6698192772234,
  -80.2595329498415,
  -79.9610753218222,
  -78.8480831969312,
  -79.8656604422387,
  -79.800838995227,
  -79.3444588854026,
  -79.2810182970627,
  1,
  0,
  -80.2545404925377,
  0.558274618011392,
  -79.5951039309723,
  -80.1211277097826,
  -79.9153550613993,
  -79.4374194038114,
  -81.0429657437832,
  -79.5036113145687,
  -80.2532412023902,
  -81.1374210633037,
  -80.5892048274861,
  -80.3081568933648,
  -80.2217382455084,
  -81.4905229032375,
  -80.5539438499341,
  -80.0768261803062,
  -80.833478489667,
  -79.8624007647878,
  -80.0121482922973,
  -80.4723279196616,
  -79.7862475840882,
  -79.8775684704035,
  1,
  0,
  -81.3753105571,
  0.473370577257571,
  -80.6532084004444,
  -81.6566740331885,
  -81.0195955986853,
  -80.6750578958245,
  -82.3064915767151,
  -81.4762799886358,
  -80.8027498085527,
  -81.6155882913801,
  -80.6540418257311,
  -81.29343317099,
  -81.7180512511273,
  -82.3125602514717,
  -81.1874020185687,
  -81.3867674441502,
  -81.4140460915126,
  -81.1569387650522,
  -81.6136799146057,
  -81.7017790774233,
  -81.4387060450661,
  -81.4231596928739,
  1,
  0,
  -82.2591104553939,
  0.371640699275297,
  -82.0203867329333,
  -82.5072643105352,
  -82.1468850711452,
  -81.712044908201,
  -83.2084590864401,
  -82.4971153810055,
  -81.9327729371186,
  -82.0558165985949,
  -82.1382526309745,
  -82.0313317842038,
  -82.524572192046,
  -82.2290656643477,
  -82.1994425069539,
  -81.8653987872792,
  -82.5035194394394,
  -81.7924451778913,
  -82.235023097541,
  -82.8958409148796,
  -82.1265829182793,
  -82.559988968069,
  1,
  0,
  -83.1409945530114,
  0.475231883781707,
  -82.4850005619332,
  -83.0726767069081,
  -83.5622378324952,
  -82.9001618793533,
  -83.7924358244353,
  -83.9548385688042,
  -82.8981402165904,
  -82.9608939176189,
  -83.2639009634682,
  -82.4636543756046,
  -83.511329005332,
  -82.5726324775691,
  -82.7882660853964,
  -82.7327751761545,
  -83.6522833472557,
  -82.5547823905531,
  -83.6201655119315,
  -83.7059942672489,
  -83.340513419712,
  -82.987208531864,
  1,
  0,
  -84.0871810179779,
  0.542828858587319,
  -83.1178000602093,
  -84.4752051803494,
  -84.9518260892261,
  -84.5050235344907,
  -84.3045221559915,
  -84.1209739549681,
  -83.5377810810712,
  -83.5374769946613,
  -84.7298604089558,
  -84.0296742827266,
  -84.6210241081844,
  -83.7447262981516,
  -83.9776319203392,
  -83.822691846143,
  -84.6533115463362,
  -82.9914598996257,
  -84.4137392855873,
  -84.3184089152372,
  -83.5504828021799,
  -84.3399999951234,
  1,
  0,
  -85.2533483279611,
  0.687657367561377,
  -84.880233530103,
  -85.5520270419974,
  -86.4210182633777,
  -85.8671474923888,
  -85.5035835775829,
  -84.7554980204925,
  -85.2153957487131,
  -84.9276356236817,
  -85.8769280289079,
  -85.1615908074152,
  -86.2139723967906,
  -83.9737896099853,
  -83.9252898822736,
  -85.5111408315492,
  -85.6225917521276,
  -84.1717024811439,
  -84.804406295959,
  -85.6692520187581,
  -85.4841367344175,
  -85.5296264215574,
  1,
  0,
  -86.9784495923134,
  0.523818506604831,
  -85.8112403280483,
  -87.1732277010759,
  -87.0487207909414,
  -86.7671986372013,
  -87.1515532465711,
  -86.8726160022202,
  -86.9576911115363,
  -87.505653885536,
  -87.1127969691986,
  -87.0221300975699,
  -87.4448650262481,
  -85.9803855721408,
  -86.2256683413576,
  -87.7078929055847,
  -87.1179011383076,
  -86.8165490834066,
  -87.1554820077951,
  -87.8674461538295,
  -87.258599804971,
  -86.5713730427287,
  1,
  0,
  -88.1060676598403,
  0.399588187187834,
  -87.3251723120826,
  -88.1679437505144,
  -88.2184732778075,
  -87.3863432946138,
  -88.4293346760982,
  -88.1005043538937,
  -88.8531249873693,
  -88.8482459686235,
  -88.2432576860612,
  -88.0669316796079,
  -87.8097584996233,
  -88.0052312251536,
  -87.8732866117571,
  -88.3695695940345,
  -88.1841452688496,
  -87.7877144281064,
  -88.1372313944191,
  -88.1440641314859,
  -88.4876159387324,
  -87.6834041179729,
  1,
  0,
  -88.8293142155,
  0.651159249256713,
  -88.5439088811795,
  -88.7916537588204,
  -88.9670058410184,
  -88.1660646117404,
  -89.0674146147306,
  -88.1918847558075,
  -89.9199748459445,
  -90.2308539877561,
  -89.1655900144374,
  -88.9284177609882,
  -87.6244347746774,
  -89.3566975742759,
  -87.8580325572911,
  -88.9142117952164,
  -88.8268272522927,
  -87.8986668185085,
  -88.8950699176318,
  -88.9308888444966,
  -89.18718738877,
  -89.1214983144173,
  1,
  0,
  -89.8069607157603,
  0.860049070512546,
  -89.2580213991174,
  -89.3728000401597,
  -90.3526509507843,
  -89.8560848089384,
  -89.6461495638105,
  -89.5273031720936,
  -91.2470843077961,
  -90.9772752372062,
  -89.9166321101222,
  -90.2306476020883,
  -89.0805372571906,
  -90.9769708190752,
  -89.333438760456,
  -89.0294129508114,
  -88.1980196430548,
  -88.0535015857301,
  -90.1253291457524,
  -90.1776207486144,
  -90.0599063434301,
  -90.7198278689737,
  1,
  0,
  -91.3569670714115,
  0.697919483985262,
  -90.7934401007527,
  -91.0850779656974,
  -91.1392540369834,
  -91.3467577037002,
  -91.0413064498042,
  -91.7670441501874,
  -92.7821160267282,
  -92.2165436849789,
  -91.7648881963747,
  -91.2955806093904,
  -90.3478123269824,
  -92.27343225955,
  -91.3347535871459,
  -90.9775284718901,
  -89.8401409432788,
  -90.4810849261817,
  -91.4965438550896,
  -92.0013956217351,
  -91.628681507603,
  -91.525959004175,
  1,
  0,
  -91.9551726926394,
  0.491761561401882,
  -91.6003920317796,
  -92.3272300655809,
  -92.3749570737915,
  -92.1267308535555,
  -91.5150303442823,
  -92.2259871352442,
  -92.929527207983,
  -92.2314153066144,
  -91.7774373156096,
  -91.4579708677895,
  -91.3655673642265,
  -93.0840521425626,
  -91.2709504377637,
  -91.6227616784294,
  -92.2881079404254,
  -91.570991042841,
  -91.9090456646996,
  -91.7798282051015,
  -91.7082460500439,
  -91.9372251244643,
  1,
  0,
  -92.6290998958044,
  0.693128353400419,
  -92.8481353059317,
  -92.5730374997765,
  -92.9625899204768,
  -92.9645237812717,
  -92.489902610133,
  -93.4470905038236,
  -93.6979785385667,
  -93.0222594362273,
  -90.9530903800244,
  -91.8260930773958,
  -92.5678455052473,
  -93.9630872214345,
  -92.6923712464828,
  -92.3960150410319,
  -92.5777317696948,
  -92.8245094831771,
  -92.255520152689,
  -91.5029727786234,
  -92.291027003251,
  -92.7262166608298,
  1,
  0,
  -92.9347900528285,
  0.683048374437113,
  -93.5348820763102,
  -92.2147502483911,
  -93.2927379070913,
  -93.2716387395889,
  -92.7231444038547,
  -93.8975397721491,
  -93.8010899927179,
  -93.5279954892016,
  -92.4832231660589,
  -92.4486758907684,
  -92.1885433578317,
  -94.5084429392976,
  -93.0454994727913,
  -92.2943547204282,
  -92.8588328469788,
  -92.5974008192135,
  -92.311812911062,
  -92.3233975449943,
  -92.0658148628925,
  -93.3060238949481,
  1,
  0,
  -93.116686129408,
  0.7537347705587,
  -93.9123531924441,
  -92.8719725989857,
  -93.5260321510044,
  -93.4282076642761,
  -93.3819694616456,
  -93.559174745958,
  -94.8876639267662,
  -93.4599757819409,
  -92.7639500349022,
  -92.6271287972002,
  -91.8610489267443,
  -94.3493581166247,
  -92.438150046534,
  -92.2381110480412,
  -93.3453015162641,
  -93.0052236579677,
  -92.401370049457,
  -92.6989902057565,
  -92.2152929572933,
  -93.3624477083534,
  1,
  0,
  -92.8453731263038,
  0.63000662186678,
  -93.7695774807479,
  -92.4503942444746,
  -93.0984254747773,
  -93.2449603151748,
  -92.8876445989012,
  -92.5971509941892,
  -93.8353940987824,
  -92.5948966392344,
  -92.9408252429895,
  -92.7226050308503,
  -91.6258063831096,
  -93.2645046938594,
  -92.5684900083367,
  -92.0271477584948,
  -94.0668633640171,
  -92.6239261083993,
  -91.7681130340056,
  -93.0992390879774,
  -92.8355664287174,
  -92.8859315390365,
  1,
  0,
  -93.3763339360516,
  0.58670504258519,
  -94.3197951073479,
  -92.6595603117114,
  -93.4726219427029,
  -93.6411095932484,
  -93.7537439751693,
  -92.8564704410153,
  -93.7274354616877,
  -93.0022826256188,
  -93.4157733527869,
  -93.1043078936962,
  -92.0589426168081,
  -93.5750581290157,
  -93.2359591661251,
  -92.8856192892074,
  -94.4962727765927,
  -93.2433626829177,
  -93.1924628452613,
  -94.0694654925914,
  -93.8990337431185,
  -92.9174012744084,
  1,
  0,
  -93.7529961206516,
  0.607802817967594,
  -94.9416547842693,
  -93.3668122138519,
  -93.9209042264616,
  -94.1837431056871,
  -93.7332312146048,
  -92.9964694059263,
  -94.8044800836203,
  -93.2273927977814,
  -93.7430493204653,
  -93.3754331223747,
  -93.5209626413596,
  -94.1553425069386,
  -92.933060140394,
  -93.2031851697499,
  -94.0803048470084,
  -93.9619524642317,
  -93.9090810414908,
  -94.4561388559903,
  -93.9160330407549,
  -92.6306914300721,
  1,
  0,
  -93.744279666132,
  0.794893642458335,
  -94.7069409851749,
  -93.3823679364027,
  -93.8836122576754,
  -94.7507697918381,
  -93.7047874839112,
  -92.2788025312492,
  -94.8045872635392,
  -93.8115980642327,
  -93.6506177752341,
  -92.6529428556556,
  -93.932751967727,
  -94.1323298599335,
  -93.6460899335284,
  -93.3867880540322,
  -94.1199604036187,
  -94.7882093604472,
  -94.0738188137747,
  -93.7729712305133,
  -93.5984295284087,
  -91.8072172257431,
  1,
  0,
  -92.8867394660165,
  0.920926763192229,
  -94.2542186908145,
  -92.6069562428852,
  -93.3620830896502,
  -94.1301070817052,
  -92.7237874528853,
  -91.1232448957518,
  -94.0140079579715,
  -92.1677665578626,
  -93.2324758243209,
  -92.0549331385398,
  -93.6582499272492,
  -93.4529849781907,
  -92.1034070710932,
  -92.5611634835901,
  -92.846096947061,
  -93.9031871227092,
  -92.84710774445,
  -93.4025313281073,
  -92.2099174355646,
  -91.0805623499273,
  1,
  0,
  -92.6915529097237,
  0.899133228654806,
  -94.2362966866125,
  -92.5475751695879,
  -93.0965354438421,
  -93.7925079876559,
  -92.3367620240893,
  -91.4645417126898,
  -93.5296519100853,
  -91.9429224098676,
  -93.700909534899,
  -92.1702508450616,
  -93.3326655535905,
  -92.0965604448367,
  -92.3109017102235,
  -92.8005678987498,
  -92.571652602264,
  -94.0550028454435,
  -91.5638750401356,
  -92.945470270207,
  -92.4319571346358,
  -90.9044509699955,
  1,
  0,
  -91.8277615118665,
  1.07135655363357,
  -94.0605322830064,
  -92.2909900728975,
  -91.6242312664493,
  -93.0254415250658,
  -92.1303467854232,
  -91.2691696326641,
  -93.5397533252064,
  -91.47963052236,
  -91.6680664740021,
  -90.3680605884311,
  -91.8715153764865,
  -90.7637683903069,
  -92.2207126169139,
  -92.1356197168508,
  -91.6831457333458,
  -92.5891127257832,
  -90.6954402263602,
  -92.2708021999215,
  -91.4774728738451,
  -89.3914179020112,
  1,
  0,
  -91.6196202886103,
  0.877948498762702,
  -93.4951562754624,
  -92.0468514597223,
  -91.7885256065357,
  -92.0445071408255,
  -91.5280328577032,
  -92.3071641393696,
  -92.5035342524331,
  -91.0895562714696,
  -91.0033282044967,
  -90.6892933128589,
  -91.5279635418912,
  -90.6311076967544,
  -92.3920394835332,
  -91.4305697569985,
  -91.101325466723,
  -92.5198265891011,
  -90.8494916067037,
  -92.1990359909131,
  -91.7026175252488,
  -89.5424785934634,
  1,
  0,
  -91.8106796772517,
  0.976771522516385,
  -94.2431496963617,
  -92.6774935754122,
  -91.9478222192199,
  -91.7425272034866,
  -91.7162534988246,
  -92.2958999658171,
  -92.324649220062,
  -91.5500997437675,
  -91.11603503647,
  -90.4773731114646,
  -91.6256209751507,
  -90.9201001052416,
  -92.1488064384116,
  -91.7585505330169,
  -91.4897285183606,
  -93.10284964589,
  -90.6941267012637,
  -92.3286041940941,
  -92.2796778557298,
  -89.774225306989,
  1,
  0,
  -91.2655032872001,
  1.04641990485182,
  -93.4132837339008,
  -91.8267348675842,
  -92.1763123637435,
  -91.3950572024754,
  -91.7615292406752,
  -91.5218669049431,
  -91.6584188190914,
  -91.4930930637036,
  -90.7381574986946,
  -89.8417007571767,
  -90.5130903245617,
  -90.3187457536784,
  -90.9386141753659,
  -91.0090105272321,
  -91.0922300694848,
  -93.098741382501,
  -90.7281674818728,
  -91.8981350810541,
  -91.1678370927547,
  -88.7193394035079,
  1,
  0,
  -91.0780471925111,
  1.20762050690714,
  -93.425362026723,
  -91.6921019817106,
  -91.9018306888762,
  -91.0950299356004,
  -91.4071208637129,
  -91.4707792380899,
  -91.710536886128,
  -91.1172869414755,
  -90.139753585286,
  -88.7752772596747,
  -90.315325510619,
  -90.2601418396223,
  -91.0480437830047,
  -90.7873931012589,
  -91.0891128481608,
  -93.0554278198288,
  -90.5863044760459,
  -91.8663609663493,
  -91.5599476344441,
  -88.2578064636107,
  1,
  0,
  -91.312734405492,
  1.17878691116363,
  -93.5520573223861,
  -92.226741090735,
  -92.221110821744,
  -91.8466303849731,
  -91.5490223898966,
  -91.53599805631,
  -91.3266883905393,
  -91.2118836425733,
  -90.0029108165991,
  -89.4670763369737,
  -90.5739800877651,
  -89.8076080878989,
  -90.9504664759275,
  -91.0286185964198,
  -91.6812412511036,
  -93.3295273228677,
  -90.7183525779349,
  -92.7436794243484,
  -91.307433742658,
  -89.1736612901854,
  1,
  0,
  -91.2713016989742,
  1.30707820892912,
  -93.7630427510047,
  -91.6173228315901,
  -91.9869899274752,
  -91.4865555770867,
  -91.369153890082,
  -91.5884521406035,
  -91.878946551048,
  -91.2853348464485,
  -90.0691091175016,
  -88.9417722671155,
  -90.5650741580027,
  -90.1024770338653,
  -91.2472259176218,
  -90.6482954097919,
  -92.0199045245937,
  -93.7026746970396,
  -90.3287465168363,
  -92.7175655649316,
  -91.3862073650805,
  -88.7211828917642,
  1,
  0,
  -91.4458355313091,
  1.38344631524294,
  -94.2623238883462,
  -92.6700789492493,
  -92.2073008955248,
  -90.7695967006836,
  -91.4179556199476,
  -92.7443196173367,
  -92.4738703211722,
  -91.3946583522986,
  -90.2491806234926,
  -90.0706456804447,
  -90.6367010803214,
  -89.3976544158147,
  -90.4576657437233,
  -91.4087237876068,
  -91.8279142857507,
  -93.8828113918865,
  -89.7283127976087,
  -92.3098017259682,
  -91.6086349853219,
  -89.3985597636837,
  1,
  0,
  -90.8185223349499,
  1.31169390060263,
  -93.9975448345531,
  -91.8828001907244,
  -91.5636913495428,
  -90.1710302660309,
  -90.0436849410643,
  -91.488107105187,
  -91.1323845256169,
  -91.2730739870587,
  -90.2002234421467,
  -90.7033371468724,
  -90.3472841697621,
  -88.7027393538363,
  -89.4762454610199,
  -91.5536199983838,
  -90.6723896114444,
  -92.4978074649458,
  -89.1162945490406,
  -92.2349101393664,
  -90.4446005939499,
  -88.868677568452,
  1,
  0,
  -90.5974179961216,
  1.32479066172705,
  -93.2107879172392,
  -91.3840673409154,
  -91.4368635203967,
  -90.7496676744093,
  -88.914224685674,
  -91.617332259955,
  -91.3963015987545,
  -91.2225649884732,
  -89.0803302107084,
  -90.5970683393789,
  -90.4215975869993,
  -88.3965255301824,
  -90.1008866693117,
  -91.3514194381124,
  -89.9712792226777,
  -92.3220915581711,
  -88.7907952262478,
  -92.1436540546262,
  -89.9125579854666,
  -88.9283441147332,
  1,
  0,
  -90.4625398375769,
  1.26278241070999,
  -93.3257219586904,
  -91.112736578558,
  -92.181517394993,
  -89.9542212349763,
  -89.220843424589,
  -91.2294768885198,
  -90.555484088947,
  -91.0904386439717,
  -88.7009382121997,
  -89.7912404498225,
  -90.556289388558,
  -88.2943715693403,
  -90.1513945216144,
  -90.6065674810715,
  -90.1471104648057,
  -92.160149620041,
  -89.6049790798049,
  -91.5998527495702,
  -90.0420563203975,
  -88.925406681068,
  1,
  0,
  -90.1958534632904,
  1.16683906367918,
  -92.1379586282069,
  -90.2286428807892,
  -91.8211006593432,
  -88.9964924791211,
  -89.0502088241231,
  -90.7498458446117,
  -90.1779718104057,
  -91.5103864465784,
  -89.0481501120183,
  -89.800067204932,
  -90.1017389576351,
  -88.4698703954244,
  -89.851229278841,
  -89.9023417163914,
  -90.9170288296694,
  -92.5902504908629,
  -90.0141604028953,
  -90.6640603364353,
  -89.3645572226057,
  -88.5210067449186,
  1,
  0,
  -89.5663524494916,
  0.992932251084082,
  -91.1280669237339,
  -88.951929807008,
  -91.51101562632,
  -88.9530298171391,
  -88.1624036902243,
  -90.161863404072,
  -89.4215831106856,
  -90.7626526725977,
  -89.53336044588,
  -89.3519730315182,
  -88.8709093325916,
  -88.8026158833165,
  -88.8644121320796,
  -89.5494373694581,
  -89.3816118439211,
  -91.427491477507,
  -88.8437511619954,
  -90.2805347360246,
  -89.0628133021998,
  -88.30559322156,
  1,
  0,
  -88.1273764001533,
  0.894925999700991,
  -88.9796057403501,
  -88.0650144620808,
  -90.4330553286265,
  -88.3047991260242,
  -86.4957038436695,
  -88.6818002137454,
  -88.7460474980769,
  -88.4610165923595,
  -88.3167147093518,
  -87.394740418938,
  -87.4324956021158,
  -87.7405240615797,
  -86.8766029678963,
  -87.4892943070321,
  -87.6643858968659,
  -89.3103525340157,
  -87.8713175902086,
  -88.829644715212,
  -87.6732800568624,
  -87.7811323380557,
  1,
  0,
  -87.1496276393718,
  1.00311852807226,
  -87.3052987816442,
  -86.6901542184734,
  -89.5786287626229,
  -86.7236011623888,
  -84.9665505054611,
  -87.2202455859293,
  -87.21400144771,
  -86.612723928921,
  -88.0983062138863,
  -86.5382892258808,
  -86.1984327712091,
  -86.8806898476024,
  -86.7346246782589,
  -86.9291564117746,
  -86.3374131502315,
  -88.6947468679544,
  -86.8438310573392,
  -88.466409156378,
  -87.7750832058092,
  -87.184365807962,
  1,
  0,
  -86.9148547367532,
  0.859766266190581,
  -86.7121504303196,
  -86.4446242798788,
  -88.4319402591018,
  -86.7773057498745,
  -84.892000629432,
  -87.3020855043236,
  -87.0415487489604,
  -86.1195476772099,
  -87.3599984831369,
  -86.4832686456059,
  -85.9177892798241,
  -87.0141145596703,
  -86.317526251429,
  -86.4105903639684,
  -86.3992193851096,
  -88.3209119024376,
  -87.0503636089279,
  -88.0463511788014,
  -87.7109807575271,
  -87.5447770395249,
  1,
  0,
  -85.0987436898058,
  0.844451405960837,
  -85.1953457882863,
  -84.6762882563803,
  -87.1546357428856,
  -84.7575295031354,
  -83.4648506485035,
  -85.0915936843048,
  -85.2618814687852,
  -85.2767356362142,
  -85.2807389279976,
  -84.6897374592326,
  -83.7775105650659,
  -84.260558717608,
  -85.1789806267281,
  -84.9651038341542,
  -84.0566915396883,
  -85.5920260848757,
  -85.6472874332282,
  -86.1200580450835,
  -85.9363812199547,
  -85.5909386140044,
  1,
  0,
  -83.4831468525212,
  0.691929892568083,
  -83.7791687289265,
  -82.9595593567976,
  -84.9784510312074,
  -83.3405965119999,
  -82.4251938316404,
  -83.7464929716608,
  -83.8748368555759,
  -83.7129929843011,
  -83.2927559863241,
  -82.8463337858094,
  -82.5642468594699,
  -82.8372586305676,
  -82.8288358722486,
  -83.6021957897758,
  -82.6494203994682,
  -83.8432622480245,
  -84.133130237523,
  -84.7177379231423,
  -83.8261942328179,
  -83.7042728131421,
  1,
  0,
  -83.1216444021642,
  0.748519715510838,
  -82.6087425720454,
  -82.3091806681534,
  -84.4914464014531,
  -83.8120974895799,
  -81.913017208044,
  -83.4413199035987,
  -83.4418634429357,
  -83.3592711186502,
  -83.2371357180193,
  -82.4806880915235,
  -82.3611061608621,
  -82.3145586488088,
  -82.2495533932717,
  -83.1811625311737,
  -82.4276416204431,
  -83.5483801341995,
  -83.4926495942872,
  -84.4765391401054,
  -83.7978044608445,
  -83.488729745284,
  1,
  0,
  -82.4283310533793,
  0.731299611278349,
  -82.2437396751496,
  -81.8086145166429,
  -83.14706781813,
  -82.6777630000613,
  -81.7610625625386,
  -82.6346679209503,
  -82.9065675902004,
  -82.3251832405607,
  -82.3989032607822,
  -81.7385493374237,
  -81.2507684644544,
  -81.4734002685193,
  -81.3057963795267,
  -83.05215546745,
  -82.050379347531,
  -83.1262574980962,
  -82.962855516421,
  -84.0908200666523,
  -82.9606033705945,
  -82.6514657659013,
  1,
  0,
  -82.468783245315,
  0.661313354115407,
  -81.5906118347061,
  -81.83021916725,
  -83.2386403515042,
  -82.7182883987111,
  -81.4241399386541,
  -82.9148252587064,
  -82.9861904126776,
  -82.087059132444,
  -83.1587922855765,
  -82.0576471259061,
  -81.3975804931255,
  -81.9142660134094,
  -81.7077479012529,
  -83.4563008905441,
  -82.8492764043751,
  -82.3952464050092,
  -82.6542242338978,
  -83.2232957509107,
  -82.7964082112359,
  -82.9749046964039,
  1,
  0,
  -82.7409149201698,
  0.556784384361563,
  -82.100916539941,
  -81.9568932688989,
  -83.3200416105137,
  -82.5023986731039,
  -81.7377623012998,
  -82.8740469451979,
  -82.9399932995053,
  -82.7812868443298,
  -83.6402814477991,
  -83.0056539375058,
  -82.080073222411,
  -82.4001222532021,
  -81.8299738395547,
  -82.9209396750118,
  -83.2198629503601,
  -82.9265121219951,
  -82.8483175729857,
  -83.0948747446289,
  -83.4689295930318,
  -83.1694175621195,
  1,
  0,
  -82.3563147778179,
  0.626382692708521,
  -81.628766788748,
  -81.519072862156,
  -82.7758779425082,
  -82.0490063700826,
  -81.0283724008222,
  -82.3905360056057,
  -82.1654994468179,
  -82.3986251948026,
  -83.3823113676352,
  -82.4815949450875,
  -82.3496219511647,
  -81.926627144159,
  -81.5075269241157,
  -82.8666556625367,
  -83.187566162547,
  -82.3550297428686,
  -82.6618336500659,
  -82.658262014256,
  -82.4184229404777,
  -83.3750860398998,
  1,
  0,
  -83.3353359778999,
  0.653387164363982,
  -82.3750113428022,
  -82.6509693456669,
  -84.6654602947359,
  -83.0247732102926,
  -82.4354568337614,
  -83.1350846059824,
  -83.5652887334624,
  -83.7622564937417,
  -84.0784223340828,
  -83.6941085801193,
  -83.1152432186446,
  -83.9324848479191,
  -82.2770592611986,
  -82.3840828141712,
  -83.9586443251329,
  -83.3853691760733,
  -83.5283736483679,
  -83.5702713704772,
  -83.4229010982169,
  -83.7454580231494,
  1,
  0,
  -83.8990619299493,
  0.770034791369627,
  -83.3556786254864,
  -83.0944558689956,
  -84.9113948385526,
  -83.6470575577013,
  -83.3733229742,
  -83.1287519258876,
  -83.7055644608892,
  -85.3637024819344,
  -84.0770745357732,
  -84.2546813569092,
  -82.8271895022708,
  -85.3749581349455,
  -83.083185436523,
  -82.8972041422597,
  -84.6852352945379,
  -83.9829546581415,
  -83.8233874647682,
  -83.7754627225041,
  -84.458661156064,
  -84.1613154606423,
  1,
  0,
  -85.3443233933269,
  0.619749023351331,
  -85.2265970024743,
  -83.9701795747931,
  -85.9413928698087,
  -85.0042636698926,
  -84.7246802564273,
  -85.4263352482809,
  -85.8352976070202,
  -86.1630850984808,
  -85.7762156854579,
  -86.2834318207355,
  -84.2966799982851,
  -85.7213902119488,
  -85.2371710949369,
  -85.1859823153025,
  -84.750429930045,
  -85.8545355887714,
  -84.8205118788402,
  -85.2744032663555,
  -85.9573230427098,
  -85.4365617059708,
  1,
  0,
  -86.8737341287399,
  0.465202407143357,
  -86.3728002788728,
  -85.5313847256462,
  -86.9230573328542,
  -86.4842147219802,
  -86.7646227663403,
  -87.3598605015695,
  -86.8536527615328,
  -87.1498262023978,
  -87.0503641835501,
  -87.3839291373532,
  -86.3343860188929,
  -86.9938863338804,
  -86.7950361642675,
  -87.0571721559312,
  -86.4980983607854,
  -87.3870476820857,
  -86.9313893894839,
  -86.9307453573103,
  -87.5642722203511,
  -87.1089362797118,
  1,
  0,
  -88.4781108039718,
  0.652792429887406,
  -88.8341852532956,
  -87.4484095913824,
  -89.1921091809334,
  -88.6219527312008,
  -88.4796129947023,
  -89.1582831295067,
  -89.1658062654699,
  -88.6438990224893,
  -88.8503833581861,
  -89.6327180063177,
  -87.894525436089,
  -87.8991400190278,
  -87.9304261885995,
  -87.7370252153672,
  -87.0603552680847,
  -88.5411513307632,
  -88.6080727137572,
  -88.6461705764694,
  -88.205283597296,
  -89.0127062004971,
  1,
  0,
  -90.151452388909,
  0.541994150930576,
  -90.7064788497792,
  -89.8420700279377,
  -90.1526056185954,
  -90.1453270852521,
  -89.7647498794102,
  -89.7995117436275,
  -90.7813069799065,
  -90.7675558420128,
  -90.4175598428734,
  -91.0638185877874,
  -89.955160486982,
  -89.6168528261926,
  -89.1262066331631,
  -91.064160076236,
  -89.570516118708,
  -89.8406734940385,
  -90.0132982877396,
  -90.5807006334641,
  -89.5480346612068,
  -90.2724601032657,
  1,
  0,
  -92.4421608936112,
  0.503315282004311,
  -92.5459202407423,
  -92.3562489810787,
  -93.1953164206791,
  -92.8685339826961,
  -92.0378919924011,
  -92.1806314213932,
  -92.5325413085744,
  -92.3846218336002,
  -92.9924213415886,
  -93.1885447374726,
  -92.5408328283989,
  -91.9435743201227,
  -91.454753180563,
  -93.1901043350342,
  -91.6749928739211,
  -92.3031685488047,
  -92.5171290199029,
  -92.7541928404183,
  -92.4011336798415,
  -91.7806639849898,
  1,
  0,
  -94.4681902156178,
  0.489825936250846,
  -94.8998474559115,
  -94.334835507319,
  -94.9416053931504,
  -94.3659153949,
  -94.5181463034552,
  -93.6338213087418,
  -94.2189570082389,
  -93.9008305453164,
  -94.5187101636614,
  -95.4628607792466,
  -94.6971739912519,
  -94.4806945947315,
  -93.5991757392387,
  -95.1303786660436,
  -94.7894614015878,
  -94.649158316631,
  -94.3460632899551,
  -94.798840860107,
  -94.3301238591895,
  -93.747203733678,
  1,
  0,
  -96.0131391293905,
  0.541306176607581,
  -94.7824503382102,
  -95.441388504928,
  -95.833996471911,
  -95.9112564509097,
  -96.1658137250831,
  -95.5642182471744,
  -95.6579887460958,
  -95.2752197784376,
  -96.4341626700002,
  -96.776558820025,
  -96.1230447934388,
  -96.0651484260252,
  -95.9835880484991,
  -96.9827334587755,
  -96.2694016160763,
  -95.732730558333,
  -96.7065849528139,
  -96.2241184339065,
  -96.5877366967647,
  -95.7446418504019,
  1,
  0,
  -97.4027541676354,
  0.652813106604772,
  -96.265853155181,
  -97.4670380172451,
  -96.971368158447,
  -97.6063908094491,
  -97.9216037903038,
  -97.6460355164666,
  -97.009227108725,
  -96.3297915184508,
  -97.3448391882567,
  -97.5441349727094,
  -96.5090265271993,
  -97.1296136715575,
  -98.5221043789755,
  -97.6507743964081,
  -97.7771499833817,
  -97.6401033684179,
  -98.7832988274921,
  -97.0438914143756,
  -97.9425191828583,
  -96.9503193668084,
  1,
  0,
  -97.2529645564463,
  0.586069351952725,
  -98.0024982427104,
  -97.8522096939917,
  -97.3977864743293,
  -96.892789662928,
  -97.629988928689,
  -97.9978788712623,
  -96.8292600369718,
  -96.7374684004349,
  -96.7775048174264,
  -96.9012500640965,
  -96.4685911622883,
  -97.8366898176759,
  -97.7242378925832,
  -97.1642096224462,
  -97.2878572926613,
  -96.4718005758682,
  -98.3565805368787,
  -96.6352190208034,
  -97.538244155798,
  -96.5572258590829,
  1,
  0,
  -97.1309438246627,
  0.514375366057366,
  -97.1317560674641,
  -97.4571577822107,
  -97.4847661950574,
  -96.9711909778802,
  -97.4677176787405,
  -97.447448730268,
  -97.7705022298722,
  -96.8794594699613,
  -97.5188625003915,
  -97.4431454348796,
  -96.6596458938133,
  -97.4366764318168,
  -95.8794276627087,
  -96.7088636527255,
  -97.3162361774437,
  -96.268668307309,
  -97.6093355366077,
  -96.3536327231437,
  -97.4863154525479,
  -97.3280675884122,
  1,
  0,
  -96.5069257227686,
  0.523281234012032,
  -96.7467671695925,
  -96.6424085265203,
  -96.3763812878887,
  -97.0130758658357,
  -95.972331890033,
  -96.6159609213077,
  -97.2776546225697,
  -96.2994064710218,
  -95.9151653197966,
  -96.6622822286991,
  -95.8705783243338,
  -97.0536910189178,
  -96.2024234561536,
  -96.7942511430282,
  -97.3927525206851,
  -95.7466441771616,
  -97.2773141965562,
  -96.417824236868,
  -95.7942593677802,
  -96.0673417106222,
  1,
  0,
  -95.9205275049126,
  0.536603004167341,
  -95.3215822996912,
  -95.5795222177954,
  -95.5323194840168,
  -96.1357624493126,
  -95.6144943624308,
  -96.3527733871717,
  -96.0454697556676,
  -95.2311958109076,
  -95.1417603094404,
  -96.8655479062696,
  -96.371946928471,
  -96.0098819496979,
  -95.8262365013447,
  -96.8155052384297,
  -96.5740740788006,
  -95.1408797925367,
  -95.7587904389464,
  -96.3840760185934,
  -95.5214739269431,
  -96.1872572417856,
  1,
  0,
  -95.0429368335613,
  0.628524514998862,
  -94.8008558529434,
  -94.7956868564519,
  -94.6259344333918,
  -94.1659893007847,
  -95.6492947700391,
  -95.6566640192352,
  -95.2406320591951,
  -93.9230324791136,
  -94.5651357414412,
  -94.9884461800061,
  -94.555875421725,
  -95.3755848079374,
  -94.761406878359,
  -96.2680526978446,
  -95.8399826233292,
  -94.0504199645337,
  -95.3045818802421,
  -95.3156351108162,
  -95.2788306727092,
  -95.6966949211275,
  1,
  0,
  -93.1549320997899,
  0.560512762703527,
  -93.2766023772751,
  -93.3205888173407,
  -93.1072958449733,
  -93.2385886504849,
  -93.3280207057287,
  -93.2427142814611,
  -92.2590785195527,
  -92.2612288941558,
  -93.0102270774751,
  -93.3220159203791,
  -92.5351561390405,
  -92.7936734764182,
  -93.3072107748886,
  -94.6054916733312,
  -93.6486486671565,
  -92.3729448730808,
  -93.6445133116641,
  -92.7802181670073,
  -93.7258426768737,
  -93.3185811475114,
  1,
  0,
  -90.797920360761,
  0.6642988666026,
  -90.2849982190698,
  -90.9329665383225,
  -91.0518049255848,
  -90.7702667599804,
  -90.9672257554898,
  -90.6193333300192,
  -90.1153773791718,
  -90.0808177109775,
  -90.6480670781738,
  -90.3563343725764,
  -90.7313807251882,
  -89.9144323065766,
  -90.8158633843793,
  -92.202949559093,
  -92.241054487358,
  -89.6628706486736,
  -91.1756251667808,
  -90.804236661414,
  -91.3908398288422,
  -91.191962377549,
  1,
  0,
  -89.1288549739951,
  0.410331902491838,
  -89.012535112191,
  -89.1710049380383,
  -89.3197354579022,
  -89.1982408150046,
  -88.6520698151028,
  -89.150697937191,
  -89.4431509414872,
  -88.2286187863031,
  -89.0117150483643,
  -89.3006927403341,
  -89.2644249212078,
  -88.9314480221549,
  -89.1505123817386,
  -90.1415415644007,
  -89.3484734415413,
  -88.5947803721694,
  -89.7555595441495,
  -88.9221694353238,
  -89.1787077192268,
  -88.8010204860705,
  1,
  0,
  -87.7034038961684,
  0.406651186788673,
  -87.5569451265363,
  -87.8470038708875,
  -87.8528799182909,
  -87.9657536908375,
  -87.3318998356277,
  -87.6733488744854,
  -87.7894726697703,
  -86.9987193946073,
  -87.4541454997986,
  -87.5731483934739,
  -87.6896855971431,
  -87.8423129372548,
  -87.7132868475847,
  -88.7569007032276,
  -87.738533906582,
  -87.9569349925418,
  -88.2401030806914,
  -86.8536105930608,
  -87.7990604860913,
  -87.4343315048746,
  1,
  0,
  -85.9670369299527,
  0.616425358755413,
  -86.0977048921586,
  -85.9432286609474,
  -86.5005937660656,
  -86.2459755154038,
  -85.4279686283908,
  -86.6183491543815,
  -86.0871102372326,
  -85.3687635597989,
  -86.2109554501023,
  -85.4141922017129,
  -85.9982686015159,
  -85.7967439837924,
  -85.6392901296087,
  -87.6121531848301,
  -85.8276985878918,
  -85.3475472856949,
  -86.4819769397337,
  -84.6480042821162,
  -85.786710897998,
  -86.2875026396784,
  1,
  0,
  -84.2468153380011,
  0.678980852878139,
  -84.6402348290489,
  -84.0067127151251,
  -84.7020440975492,
  -84.6394923857764,
  -84.2984082408243,
  -84.2688558536791,
  -84.4226055157147,
  -83.5919696770694,
  -84.3693246815604,
  -84.666470863417,
  -84.4081144328819,
  -83.5572057271096,
  -83.8720809292125,
  -85.9299967402391,
  -83.5523817462794,
  -83.797779881557,
  -85.1532038289882,
  -82.8174412927078,
  -83.6330635146634,
  -84.608919806618,
  1,
  0,
  -83.4654013406077,
  0.504158618540316,
  -83.43615683965,
  -83.2231649367878,
  -84.1666923372488,
  -82.9409893193499,
  -83.623598878262,
  -83.2883203925456,
  -83.2512050107975,
  -83.6154984051146,
  -82.9978160494365,
  -83.3626278361536,
  -84.0012884919007,
  -82.9597999083523,
  -83.4487922318538,
  -84.6586769418291,
  -83.3662830852605,
  -83.052386185786,
  -84.4317439389523,
  -82.7279832957285,
  -83.4428747441822,
  -83.3121279829631,
  1,
  0,
  -83.5926373364373,
  0.340838266010795,
  -83.1717258071961,
  -83.7702303685241,
  -83.4393382390514,
  -83.8124530350813,
  -83.6058668407857,
  -83.1930841993116,
  -83.1690712847679,
  -83.859739772394,
  -83.3270144985789,
  -83.8638088061888,
  -83.6524214910196,
  -83.9932145214825,
  -83.7179942319193,
  -83.9041679815047,
  -83.4622875012006,
  -83.2125930622622,
  -84.0137320182392,
  -82.8861259936835,
  -83.712239871972,
  -84.0856372035828,
  1,
  0,
  -83.6783118229908,
  0.422649391598523,
  -83.5199225034034,
  -83.2797189006197,
  -83.3886881435857,
  -83.5472620134242,
  -83.937552157436,
  -83.8485079078775,
  -82.6846798306751,
  -84.0662722978086,
  -83.7744732005269,
  -84.4847067010024,
  -84.047551066071,
  -84.3555300854735,
  -83.3818410191538,
  -83.8732945173001,
  -83.4473379484045,
  -83.9720544812979,
  -83.8860842121865,
  -83.3488393727354,
  -83.3912385959469,
  -83.3306815048871,
  1,
  0,
  -84.0199877990545,
  0.490828561758972,
  -83.9964400600387,
  -82.9323630193157,
  -83.1463661092985,
  -84.1005038979752,
  -84.4277392694735,
  -84.6147200831895,
  -84.0523247164694,
  -84.6915912964186,
  -83.4748016646019,
  -84.3958750868231,
  -83.9325823837623,
  -84.8474679426462,
  -84.2822225469726,
  -83.7522034323282,
  -84.2463273121007,
  -83.7601830272052,
  -84.2787007792148,
  -83.965289616916,
  -83.904984924622,
  -83.5970688117189,
  1,
  0,
  -85.0560993449489,
  0.609348749779633,
  -84.9344634909765,
  -84.6209606687717,
  -83.1178416876808,
  -84.9339004807394,
  -84.9238849246688,
  -84.9837580277361,
  -85.7262756631681,
  -85.4725778651675,
  -85.3547619441617,
  -84.9580079695846,
  -85.498698856814,
  -85.6027011970056,
  -85.5772105711179,
  -85.059587527782,
  -85.9772207417043,
  -85.3766081918011,
  -85.1550496612367,
  -84.638319374756,
  -84.7194742182708,
  -84.4906838358338,
  1,
  0,
  -86.8987170193109,
  0.555685830213173,
  -86.4072530704543,
  -86.584969100646,
  -86.4061737703146,
  -86.736468138288,
  -85.734733537888,
  -86.4700688989242,
  -87.4318852176892,
  -87.0369906057613,
  -87.7295132739805,
  -87.0050719559291,
  -86.8823608128868,
  -87.597162921181,
  -87.0799158451855,
  -86.3822267436665,
  -87.974243963964,
  -87.2744459310538,
  -86.8268238305576,
  -86.2038714987666,
  -87.2720549728473,
  -86.9381062962346,
  1,
  0,
  -89.1551242203687,
  0.564800970936294,
  -88.8115393223465,
  -88.960280073152,
  -88.6935366714504,
  -89.0584076567008,
  -88.3172429717427,
  -89.2340271152128,
  -89.5734847235696,
  -88.5239073603857,
  -89.1380571871227,
  -88.8571449398955,
  -89.8429936654219,
  -90.3757356351261,
  -89.8962439063456,
  -88.9526555581264,
  -89.8960482128249,
  -88.3577105170629,
  -88.9788996258324,
  -88.8377657622059,
  -88.9962376960649,
  -89.8005658067831,
  1,
  0,
  -91.2499919392495,
  0.520933559335634,
  -90.3627494679593,
  -91.0310153890558,
  -91.4532320361286,
  -91.2243274806738,
  -90.0841311621307,
  -91.5513100316936,
  -91.7085559724402,
  -90.6591891182514,
  -91.6833141038904,
  -91.523764032031,
  -91.4853385138584,
  -92.1715037995136,
  -91.7124217914069,
  -91.2320678493776,
  -91.3503609348771,
  -91.0128380444068,
  -91.3406589002987,
  -91.4977862513202,
  -90.4185356867533,
  -91.4967382189223,
  1,
  0,
  -93.7665586232737,
  0.592726278688507,
  -93.6084731235273,
  -92.7150266004671,
  -92.93662791035,
  -94.2427758813399,
  -92.9513221237336,
  -94.4782205484395,
  -93.4613965920604,
  -94.0519445896766,
  -93.8761270235257,
  -93.4540450003474,
  -94.2260658993084,
  -94.4551693957828,
  -94.3474574847874,
  -93.11422009488,
  -93.5865244705668,
  -93.6363595399861,
  -94.3980585032324,
  -94.2898218351836,
  -93.0426741487504,
  -94.4588616995288,
  1,
  0,
  -96.1683396948662,
  0.622953766013833,
  -96.5584839836625,
  -96.1241593033676,
  -96.5205142527506,
  -96.2875253455179,
  -97.1876481290421,
  -96.3134323808315,
  -95.5629710083224,
  -94.701706167572,
  -95.814897479066,
  -95.4053999693226,
  -96.7341638200332,
  -96.5788905496676,
  -95.9597899302858,
  -95.4371766366835,
  -95.9252272427045,
  -96.7816942315876,
  -97.1571834666335,
  -96.2639775421938,
  -95.6607142650501,
  -96.39123819303,
  1,
  0,
  -98.7314389658309,
  0.567859858623292,
  -98.8282039731593,
  -98.7348939012964,
  -98.6542908886487,
  -98.3076481552789,
  -98.519819507209,
  -99.4080647667658,
  -99.1713900237743,
  -97.9621711524758,
  -98.7901870710625,
  -98.1369568632704,
  -100.257488612278,
  -99.2802381207205,
  -98.748747379414,
  -98.0030837353874,
  -98.228890338373,
  -98.7937647706946,
  -99.3445050903989,
  -98.057588763482,
  -98.8382880280675,
  -98.5625581748605,
  1,
  0,
  -100.665457367462,
  0.383041652768932,
  -100.509024485223,
  -100.643521547079,
  -100.048556694122,
  -100.725772237257,
  -101.227577911903,
  -100.651954363235,
  -100.172127439291,
  -99.9405766907495,
  -101.152289184635,
  -100.995014460609,
  -101.021040195193,
  -100.760224759532,
  -101.12126835372,
  -100.818614144447,
  -100.12823163403,
  -100.652046700195,
  -100.462618641444,
  -100.389573551038,
  -101.043193676916,
  -100.845920678617,
  1,
  0,
  -101.726767953154,
  0.501521912709643,
  -102.079645562366,
  -100.954098620299,
  -102.185786749819,
  -102.453423919938,
  -101.933134471992,
  -101.246037484385,
  -101.028114933304,
  -101.952559690148,
  -102.632716853679,
  -101.690859809492,
  -101.496391958799,
  -101.67551940985,
  -102.103552027602,
  -101.90272608725,
  -101.102382461073,
  -101.964078901428,
  -101.087284703001,
  -101.128012329561,
  -102.217665080474,
  -101.701368008625,
  1,
  0,
  -102.827369920447,
  0.42612035440906,
  -102.053361580033,
  -102.961205826604,
  -102.486337494603,
  -103.681560914865,
  -103.036693592173,
  -102.229604655231,
  -103.17535178894,
  -102.976606949722,
  -103.510900911177,
  -102.70944467484,
  -103.116561028695,
  -102.165920958213,
  -102.442886821632,
  -102.567663111135,
  -102.988174318886,
  -102.924710253757,
  -103.018680494225,
  -102.521727429227,
  -102.931898584947,
  -103.048107020042,
  1,
  0,
  -103.007822721622,
  0.473950603435172,
  -102.201194579583,
  -103.320873435134,
  -103.875744301669,
  -103.788241461323,
  -102.673886984171,
  -102.820861667003,
  -102.806780853534,
  -103.20285335464,
  -103.783764268451,
  -102.921643006883,
  -103.196177282112,
  -102.423737142067,
  -102.837788768713,
  -102.469267209819,
  -103.341735503913,
  -103.325102120121,
  -102.550797207508,
  -102.902662732867,
  -102.583583934055,
  -103.129758618876,
  1,
  0,
  -102.568393472994,
  0.406816704733441,
  -102.545224513523,
  -103.065103563999,
  -103.154875847119,
  -102.379421179435,
  -102.808833290975,
  -103.075212720933,
  -102.296079004832,
  -102.224105271424,
  -102.743424837758,
  -101.733194428369,
  -102.487663887252,
  -101.751556725415,
  -102.214957281131,
  -102.316496244328,
  -102.988805689988,
  -103.00074674737,
  -102.715269905927,
  -102.746177429587,
  -102.522193700744,
  -102.598527189775,
  1,
  0,
  -101.509919246011,
  0.59026793052821,
  -101.599952453863,
  -101.945053329612,
  -101.376889509667,
  -101.446521204779,
  -101.284961784003,
  -102.521128007487,
  -101.960615770018,
  -101.543092409126,
  -101.265456976879,
  -99.9536316459257,
  -101.84139102858,
  -101.214446846441,
  -101.370606881254,
  -101.642604043292,
  -102.050693500545,
  -100.466296516737,
  -101.195543662459,
  -101.867815548695,
  -101.278455894244,
  -102.373227906615,
  1,
  0,
  -100.704046705314,
  0.483778333110551,
  -100.224596329133,
  -100.39638521942,
  -99.7880984567095,
  -100.565631771387,
  -100.823987153071,
  -101.475681450666,
  -99.9952799147803,
  -101.068163760299,
  -100.614984557645,
  -100.445152188837,
  -100.493030706594,
  -100.551576361912,
  -101.233052911146,
  -100.914101715738,
  -100.911859411499,
  -100.608802260268,
  -100.978718044442,
  -100.400034315941,
  -100.733762210603,
  -101.858035366193,
  1,
  0,
  -99.4816219675011,
  0.571988246745464,
  -98.6781514481637,
  -99.4308666304492,
  -98.7112539280284,
  -100.258683615382,
  -99.6734845855623,
  -99.3145676628071,
  -99.1355317626969,
  -100.400069510187,
  -99.2406838237357,
  -99.7575026598027,
  -99.5963523826452,
  -99.9481685480347,
  -99.6348405170254,
  -99.8851788865157,
  -98.2631079373922,
  -98.9844760032606,
  -100.228471867984,
  -99.1124762650159,
  -100.062922234,
  -99.3156490813323,
  1,
  0,
  -97.8728625215172,
  0.429027730426218,
  -97.6829728283837,
  -98.3834195334528,
  -97.8736676513898,
  -97.3847781200609,
  -98.2358551978017,
  -97.3172952014457,
  -98.3695844043718,
  -97.6626656455543,
  -97.8671315517909,
  -98.549568228199,
  -98.1764375586804,
  -97.677266547539,
  -97.5023090364022,
  -97.210706167914,
  -97.6310216885857,
  -98.1293140750917,
  -98.0711869071095,
  -97.2140920035173,
  -97.9665420297083,
  -98.5514360533455,
  1,
  0,
  -96.8819566048715,
  0.332196716045807,
  -96.3558978499601,
  -97.0903627199993,
  -96.5434572542588,
  -96.9137514533108,
  -97.6244401435996,
  -96.8494154909959,
  -96.871588043287,
  -96.2153957632778,
  -97.1783681397848,
  -97.0041780142586,
  -96.8173418922752,
  -96.6564056219113,
  -97.1112470491925,
  -96.7431268090914,
  -96.6714505380968,
  -97.2207666573979,
  -97.3786710118827,
  -96.8678180755114,
  -96.7684979908245,
  -96.7569515785137,
  1,
  0,
  -96.0462692637524,
  0.577226343845158,
  -95.3034923608032,
  -97.1254122411277,
  -95.3993104125053,
  -95.7638409687622,
  -96.6452779557148,
  -96.1275822739427,
  -96.9188845738057,
  -95.9269402114945,
  -95.168839360957,
  -96.1316496864892,
  -95.5016600219004,
  -95.4871604473047,
  -95.7379584837444,
  -95.6275501725919,
  -96.2475543067942,
  -96.2099342051652,
  -96.2908160102495,
  -96.1449461741761,
  -96.033501298814,
  -97.133074108705,
  1,
  0,
  -95.8832436348052,
  0.5122227189872,
  -95.7707076940399,
  -96.3728326946224,
  -95.3661672204631,
  -95.0464532449982,
  -95.4473536963958,
  -95.522951028142,
  -96.6632437680644,
  -94.975391555998,
  -95.8022147041437,
  -96.1451931892319,
  -95.5874620384595,
  -95.528663780452,
  -95.4303446842839,
  -96.4420525554374,
  -96.3041293929457,
  -96.4018157181535,
  -95.98121938481,
  -96.1529019805726,
  -96.6938194466545,
  -96.0299549182358,
  1,
  0,
  -95.9657608171274,
  0.517253902440082,
  -95.9294997422396,
  -95.8821243298236,
  -96.149949239725,
  -96.5445795474535,
  -95.86858292037,
  -95.1686044392758,
  -97.0441321872423,
  -95.555223841694,
  -95.6914664447506,
  -96.0672496919783,
  -95.3042511135667,
  -95.4530843011578,
  -95.4050599377029,
  -95.8800587782649,
  -96.3221784521549,
  -96.4897030018788,
  -95.5856988383172,
  -96.9744312281344,
  -96.1677094829992,
  -95.8316288238195,
  1,
  0,
  -96.8902786876931,
  0.747905286658959,
  -97.5944347848562,
  -96.4393702081889,
  -97.1695436085571,
  -96.7162651300914,
  -96.8270611038207,
  -96.4145735044847,
  -98.9260426696898,
  -97.0919370832481,
  -96.5999585311921,
  -96.0150590911856,
  -95.6818295499523,
  -96.3847632273415,
  -96.7886873690319,
  -97.7691887563088,
  -96.4001726564552,
  -98.1344163850249,
  -96.7986995723008,
  -96.8077478430972,
  -96.3884737876011,
  -96.8573488914328,
  1,
  0,
  -98.3112749593773,
  0.651584644231116,
  -99.1635087407518,
  -97.5225928276016,
  -98.6181781291556,
  -97.7735953129782,
  -98.7309492594147,
  -97.7343845646883,
  -99.294623231998,
  -98.2635787956637,
  -98.7487716696008,
  -98.2388729143493,
  -98.2594335340573,
  -98.6865925401596,
  -98.3668945348982,
  -98.2235681372934,
  -98.2275675795508,
  -99.1468144522984,
  -97.8751074679265,
  -97.1877327686893,
  -97.0224803337955,
  -99.1402523926744,
  1,
  0,
  -100.735562475128,
  0.633479402433959,
  -101.464432957355,
  -100.476330077563,
  -99.8584255820708,
  -101.554338339484,
  -100.603176262596,
  -99.9036547057363,
  -101.18687799872,
  -101.189587791772,
  -101.874028149394,
  -100.249360213198,
  -100.545953738519,
  -100.688558884885,
  -100.57790185735,
  -101.241783239786,
  -100.47988392064,
  -100.916766812569,
  -101.549498601657,
  -99.9698463988276,
  -99.6099742825081,
  -100.770869687925,
  1,
  0,
  -103.668153063479,
  0.524663238553375,
  -103.447114067931,
  -103.58808406918,
  -102.940681529471,
  -104.195140787015,
  -103.481767645905,
  -104.737526692968,
  -103.936281389487,
  -103.494146408983,
  -103.932469350452,
  -102.797856056038,
  -104.234918715107,
  -104.397155562706,
  -102.935226837242,
  -103.906742617131,
  -104.051374066811,
  -103.784986605951,
  -103.50125434272,
  -102.896459225227,
  -103.516250032339,
  -103.58762526692,
  1,
  0,
  -106.261986080793,
  0.525431593355776,
  -106.436080386893,
  -106.243139895472,
  -105.932927812815,
  -106.593767753971,
  -105.983512585247,
  -106.660758237278,
  -105.809186254795,
  -106.429319345565,
  -106.292438891041,
  -105.581181767039,
  -106.727677735991,
  -107.652665796813,
  -105.331474663056,
  -106.406117356357,
  -106.509982900972,
  -106.436735547763,
  -105.695670101298,
  -105.554421827187,
  -106.393752575256,
  -106.568910181044,
  1,
  0,
  -108.421330759647,
  0.468610771785669,
  -108.753392763996,
  -109.247541890774,
  -108.049159760633,
  -108.352249541699,
  -108.478820469151,
  -107.773873631112,
  -108.159377325207,
  -107.884503487351,
  -108.421762964718,
  -108.095783170786,
  -108.072368737264,
  -109.238364431548,
  -108.524626753988,
  -107.643271321697,
  -108.560425890812,
  -108.487362947444,
  -108.627962749439,
  -108.810896106545,
  -109.190961874365,
  -108.053909374418,
  1,
  0,
  -110.397364884295,
  0.569562388318629,
  -110.899152422921,
  -110.86354036394,
  -110.095763250423,
  -110.074647643198,
  -110.560285841023,
  -110.269831588696,
  -110.119090427302,
  -109.733976892675,
  -110.833508760142,
  -110.198359645634,
  -108.906855311739,
  -109.973875672141,
  -111.2718812599,
  -109.810366346295,
  -110.504846050263,
  -111.096026246134,
  -111.049950045791,
  -110.829120388455,
  -110.2218415268,
  -110.634378002421,
  1,
  0,
  -112.761293937123,
  0.739117621555885,
  -113.192337714718,
  -112.363221321844,
  -112.666579351441,
  -112.81332223282,
  -113.916341449047,
  -112.476026750343,
  -111.860333819521,
  -112.104313708277,
  -112.608316741938,
  -112.810461568394,
  -112.044863460964,
  -113.191483106881,
  -113.995958986578,
  -112.101223640721,
  -113.175750699074,
  -112.850201937124,
  -111.059046216041,
  -112.745500949822,
  -113.390804410274,
  -113.859790676641,
  1,
  0,
  -114.441580061888,
  0.774888711398031,
  -115.531445913785,
  -114.670756950175,
  -115.473741958817,
  -114.385123789049,
  -115.821875022266,
  -114.24200231859,
  -113.490933249805,
  -113.872655607098,
  -113.90109290159,
  -114.199323659994,
  -113.622769055719,
  -114.058893133529,
  -114.317546315126,
  -113.860467600759,
  -115.36799246992,
  -115.830491536102,
  -113.26806890074,
  -114.454785918392,
  -113.954211375115,
  -114.507423561183,
  1,
  0,
  -115.817959126574,
  0.456492943547543,
  -116.792849827018,
  -115.964281433283,
  -115.98223662248,
  -116.165913568681,
  -115.552391498172,
  -115.329640625018,
  -115.802003136781,
  -116.324958327081,
  -115.278685638513,
  -115.161807521716,
  -116.160768001874,
  -116.050777630103,
  -115.597899403714,
  -115.634672996546,
  -115.67868816042,
  -115.68425205075,
  -115.018470174635,
  -115.858942665838,
  -116.599283781901,
  -115.720659466946,
  1,
  0,
  -116.3919544481,
  0.707253567703365,
  -117.304646364893,
  -116.377638365284,
  -117.49085461924,
  -116.84061917187,
  -115.731794626652,
  -115.97920953659,
  -116.758188315265,
  -115.676631350431,
  -116.309113762358,
  -116.277442447514,
  -116.850250719247,
  -115.166479681638,
  -116.9356279348,
  -116.805604460499,
  -117.677076777287,
  -115.969524110618,
  -116.336563432284,
  -116.481716837438,
  -115.698633327025,
  -115.171473121067,
  1,
  0,
  -117.207898985147,
  0.606665032121602,
  -118.492099604015,
  -117.666187419807,
  -116.933688819566,
  -116.104863966539,
  -117.080967320668,
  -117.157945022934,
  -116.775241058274,
  -116.902130473978,
  -116.932524700977,
  -117.020963579582,
  -117.537383455588,
  -116.355025280208,
  -117.654358754613,
  -116.929479651006,
  -117.014660261558,
  -117.202956322887,
  -117.266552206922,
  -117.379928284088,
  -118.699237700987,
  -117.05178581875,
  1,
  0,
  -117.318506070392,
  0.514349537005558,
  -117.80684935736,
  -118.208137562892,
  -117.150556292348,
  -117.829745726472,
  -118.218770457003,
  -117.575718238827,
  -116.865897153931,
  -116.887305681414,
  -117.251887711568,
  -117.508449953562,
  -117.112837297727,
  -117.003550642041,
  -117.078174523158,
  -117.332583672664,
  -116.605417762894,
  -116.393727208043,
  -117.542872971947,
  -117.083382268864,
  -116.868954708656,
  -118.045302216477,
  1,
  0,
  -117.11657837434,
  0.596429661938693,
  -117.664285591674,
  -117.715175437412,
  -117.095358244831,
  -117.46634833677,
  -116.496423498313,
  -117.936238050847,
  -115.726019698122,
  -117.144303728446,
  -116.499491917917,
  -117.211970760105,
  -117.257717593359,
  -117.035992250587,
  -117.460518527683,
  -117.948912445226,
  -116.010195860252,
  -117.082822000276,
  -116.779573715312,
  -117.549443946502,
  -116.783931511042,
  -117.466844372128,
  1,
  0,
  -116.322440738394,
  0.592280588347771,
  -115.929292993634,
  -117.114639589426,
  -115.94535402613,
  -116.473390963864,
  -116.632961949903,
  -116.649285478772,
  -115.813705691598,
  -117.65662728939,
  -116.710544567348,
  -115.592531263828,
  -116.020229061804,
  -116.046664531086,
  -115.964189067315,
  -115.908919673481,
  -115.617211158916,
  -116.233158729555,
  -115.620644575816,
  -117.296880249612,
  -116.936505734628,
  -116.286078171765,
  1,
  0,
  -115.46803604777,
  0.571745150484217,
  -114.959372128304,
  -114.908404135482,
  -115.116829206398,
  -116.11912191022,
  -114.951326825468,
  -115.525095658087,
  -116.248095508271,
  -115.814704605847,
  -116.281670287924,
  -115.079452057082,
  -116.127650573511,
  -116.110327563646,
  -115.349935550841,
  -115.706897223822,
  -115.112012218144,
  -114.3871892081,
  -115.579230844484,
  -116.137019774124,
  -114.843722915195,
  -115.002662760439,
  1,
  0,
  -114.036518473936,
  0.702735143833195,
  -114.526225255613,
  -113.322998046308,
  -113.552189183885,
  -114.220325424094,
  -113.547829762264,
  -114.258921174233,
  -113.741860527493,
  -112.811707522611,
  -114.72510872254,
  -112.903907684638,
  -115.082330034588,
  -113.982513326312,
  -113.580858461072,
  -113.61239925725,
  -114.587099588631,
  -115.062058814181,
  -115.361636577825,
  -114.088737311207,
  -113.671990979601,
  -114.089671824373,
  1,
  0,
  -113.087106173794,
  0.467436931785377,
  -113.4686779178,
  -113.640366452914,
  -112.664255466759,
  -113.473778640741,
  -113.016733818639,
  -113.004831243238,
  -112.522308160774,
  -112.61131652223,
  -113.09361043543,
  -112.91788281751,
  -113.736251414254,
  -112.224202789297,
  -112.911213700048,
  -113.520020504946,
  -112.871717615901,
  -113.641603554489,
  -112.421989965509,
  -113.839674546844,
  -112.94184433042,
  -113.21984357813,
  1,
  0,
  -112.637391008694,
  0.602899239314587,
  -113.114299740348,
  -113.167160362112,
  -112.596534149343,
  -112.322614626502,
  -112.669671696858,
  -112.704021447298,
  -111.048216011003,
  -112.15128231594,
  -111.809884861448,
  -112.73436514365,
  -112.896583943915,
  -112.952349227544,
  -112.157950889863,
  -113.115903180424,
  -113.322997378358,
  -112.546374636721,
  -112.747457228409,
  -113.20254042475,
  -111.913665768861,
  -113.573947140524,
  1,
  0,
  -112.970154215244,
  0.614427114927017,
  -113.499045597992,
  -113.376450360654,
  -113.746817276102,
  -112.24041779486,
  -113.002856017116,
  -113.541429234354,
  -112.338255432545,
  -111.931368208818,
  -112.394789014235,
  -113.51992014896,
  -112.978171304223,
  -112.936306451619,
  -113.700873072598,
  -111.985758224669,
  -112.532945865737,
  -113.307101619572,
  -112.641285160783,
  -113.310314970871,
  -112.500272126717,
  -113.918706422452,
  1,
  0,
  -113.074079041855,
  0.640763535719605,
  -113.083015224459,
  -112.755434637307,
  -112.757531812416,
  -112.798348658342,
  -111.748739634702,
  -114.020018844661,
  -112.679063611269,
  -113.776635323534,
  -112.317773397721,
  -113.881738937686,
  -113.015282924347,
  -112.716968377731,
  -113.076684666914,
  -113.252182827301,
  -113.646146828557,
  -113.215428979991,
  -112.011634423972,
  -112.975665959312,
  -114.051613732917,
  -113.701672033962,
  1,
  0,
  -114.324501022091,
  0.561697095203742,
  -115.314470217772,
  -114.86407291297,
  -113.737273234568,
  -113.535806037798,
  -114.710862944789,
  -114.617150354445,
  -113.817992198473,
  -114.08343766483,
  -114.485031588627,
  -113.62693390098,
  -114.102587203975,
  -113.636855953791,
  -114.77481611648,
  -114.268720513406,
  -113.523791237234,
  -114.235391955355,
  -114.919832024081,
  -114.736484271942,
  -115.214287085439,
  -114.284223024867,
  1,
  0,
  -115.835710225481,
  0.67127531077984,
  -117.075161306181,
  -115.826397700452,
  -115.305167215481,
  -115.390040040095,
  -116.264633184043,
  -115.997117893299,
  -114.990492714871,
  -116.627332313786,
  -115.793323578873,
  -115.744189167774,
  -114.90194742078,
  -116.476930735389,
  -116.081505526047,
  -115.889374688122,
  -115.513229922901,
  -116.306311087598,
  -115.916085629616,
  -114.504347702958,
  -115.207766338061,
  -116.902850343301,
  1,
  0,
  -117.427743175893,
  0.50501369414957,
  -117.187442935354,
  -117.355085039024,
  -117.673167552483,
  -117.885662017991,
  -116.350426778965,
  -117.648255819361,
  -117.296536685894,
  -117.958984332972,
  -117.0850399471,
  -117.014639342715,
  -117.242654488538,
  -117.228160070635,
  -117.773740235906,
  -117.671617301216,
  -117.645546125007,
  -117.50264656078,
  -117.36930465956,
  -116.801639825878,
  -117.064571960983,
  -118.799741837506,
  1,
  0,
  -119.858242298354,
  0.667962646272678,
  -119.616059536425,
  -119.512588206467,
  -118.825435703653,
  -119.364860168008,
  -120.271883098727,
  -120.468806638362,
  -119.684544272421,
  -120.225032946629,
  -118.557171895513,
  -119.089342505371,
  -119.392127252463,
  -120.71167289778,
  -119.888418604067,
  -120.898330133954,
  -120.234136228745,
  -120.607534528583,
  -119.821059803154,
  -120.206385570741,
  -119.139680275539,
  -120.649775700474,
  1,
  0,
  -121.716741701709,
  0.6236129031678,
  -121.916875444564,
  -122.497130746201,
  -122.022271718196,
  -121.003750539533,
  -122.071305571734,
  -122.085469193702,
  -122.178552207815,
  -122.490343772007,
  -120.751197787881,
  -122.150260139569,
  -121.0381140275,
  -121.703735301752,
  -122.575803994272,
  -122.061283994352,
  -120.654633383932,
  -121.913849474729,
  -121.297064838838,
  -120.896284052813,
  -122.027421640546,
  -120.999486204239,
  1,
  0,
  -123.398666146951,
  0.67282258080477,
  -123.157137024778,
  -123.929673473166,
  -123.707151585462,
  -122.927809722143,
  -123.459837688809,
  -122.636548278345,
  -123.007443714423,
  -123.956676826983,
  -123.821459811515,
  -124.832445907493,
  -123.710196297994,
  -124.317595471656,
  -123.816595417877,
  -123.021913829818,
  -123.39127201075,
  -121.956664199803,
  -123.169711127613,
  -122.279123970079,
  -123.521330299519,
  -123.352736280801,
  1,
  0,
  -125.554418264201,
  0.743644635501247,
  -126.910073156493,
  -126.169566397721,
  -125.90924702578,
  -125.485135572125,
  -125.486267460297,
  -124.564368868878,
  -125.526603067813,
  -125.001269360597,
  -125.839261725009,
  -125.070279871016,
  -126.483607123121,
  -124.57851563885,
  -125.781927362443,
  -126.124060834546,
  -126.887071692972,
  -125.152477786917,
  -125.981148154634,
  -124.437045330904,
  -124.874179441673,
  -124.826259412228,
  1,
  0,
  -127.508548797848,
  0.561064609835011,
  -127.636017052393,
  -127.157055313624,
  -128.175756372965,
  -128.503277600513,
  -127.030232531691,
  -127.106762981589,
  -127.079771729131,
  -127.365066357773,
  -127.665904827338,
  -127.230543661782,
  -128.052966560851,
  -126.341994707129,
  -126.778233463044,
  -127.808835470703,
  -128.356938185033,
  -127.884215524193,
  -127.833919025048,
  -127.558541728087,
  -127.735463124503,
  -126.869479739565,
  1,
  0,
  -129.061601546235,
  0.62574280541541,
  -128.880480428657,
  -128.158452131662,
  -129.636511744996,
  -129.297612176542,
  -128.111858356722,
  -129.374339881603,
  -129.115789899323,
  -128.378306082224,
  -129.349592119967,
  -129.697377707872,
  -129.230534046051,
  -128.6195997038,
  -129.976857742777,
  -128.544984600499,
  -130.313959049719,
  -128.388729018652,
  -128.533238510154,
  -129.351581094099,
  -128.624245615147,
  -129.647981014233,
  1,
  0,
  -129.703213514821,
  0.696414116954859,
  -129.890694558264,
  -129.180114833712,
  -129.551724089716,
  -129.285772884427,
  -129.701334994094,
  -129.358593102969,
  -129.671995027445,
  -129.920189259281,
  -131.222612361792,
  -130.193408318807,
  -130.357655744316,
  -130.083354872614,
  -129.622320846289,
  -127.856039771164,
  -130.547728979987,
  -130.017010549021,
  -129.7499305014,
  -129.383556192017,
  -128.66611535375,
  -129.804118055362,
  1,
  0,
  -129.851171980054,
  0.525035093058829,
  -129.454823790709,
  -129.18227414044,
  -129.906648200808,
  -129.7481604568,
  -129.785359538104,
  -129.239579073008,
  -129.365986242264,
  -130.071479301698,
  -130.128299857238,
  -129.587620739656,
  -129.420709491977,
  -131.574963057088,
  -129.795293354092,
  -129.76299210281,
  -130.132145642496,
  -129.962422992515,
  -130.41522662255,
  -129.846912616599,
  -129.480790266976,
  -130.161752113257,
  1,
  0,
  -129.269364206108,
  0.855525333712884,
  -129.738681735277,
  -127.426294245011,
  -127.840810562567,
  -129.819327524255,
  -129.080858704145,
  -129.984956453949,
  -129.118613590832,
  -130.728181032791,
  -129.960455137354,
  -129.82823945339,
  -129.323499261505,
  -130.529351351435,
  -128.67382617528,
  -129.702981509604,
  -129.03794513491,
  -128.460721584407,
  -129.394127353804,
  -128.112222327436,
  -128.953431177152,
  -129.672759807065,
  1,
  0,
  -128.551414839308,
  0.574718628812939,
  -128.691560263334,
  -128.615691279838,
  -128.700196890787,
  -129.358707309526,
  -128.804807343391,
  -129.755538632383,
  -127.846707229367,
  -129.320696389693,
  -127.95861251483,
  -128.525540155536,
  -128.153374058645,
  -128.426571439256,
  -127.789733476517,
  -129.27097660959,
  -127.981007973777,
  -128.416640786142,
  -128.250533888142,
  -129.133149893563,
  -128.04330708163,
  -127.984943570214,
  1,
  0,
  -128.013011086853,
  0.71230821629712,
  -127.721768814492,
  -127.573382802309,
  -127.779957800912,
  -128.041787082332,
  -127.720425765372,
  -127.029657138953,
  -127.529093154967,
  -128.495110632296,
  -128.878664198524,
  -127.587384789263,
  -128.045646696014,
  -127.256259522911,
  -128.036327068439,
  -128.604488499538,
  -129.650883235661,
  -127.016625424092,
  -127.563750679518,
  -127.966185874905,
  -129.403683780712,
  -128.359138775858,
  1,
  0,
  -126.656326795667,
  0.587610827348444,
  -126.893430118266,
  -127.00831618229,
  -127.174184593121,
  -126.269013831404,
  -126.783760712186,
  -127.372914071477,
  -125.76279187474,
  -125.48752779528,
  -126.763597063754,
  -127.378301177018,
  -127.17713177323,
  -127.371775073538,
  -126.53754422818,
  -127.109621407507,
  -126.719806260747,
  -126.334975133391,
  -126.651803980625,
  -125.419789152858,
  -126.36806590418,
  -126.542185579552,
  1,
  0,
  -124.781007131589,
  0.61485596564136,
  -125.523525617421,
  -125.207863182511,
  -125.779736812233,
  -125.215907579455,
  -123.696298868086,
  -125.585256130354,
  -124.463447489316,
  -124.753112890422,
  -123.768765449943,
  -125.332400558715,
  -124.220506533639,
  -123.836979828676,
  -124.521099677104,
  -124.878845805974,
  -124.878831592214,
  -124.481851074502,
  -125.010208983715,
  -125.091341769495,
  -125.167211393372,
  -124.206951394635,
  1,
  0,
  -123.531330832396,
  0.56131531144717,
  -123.974173636683,
  -124.239447245673,
  -123.633479739126,
  -122.92617157033,
  -122.884715243521,
  -123.081493081613,
  -124.101969283275,
  -123.910850178996,
  -122.286499563398,
  -123.933052675092,
  -123.202471095857,
  -123.400497485142,
  -124.439693772866,
  -123.900110192149,
  -123.241019608139,
  -123.851048938003,
  -122.787909481856,
  -124.032130530404,
  -123.389263292666,
  -123.410620033127,
  1,
  0,
  -123.033182329361,
  0.774574770709346,
  -123.050142242225,
  -122.362119042299,
  -122.544208718761,
  -123.571886939793,
  -122.386104978634,
  -123.088423474721,
  -123.892676390396,
  -123.563120658782,
  -122.412875537742,
  -123.478268874734,
  -124.272597994591,
  -122.132293824919,
  -122.661617437223,
  -124.156133766126,
  -124.206762304862,
  -121.383842270663,
  -122.875663226298,
  -122.385577314105,
  -122.905623127807,
  -123.333708462533,
  1,
  0,
  -122.226615633053,
  0.574712973199319,
  -122.060826856824,
  -122.212448857926,
  -122.247204953982,
  -121.864908153391,
  -121.122323722497,
  -121.874955881429,
  -122.955603005848,
  -122.849977515433,
  -122.501864338445,
  -122.500466622706,
  -121.383767554477,
  -122.211306705208,
  -122.529367177333,
  -122.570029743192,
  -123.077348601993,
  -122.977964237765,
  -121.070077377404,
  -122.488475870153,
  -122.018322556379,
  -122.015072928671,
  1,
  0,
  -121.369682642115,
  0.599031717260762,
  -121.565186952579,
  -120.496503880472,
  -121.542583435199,
  -120.562886989419,
  -121.179182621417,
  -121.982578477472,
  -121.275998116142,
  -122.498259919992,
  -120.591570651951,
  -120.949729973712,
  -120.619398672894,
  -121.322149418017,
  -121.188935999883,
  -122.515488512527,
  -120.784956839964,
  -122.002382654445,
  -121.733903197588,
  -121.530700377625,
  -121.532325138513,
  -121.518931012484,
  1,
  0,
  -121.476591421585,
  0.764486178950418,
  -122.083033570287,
  -119.470721476722,
  -121.102581571076,
  -121.748544642167,
  -121.276261764847,
  -121.815360131539,
  -121.658693748031,
  -121.534757151993,
  -121.328599402159,
  -121.85870733778,
  -121.808985554152,
  -122.359793320751,
  -120.974781948987,
  -121.954592511067,
  -120.5436510154,
  -122.783139558205,
  -122.348017046896,
  -120.339868645195,
  -121.437332656183,
  -121.104405378271,
  1,
  0,
  -122.005287830001,
  0.706384153024943,
  -121.487498120935,
  -121.196536344087,
  -121.289400647168,
  -122.223500233683,
  -121.479973123605,
  -122.499278764771,
  -121.393150668735,
  -122.206349845142,
  -121.750500049226,
  -122.684186031047,
  -121.93126224814,
  -122.364315677402,
  -122.172595071571,
  -121.832353365469,
  -123.683749070513,
  -121.696306788821,
  -120.513081439726,
  -122.626092506027,
  -122.893573923958,
  -122.18205268,
  1,
  0,
  -123.045075712997,
  0.498483146261414,
  -123.315576547664,
  -123.006562457811,
  -122.94177887781,
  -122.530041801025,
  -122.434678734375,
  -122.86394822994,
  -123.368702697996,
  -122.764682299121,
  -122.128621981313,
  -123.643606411351,
  -122.568115479156,
  -122.178233319581,
  -123.120238896858,
  -122.996316727808,
  -123.534448890334,
  -123.805002645439,
  -123.156953944257,
  -123.627796751736,
  -123.250026063088,
  -123.666181503277,
  1,
  0,
  -124.365300370462,
  0.638587525227558,
  -125.522374514515,
  -124.047373654634,
  -125.467177958378,
  -124.465305546593,
  -123.964760722129,
  -124.182133545228,
  -124.047273992578,
  -123.78993067996,
  -123.322570369441,
  -123.998857077958,
  -123.757223326212,
  -124.642930150684,
  -124.089057252738,
  -123.988447566728,
  -124.668124410788,
  -123.671374217399,
  -124.195030513387,
  -125.014549904482,
  -125.362268086621,
  -125.109243918782,
  1,
  0,
  -125.629239865845,
  0.548083170694839,
  -125.626877092459,
  -125.33135604797,
  -125.121146047006,
  -125.9807219411,
  -125.822995776656,
  -124.898442295222,
  -125.367616316597,
  -125.48293348492,
  -125.391681537847,
  -126.403504104797,
  -125.433869463002,
  -125.149271400328,
  -124.965277162461,
  -125.887380682799,
  -125.840918341264,
  -124.661925140018,
  -125.948760486639,
  -126.520184038321,
  -126.653416343323,
  -126.096519614174,
  1,
  0,
  -127.261128725433,
  0.616272627011083,
  -128.311109011234,
  -126.933436558329,
  -126.668564831253,
  -126.445362754228,
  -127.965714380475,
  -126.835945781065,
  -127.592194058734,
  -126.795821252892,
  -127.530366437643,
  -127.87201624273,
  -126.644730286571,
  -126.505920794519,
  -126.472818225547,
  -128.153679450488,
  -126.993863307714,
  -127.22572727346,
  -127.748432512375,
  -127.433438026122,
  -126.968242738801,
  -128.125190584487,
  1,
  0,
  -128.119617929503,
  0.599386636524668,
  -128.494389185081,
  -128.470130287128,
  -128.305519439239,
  -127.752778746152,
  -128.645986691333,
  -128.073951844153,
  -127.721100141215,
  -128.276397283613,
  -127.508392226697,
  -129.634369999873,
  -128.153439388838,
  -127.813468468892,
  -128.80143934376,
  -126.705746082692,
  -128.071532628445,
  -127.949007105155,
  -127.971525458403,
  -127.480443279265,
  -127.973186887423,
  -128.589554102708,
  1,
  0,
  -129.177133996621,
  0.651269405417225,
  -129.737319202173,
  -129.436489177729,
  -128.972557937148,
  -128.155758008434,
  -128.477897977703,
  -129.094524453918,
  -128.671539680385,
  -129.851217406093,
  -128.435538811783,
  -129.384442942309,
  -130.136606974116,
  -129.422498733925,
  -129.518293774816,
  -129.645510655922,
  -129.322253740341,
  -128.891491891663,
  -130.096280569085,
  -127.667782445645,
  -129.640438005871,
  -128.984237543362,
  1,
  0,
  -129.566689071927,
  0.512148743117158,
  -128.940450580461,
  -129.461742915561,
  -129.164595804117,
  -129.382761172406,
  -129.7775343054,
  -129.006421833273,
  -129.279082655157,
  -129.889767149823,
  -128.805309954415,
  -130.533289762716,
  -130.459162164881,
  -129.678963714077,
  -130.22646578346,
  -129.391602574475,
  -129.237518361362,
  -129.232888699482,
  -129.233476019977,
  -130.265682248758,
  -130.002663495855,
  -129.364402242886,
  1,
  0,
  -129.49301241609,
  0.459439888012748,
  -129.23601461473,
  -130.149873393063,
  -129.388355033029,
  -129.007119902649,
  -129.997805101096,
  -129.476895451687,
  -129.194135386637,
  -129.751724833062,
  -128.914930314855,
  -129.465887707788,
  -129.297080852389,
  -128.956569711348,
  -129.494589433312,
  -129.625802628219,
  -130.180560490869,
  -130.395442253029,
  -129.546718278829,
  -129.59007208805,
  -129.624632169665,
  -128.566038677503,
  1,
  0,
  -128.649047773072,
  0.652518917899897,
  -129.659304511709,
  -128.713700564804,
  -128.450901381077,
  -127.795328699304,
  -128.529838413923,
  -128.268626646659,
  -128.050212669717,
  -129.74794693107,
  -128.682191411941,
  -128.033912343189,
  -128.768418230089,
  -128.929795972662,
  -129.400118422218,
  -128.260065357726,
  -127.894896573161,
  -129.018238565612,
  -127.595041841236,
  -128.22358438456,
  -129.416820666006,
  -129.542011874777,
  1,
  0,
  -127.724016009041,
  0.464702552266715,
  -127.837041470376,
  -128.550090078916,
  -127.542313566871,
  -127.985819552776,
  -128.27783553402,
  -127.351608802174,
  -127.199507840268,
  -127.554024992458,
  -127.060179832241,
  -127.758526987567,
  -127.825969082395,
  -127.127397642944,
  -127.969112815382,
  -128.410787897823,
  -127.549894574288,
  -127.434870594268,
  -127.199541069138,
  -128.230873696359,
  -128.335244159287,
  -127.279679991269,
  1,
  0,
  -126.590368968964,
  0.495122281059017,
  -126.768402633976,
  -126.628042678939,
  -125.87963364508,
  -126.154510195235,
  -126.97332071267,
  -126.781299234355,
  -125.82440525723,
  -126.63379119845,
  -126.258055061473,
  -126.244110681786,
  -127.416753274279,
  -126.743081786921,
  -127.012701437608,
  -127.562345652799,
  -126.812857435959,
  -126.644421529629,
  -126.199082801897,
  -125.792724666293,
  -127.064717624132,
  -126.413121870569,
  1,
  0,
  -125.024486624781,
  0.590412821024385,
  -124.413359113975,
  -125.358891747863,
  -124.457776981873,
  -125.423577392386,
  -125.570839750747,
  -124.862169085908,
  -123.846731446473,
  -125.272045262733,
  -125.650817048006,
  -125.546333192572,
  -125.651409565988,
  -126.187970274596,
  -125.374599257859,
  -124.45044441471,
  -124.915848770949,
  -125.07757023952,
  -124.131093169631,
  -124.730960848667,
  -124.729792520927,
  -124.837502410246,
  1,
  0,
  -123.697795409273,
  0.575460757880197,
  -123.943365404815,
  -124.531814037838,
  -123.408900304266,
  -124.151553708721,
  -123.400605928681,
  -123.223637277577,
  -123.751641430128,
  -123.313545723838,
  -124.131851515334,
  -124.05705485296,
  -123.48209648535,
  -123.345939021617,
  -124.128067057754,
  -123.457017392294,
  -122.05538132331,
  -124.661591664916,
  -123.523834450581,
  -123.788299664944,
  -124.227863207829,
  -123.371847732712,
  1,
  0,
  -121.645392310806,
  0.726991604787315,
  -122.456662852274,
  -121.388002911265,
  -121.230085935534,
  -122.33165011839,
  -121.954928776945,
  -121.649379180894,
  -121.662355022019,
  -121.515045056361,
  -121.010574386816,
  -122.100903231772,
  -120.808912323464,
  -120.577381378964,
  -121.953463155063,
  -121.849216066826,
  -120.015710727637,
  -122.579900154192,
  -122.653091043362,
  -122.431585441754,
  -120.795637466483,
  -121.9433609861,
  1,
  0,
  -119.934446371953,
  0.586562050927714,
  -120.493972864393,
  -120.548505149575,
  -120.018542349882,
  -119.375976850224,
  -120.327069323586,
  -119.987470016464,
  -119.950973584376,
  -120.803544815057,
  -120.348053123517,
  -118.981278549449,
  -120.02179860515,
  -119.261290710816,
  -119.503449625856,
  -119.971475755113,
  -121.116202018812,
  -119.61541752469,
  -120.167579393077,
  -119.702042305596,
  -118.837009437737,
  -119.657275435696,
  1,
  0,
  -118.505333775081,
  0.646387435855185,
  -118.581449043247,
  -118.713073027506,
  -118.571410558204,
  -117.699112915898,
  -118.457174892255,
  -119.183297861986,
  -118.694944013375,
  -117.654437133935,
  -119.263559847009,
  -119.313859859153,
  -118.487375782202,
  -118.763216568005,
  -117.391175941594,
  -117.577063563446,
  -119.368924704207,
  -118.752054371501,
  -118.522026331146,
  -118.058083232368,
  -119.423562783834,
  -117.630873070745,
  1,
  0,
  -117.754740079599,
  0.643245605556785,
  -117.80772353186,
  -118.428594661453,
  -118.74875723905,
  -117.210179571771,
  -118.443335725512,
  -118.197857758535,
  -117.946915629507,
  -116.754991170945,
  -118.297607586086,
  -117.881052291055,
  -117.591292497981,
  -117.090262582783,
  -117.312669783432,
  -118.323000469319,
  -118.057861371741,
  -116.950066386351,
  -117.813989230602,
  -116.750126525711,
  -118.569931541564,
  -116.918586036725,
  1,
  0,
  -116.970534060309,
  0.573096799767682,
  -117.399154354887,
  -116.656851540081,
  -116.329805331847,
  -116.228312326086,
  -117.707392192365,
  -116.871007720485,
  -116.288866775332,
  -116.1366864294,
  -117.688706865364,
  -117.784265615422,
  -116.92570060985,
  -117.271288897447,
  -116.588516350088,
  -117.045390258909,
  -117.004740690961,
  -116.631453687435,
  -117.150581423983,
  -118.008740604118,
  -116.296656493962,
  -117.396563038151,
  1,
  0,
  -116.496061133548,
  0.481481293775507,
  -116.443103606845,
  -115.842234231319,
  -116.969670123739,
  -116.683124336494,
  -116.906278949765,
  -117.281335396157,
  -116.661360878115,
  -116.749838955678,
  -116.46046355999,
  -116.391199005863,
  -117.038622449842,
  -115.896262084523,
  -116.66664640599,
  -116.301539367262,
  -116.882255032802,
  -116.497715107683,
  -116.144617308042,
  -116.847585082412,
  -115.309184146185,
  -115.948186642265,
  1,
  0,
  -116.462158515969,
  0.572184630458611,
  -116.235916613615,
  -117.150619029263,
  -115.544835973526,
  -116.384783834204,
  -115.648299130085,
  -116.995498047975,
  -116.639090956967,
  -117.017616265559,
  -116.583335817501,
  -116.392109264513,
  -117.316499680278,
  -115.771142339454,
  -116.290361052357,
  -116.395410974447,
  -116.369830794992,
  -116.763403607231,
  -115.842725317065,
  -117.607758138317,
  -115.755687347291,
  -116.538246134741,
  1,
  0,
  -116.567712731209,
  0.795865926039,
  -116.732621644931,
  -118.078384976247,
  -115.685757561641,
  -115.136667560277,
  -115.210934700563,
  -117.265485608373,
  -115.332055667656,
  -117.465230340465,
  -116.254682890713,
  -117.14192151853,
  -117.270148642583,
  -116.414705885715,
  -116.840267573956,
  -117.465820558415,
  -116.812063936375,
  -116.072647790299,
  -116.582109011152,
  -116.285077532251,
  -116.738489887408,
  -116.56918133663,
  1,
  0,
  -116.495347850122,
  0.43177424670301,
  -116.226744069429,
  -116.63418439677,
  -115.796635294744,
  -115.570696900433,
  -116.613787935187,
  -117.055463659465,
  -116.622634560713,
  -116.872803425047,
  -116.838077991223,
  -115.839491655303,
  -116.504513303244,
  -116.267783191858,
  -116.832531317297,
  -116.712541932267,
  -116.703012552182,
  -116.852924892857,
  -115.786522922412,
  -116.69353197817,
  -116.857414788581,
  -116.625660235261,
  1,
  0,
  -117.386495103529,
  0.5122856834882,
  -117.410286638254,
  -117.668481692755,
  -117.438248137392,
  -117.673379277746,
  -116.957453720474,
  -117.433928861672,
  -117.401055831248,
  -117.576325542278,
  -117.505632622209,
  -117.635136738956,
  -116.887505902345,
  -117.898056176444,
  -117.72134647343,
  -116.960539527183,
  -116.261184472054,
  -118.039151263407,
  -117.563814772844,
  -118.346929874547,
  -116.499887035005,
  -116.851557510333,
  1,
  0,
  -117.879403481579,
  0.488048064054362,
  -117.603675123344,
  -117.346568656791,
  -117.709173405382,
  -117.789321678711,
  -117.862022147203,
  -118.793863978172,
  -118.459930667247,
  -117.817606898704,
  -117.560514611623,
  -118.249656738543,
  -117.756090026156,
  -117.432084570675,
  -117.533476033813,
  -119.197639740226,
  -117.623470223497,
  -117.720602928412,
  -117.925019184641,
  -117.977265891329,
  -117.169182455747,
  -118.060904671356,
  1,
  0,
  -118.127893918439,
  0.579836246887522,
  -117.734021192518,
  -117.963640512716,
  -118.860504826094,
  -117.392226364942,
  -118.644640050491,
  -118.397333210764,
  -117.272478263679,
  -118.716867894024,
  -117.225688800706,
  -118.603748382351,
  -117.696208580599,
  -117.64010691539,
  -117.160309518839,
  -118.653308096911,
  -118.795100853585,
  -118.510189233905,
  -118.515086677277,
  -118.229697867095,
  -118.618905695146,
  -117.927815431742,
  1,
  0,
  -118.577292677144,
  0.699418312957747,
  -118.25810249383,
  -118.926602732733,
  -117.742567054988,
  -118.893128671174,
  -119.409219751796,
  -117.519742744397,
  -118.209355279705,
  -119.321458213484,
  -119.059184510061,
  -119.409537486496,
  -118.835864687087,
  -117.901639237336,
  -118.640975252058,
  -119.668492322363,
  -117.947451962448,
  -118.311438390543,
  -118.096247909644,
  -119.670987000752,
  -117.535578262005,
  -118.188279579988,
  1,
  0,
  -118.77999384455,
  0.597531878598327,
  -119.444171737572,
  -118.963449247657,
  -118.474294970434,
  -118.991533288465,
  -120.000179864365,
  -118.263657555788,
  -118.302230887901,
  -118.920714388461,
  -118.874976020874,
  -119.425493424349,
  -119.257993988122,
  -118.591881665309,
  -117.477295944015,
  -119.690875351371,
  -118.979125957369,
  -118.440094982673,
  -118.382332777439,
  -118.227786239914,
  -118.679935830407,
  -118.211852768522,
  1,
  0,
  -118.514314191494,
  0.549712824363236,
  -118.599970472086,
  -119.057481687297,
  -118.734586262663,
  -119.658542949542,
  -117.768293872004,
  -118.680689567847,
  -117.446114901595,
  -118.222103668544,
  -118.260907380476,
  -118.90430981016,
  -119.424623039918,
  -118.287465569839,
  -118.544120754309,
  -118.868955752547,
  -117.999151448322,
  -118.702456764644,
  -118.033670366822,
  -118.26601790147,
  -117.947700250235,
  -118.879121409554,
  1,
  0,
  -118.302902202709,
  0.85222323837047,
  -118.40485913469,
  -118.926054981267,
  -116.48078575495,
  -119.51191863988,
  -118.262421315045,
  -116.990618343555,
  -116.774456272984,
  -119.183327282435,
  -118.41331499978,
  -119.293277171534,
  -118.946889288,
  -118.79597240374,
  -118.67472550089,
  -118.645149995602,
  -118.600924008301,
  -117.184009059409,
  -118.798497859739,
  -117.998073993973,
  -117.857750871158,
  -118.315017177249,
  1,
  0,
  -117.19988725228,
  0.778895292866795,
  -116.76619245982,
  -118.12902457668,
  -117.364999991965,
  -117.675099209381,
  -116.181895397036,
  -116.680884255981,
  -116.585346488696,
  -117.69374703993,
  -116.606291328067,
  -117.117284325765,
  -119.418415422647,
  -116.128824929353,
  -116.58776236468,
  -117.115124402544,
  -117.244276524863,
  -117.582652927325,
  -116.412215663626,
  -117.378779727236,
  -118.019780396367,
  -117.309147613635,
  1,
  0,
  -116.451228655988,
  0.405869576912236,
  -116.358133403866,
  -117.032752935056,
  -116.250938225785,
  -116.29340721465,
  -116.168107439689,
  -116.438361204339,
  -116.992027281778,
  -115.927255269728,
  -115.786069684397,
  -115.797927444304,
  -116.928664269133,
  -116.612580305731,
  -116.343086452031,
  -116.835210910062,
  -116.707922220026,
  -116.367632211234,
  -115.949997298092,
  -116.55081646862,
  -116.568771659833,
  -117.114911221398,
  1,
  0,
  -115.368202812258,
  0.698973251782415,
  -115.842751529936,
  -115.654144923382,
  -114.991022576047,
  -115.273888491743,
  -114.371624989026,
  -115.200691043272,
  -116.700525530866,
  -114.941559319202,
  -114.34929547719,
  -114.491646575563,
  -115.205451744322,
  -115.175083816106,
  -114.700721535957,
  -115.533291500064,
  -116.669535620639,
  -116.382471208902,
  -115.833529895747,
  -114.895418891939,
  -115.218776849833,
  -115.932624725428,
  1,
  0,
  -113.755462751562,
  0.472477096246071,
  -113.961825950532,
  -114.484668018337,
  -114.649453212647,
  -113.934013342369,
  -113.719074382452,
  -113.603545662604,
  -114.413512730542,
  -113.501923346674,
  -113.378883947971,
  -113.625154877284,
  -113.369655333962,
  -113.590730389071,
  -112.98675117764,
  -114.107453234232,
  -113.549746010361,
  -114.208233695414,
  -113.402400536231,
  -113.813342744354,
  -113.971441132608,
  -112.837445305951,
  1,
  0,
  -112.013205609684,
  0.551961068780811,
  -111.761740508453,
  -112.605653718857,
  -110.830760851179,
  -112.194145739643,
  -111.935189739238,
  -112.164257235076,
  -111.97349044422,
  -112.800928768191,
  -111.820298511049,
  -111.944037027274,
  -111.634330541436,
  -112.129147711564,
  -112.360272694065,
  -112.967789483915,
  -112.055626022441,
  -111.387823178758,
  -111.285830962761,
  -111.299673503942,
  -112.414806521022,
  -112.698309030601,
  1,
  0,
  -110.455011228269,
  0.443679508914218,
  -110.16539478463,
  -110.76875973208,
  -110.382064579965,
  -110.792243288422,
  -110.285527929471,
  -110.188191600947,
  -109.996172819792,
  -111.261397281129,
  -110.606622816034,
  -111.000496006355,
  -109.942789608982,
  -110.658128226096,
  -110.777360999583,
  -110.581179520954,
  -110.30232298607,
  -110.837237869242,
  -109.957498874029,
  -109.875410787642,
  -109.666643982562,
  -111.054780871395,
  1,
  0,
  -109.330500665604,
  0.579129386050436,
  -108.232250711232,
  -109.733518374186,
  -109.664211638909,
  -109.601658313145,
  -109.762619892202,
  -109.878209450755,
  -108.896062761215,
  -108.718790717526,
  -110.232810887819,
  -109.199051696196,
  -109.300424473454,
  -110.110939369296,
  -108.931758775719,
  -108.603716104223,
  -108.978047540008,
  -109.947171203032,
  -109.806327302531,
  -108.701851525409,
  -108.679286406979,
  -109.631306168252,
  1,
  0,
  -108.168040881831,
  0.713523300499198,
  -107.437703828902,
  -108.81826027015,
  -108.170414337147,
  -109.879336494114,
  -107.5793860684,
  -108.159473065746,
  -108.351433420446,
  -107.752404410884,
  -107.465329316214,
  -108.720729585296,
  -107.734427158852,
  -109.116738313196,
  -108.235918744025,
  -108.885455790011,
  -107.039026270377,
  -108.999532447914,
  -107.652251344627,
  -107.846339639957,
  -108.03902915656,
  -107.477627973802,
  1,
  0,
  -106.761824822801,
  0.551918208916202,
  -105.860994569044,
  -106.982411710699,
  -106.330122253614,
  -106.397685895861,
  -107.131860289388,
  -106.638636018786,
  -107.488504589659,
  -106.788628993579,
  -106.492503683379,
  -107.25260408281,
  -106.782145830903,
  -106.468430336908,
  -106.260879694927,
  -107.206005292339,
  -105.857506538515,
  -107.292027401222,
  -106.812662088947,
  -106.038572284862,
  -107.827562618465,
  -107.326752282105,
  1,
  0,
  -105.879496413021,
  0.429845672147931,
  -105.810784972569,
  -106.112268342693,
  -105.473846077056,
  -105.491486775136,
  -105.829114691921,
  -106.312612292948,
  -106.554854708657,
  -105.996276235333,
  -105.506629111696,
  -106.085887084427,
  -105.365358801442,
  -105.437699130679,
  -105.243850149487,
  -106.084422781545,
  -105.89919459257,
  -105.767529024575,
  -105.489009975729,
  -106.306393155274,
  -106.89926595522,
  -105.923444401457,
  1,
  0,
  -105.380491644572,
  0.533624773278141,
  -105.317233361763,
  -105.199229236189,
  -105.730327625948,
  -104.890898705828,
  -105.438366264276,
  -105.616737546166,
  -106.661001272152,
  -105.845632562632,
  -105.111516884324,
  -105.004260040954,
  -105.291383912625,
  -105.097190071787,
  -105.386317850597,
  -106.464711717225,
  -104.729737820085,
  -105.003049889538,
  -104.766857465231,
  -105.57424871843,
  -104.693148750817,
  -105.787983194884,
  1,
  0,
  -105.833986635796,
  0.560710791385377,
  -105.029143410722,
  -106.657603541699,
  -106.263588019496,
  -105.672903768047,
  -105.816276778085,
  -105.410359109935,
  -104.974038385059,
  -106.974948763412,
  -106.015841324867,
  -105.98817160117,
  -106.235160742077,
  -105.654627924559,
  -106.269561856411,
  -105.429512040913,
  -105.399196789993,
  -105.298548945223,
  -106.331490296996,
  -105.955249723155,
  -105.016071646332,
  -106.287438047769,
  1,
  0,
  -106.369824015592,
  0.467571019974265,
  -106.210858362546,
  -107.069666213644,
  -107.048449376215,
  -106.035710183716,
  -106.278169464949,
  -105.795505038112,
  -106.749410687956,
  -106.83712388155,
  -105.974751599278,
  -105.332509110065,
  -106.923080549206,
  -105.854798679196,
  -106.235730978685,
  -106.292662441731,
  -106.945373982735,
  -106.202316272283,
  -106.626118480865,
  -106.480500718423,
  -106.060224549878,
  -106.443519740804,
  1,
  0,
  -106.824164705793,
  0.482895364205709,
  -106.920965386545,
  -106.623037669454,
  -107.437531813254,
  -106.409765322025,
  -107.070490814486,
  -106.534359100158,
  -107.635679960242,
  -107.074652883118,
  -106.807633736052,
  -105.882097884854,
  -105.655338169935,
  -107.408065776261,
  -107.015545556151,
  -107.10533901792,
  -106.592919656904,
  -107.125471349062,
  -107.008417030866,
  -106.659518070279,
  -106.61283509431,
  -106.903629823973,
  1,
  0,
  -107.564306074419,
  0.540906657895244,
  -107.872505328686,
  -107.589275578882,
  -108.090136919086,
  -107.910364561406,
  -108.226902958671,
  -107.481932901717,
  -108.371294957176,
  -107.271143037181,
  -107.575853057148,
  -106.416040322836,
  -106.819778651567,
  -107.954034342158,
  -107.514048543463,
  -108.458897955993,
  -107.101679116092,
  -106.926694671282,
  -107.915590527477,
  -107.101473843686,
  -107.317446625502,
  -107.371027588369,
  1,
  0,
  -108.62048962358,
  0.469685019805916,
  -108.833098068361,
  -108.456247383181,
  -107.970871665594,
  -108.58330947259,
  -109.168163715104,
  -108.184699971616,
  -108.453926340622,
  -109.466318762728,
  -108.680872774665,
  -107.847475497944,
  -108.616635696167,
  -108.441492730707,
  -108.87434597975,
  -109.167230227239,
  -108.278832544007,
  -107.919109970189,
  -109.253196734774,
  -108.716612056581,
  -109.204295951461,
  -108.293056928317,
  1,
  0,
  -109.533748340344,
  0.548055843717745,
  -110.52198095849,
  -108.811132734287,
  -109.120500734571,
  -110.276256457067,
  -110.060022322005,
  -108.906208104298,
  -108.76353375555,
  -109.7977998233,
  -109.834828974754,
  -109.161350648853,
  -110.364325925745,
  -109.159269771686,
  -109.792963528101,
  -108.864683256614,
  -109.809837105282,
  -109.320069905037,
  -108.966212920198,
  -109.623444110786,
  -109.652037538438,
  -109.868508231828,
  1,
  0,
  -110.624392901088,
  0.661191681334314,
  -110.389382601986,
  -110.011078923011,
  -110.690538813621,
  -111.09974996805,
  -111.514435287596,
  -110.627270254425,
  -110.456015534694,
  -109.963164309789,
  -111.037533932896,
  -109.854602920035,
  -110.480471886173,
  -111.26232722823,
  -111.263717796816,
  -111.180091852078,
  -110.192451971937,
  -110.818096923783,
  -110.534260375579,
  -109.017272335232,
  -111.855451054871,
  -110.239944050962,
  1,
  0,
  -111.230833943846,
  0.534992180086868,
  -111.121164042562,
  -111.609690877763,
  -111.20069680179,
  -111.516715665792,
  -111.648761350766,
  -111.360823061751,
  -111.067169238176,
  -112.226408967121,
  -112.485473174969,
  -110.516082669779,
  -110.587687641111,
  -111.020553985406,
  -111.488332610237,
  -110.922502746092,
  -110.812045296116,
  -110.620744308543,
  -110.95122948177,
  -110.505293064183,
  -111.399658907583,
  -111.555644985415,
  1,
  0,
  -111.328901853732,
  0.47412714395656,
  -111.14616724221,
  -111.746291151169,
  -111.123010049831,
  -111.787822023892,
  -111.25123362636,
  -110.505224581355,
  -112.003136812273,
  -111.929483364069,
  -111.491929680466,
  -111.924358145825,
  -110.742127441448,
  -111.435955622011,
  -110.745327884063,
  -110.725591799601,
  -112.016661438112,
  -111.133868600569,
  -111.447670170731,
  -111.515835532409,
  -111.069060202013,
  -110.837281706223,
  1,
  0,
  -110.642833949014,
  0.50474156360455,
  -111.389775195513,
  -110.3153539618,
  -110.668736268515,
  -110.898337906619,
  -110.811708187257,
  -110.056640766177,
  -109.712813138879,
  -111.149474549241,
  -110.18622941581,
  -110.751234370731,
  -110.812675872776,
  -110.569323285299,
  -110.964486254849,
  -110.138754049181,
  -110.841602275296,
  -111.357608859125,
  -110.588832742834,
  -111.21059481184,
  -110.834293421261,
  -109.598203647277,
  1,
  0,
  -110.185594427494,
  0.610513193802253,
  -110.383377714865,
  -110.048910598757,
  -110.366054142714,
  -110.833326529555,
  -110.839853662714,
  -110.276246753586,
  -109.478260852936,
  -110.59202932413,
  -110.348582656181,
  -110.051394157827,
  -108.765650377954,
  -109.947222912918,
  -110.297514057615,
  -109.455972428507,
  -110.863104727223,
  -111.460056080128,
  -110.160417345793,
  -109.846780428367,
  -110.285434497542,
  -109.41169930056,
  1,
  0,
  -109.824080935962,
  0.607485570630246,
  -110.073092261915,
  -110.647052738437,
  -109.755199398227,
  -110.172382944572,
  -110.019869962522,
  -110.385458661612,
  -110.17018216521,
  -110.145512826114,
  -109.958861048149,
  -109.110386195017,
  -108.484065838535,
  -109.028940373998,
  -109.346040470671,
  -109.483864332653,
  -110.082773369637,
  -110.372749994083,
  -109.601878948531,
  -109.270955430759,
  -110.987616219971,
  -109.384735538635,
  1,
  0,
  -108.398064416704,
  0.572796873284796,
  -108.929563606923,
  -108.500085199099,
  -107.239608845619,
  -108.063725247342,
  -108.649982311191,
  -108.901833393782,
  -108.68201542247,
  -108.86251012374,
  -108.302726288484,
  -107.670105844525,
  -108.334931192364,
  -108.659944593879,
  -108.18994229482,
  -108.44752767019,
  -108.567616086113,
  -108.996336962551,
  -107.513787855772,
  -109.166174508931,
  -108.955643391201,
  -107.327227495093,
  1,
  0,
  -107.284037755274,
  0.599680269950074,
  -106.822436273788,
  -107.277927821693,
  -106.917243405496,
  -107.283461070195,
  -106.92210401737,
  -107.793738601066,
  -107.468707679567,
  -106.564312641467,
  -106.41123332957,
  -107.653598376433,
  -106.38478680584,
  -107.825202128117,
  -107.797030383436,
  -108.430497705974,
  -107.560791064236,
  -107.035741582174,
  -107.038767457816,
  -106.995223602056,
  -108.539737145126,
  -106.958214014051,
  1,
  0,
  -105.924818151284,
  0.593915272773335,
  -105.98491841126,
  -105.152905821673,
  -105.915828698132,
  -106.204273274416,
  -106.814892443734,
  -106.212902511576,
  -105.422430176453,
  -105.582345164725,
  -105.499701319857,
  -106.838497167103,
  -104.70805520106,
  -105.81366328818,
  -106.900212286386,
  -105.748012866464,
  -105.659505335718,
  -105.890980815391,
  -106.089319341374,
  -106.087907667106,
  -106.745247033528,
  -105.224764201537,
  1,
  0,
  -104.283506883483,
  0.462207936292455,
  -103.457045982256,
  -104.24379597974,
  -104.451707227594,
  -104.319253900141,
  -104.388157915852,
  -104.290971269076,
  -105.433979971283,
  -103.944271014197,
  -104.408261553939,
  -104.749526574935,
  -104.799227347265,
  -103.601451994093,
  -104.483273688245,
  -103.974905615579,
  -103.821053800996,
  -104.104882647245,
  -104.721765985257,
  -103.810769306812,
  -104.587845790068,
  -104.077990105095,
  1,
  0,
  -103.509339520928,
  0.458314267675272,
  -103.394537593655,
  -103.876800067968,
  -104.0034980398,
  -103.899489103275,
  -103.900101797756,
  -104.214515038157,
  -103.262348341103,
  -103.384886497853,
  -103.267504415128,
  -103.663584786703,
  -104.212558200077,
  -102.838059412996,
  -103.694406442808,
  -103.14476716339,
  -103.027886065694,
  -103.60073344511,
  -102.754401554258,
  -102.748241206156,
  -103.869285926284,
  -103.429185320388,
  1,
  0,
  -102.166578585361,
  0.515779319864713,
  -101.84521294551,
  -102.516614596234,
  -102.948985039314,
  -102.105901488802,
  -102.114883107631,
  -103.266322054661,
  -101.815963942551,
  -102.184945011048,
  -100.938980401225,
  -102.397153511552,
  -102.152927756622,
  -102.175091587132,
  -101.726937354634,
  -101.414853597485,
  -102.043224231212,
  -102.149987200741,
  -102.256022938557,
  -102.311483266393,
  -102.879233577997,
  -102.086848097924,
  1,
  0,
  -101.932425207852,
  0.537190449773083,
  -101.027567757834,
  -102.308899842672,
  -102.226071108571,
  -101.879425893494,
  -101.341193989036,
  -102.443621920039,
  -101.768619807385,
  -101.678468680606,
  -101.722413024511,
  -101.536553463649,
  -101.731782005627,
  -102.261625874945,
  -101.691419790379,
  -101.240042306271,
  -102.910840296335,
  -102.50965372073,
  -102.611338185204,
  -102.696069546483,
  -101.838125331791,
  -101.224771611468,
  1,
  0,
  -102.009884670576,
  0.422134025529866,
  -102.090666287306,
  -101.605695890216,
  -102.192231529091,
  -101.667799052667,
  -102.828832611251,
  -101.653305425237,
  -102.19671815897,
  -102.242973161477,
  -101.898112308273,
  -102.033853159305,
  -101.82929408005,
  -101.425294328486,
  -101.955287948471,
  -102.60260241129,
  -102.806604545042,
  -101.840862981409,
  -101.243983361315,
  -102.378527842643,
  -101.825716973728,
  -101.87933135529,
  1,
  0 ;
}
