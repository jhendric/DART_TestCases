netcdf perfect_input {
dimensions:
	member = 1 ;
	metadatalength = 32 ;
	location = 2 ;
	time = UNLIMITED ; // (1 currently)
variables:

	char MemberMetadata(member, metadatalength) ;
		MemberMetadata:long_name = "description of each member" ;

	double location(location) ;
		location:short_name = "loc1d" ;
		location:long_name = "location on a unit circle" ;
		location:dimension = 1 ;
		location:valid_range = 0., 1. ;

	double state(time, member, location) ;
		state:long_name = "the model state" ;

	double time(time) ;
		time:long_name = "valid time of the model state" ;
		time:axis = "T" ;
		time:cartesian_axis = "T" ;
		time:calendar = "none" ;
		time:units = "days" ;

// global attributes:
		:title = "true state from control" ;
                :version = "$Id: perfect_input.cdl 11431 2017-04-04 17:11:44Z hendric@ucar.edu $" ;
		:model = "ikeda" ;
		:history = "identical to original perfect_ics r2738 (circa March 2007)" ;

data:

 MemberMetadata =
  "true state" ;

 location =  0, 0.5 ;

 state = 0.136904671112630,
        -0.796420439480318 ;

 time = 124.958333333333333 ;
}
