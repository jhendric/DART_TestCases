netcdf wc13_obs {
dimensions:
	survey = 13 ;
	state_variable = 7 ;
	datum = 6815 ;
variables:
	int spherical ;
		spherical:long_name = "grid type logical switch" ;
		spherical:flag_values = 0, 1 ;
		spherical:flag_meanings = "Cartesian spherical" ;
	int Nobs(survey) ;
		Nobs:long_name = "number of observations with the same survey time" ;
	double survey_time(survey) ;
		survey_time:long_name = "survey time" ;
		survey_time:units = "days since 1968-05-23 00:00:00 GMT" ;
		survey_time:calendar = "gregorian" ;
	double obs_variance(state_variable) ;
		obs_variance:long_name = "global time and space observation variance" ;
	int obs_type(datum) ;
		obs_type:long_name = "model state variable associated with observation" ;
		obs_type:flag_values = 1, 2, 3, 4, 5, 6, 7 ;
		obs_type:flag_meanings = "zeta ubar vbar u v temperature salinity" ;
	int obs_provenance(datum) ;
		obs_provenance:long_name = "observation origin" ;
		obs_provenance:flag_values = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11 ;
		obs_provenance:flag_meanings = "gridded_AVISO_SLA blended_SST XBT_Met_Office CTD_temperature_Met_Office CTD_salinity_Met_Office ARGO_temperature_Met_Office ARGO_salinity_Met_Office CTD_temperature_CalCOFI CTD_salinity_CalCOFI CTD_temperature_GLOBEC CTD_salinity_GLOBEC" ;
	double obs_time(datum) ;
		obs_time:long_name = "time of observation" ;
		obs_time:units = "days since 1968-05-23 00:00:00 GMT" ;
		obs_time:calendar = "gregorian" ;
	double obs_depth(datum) ;
		obs_depth:long_name = "depth of observation" ;
		obs_depth:units = "meter" ;
		obs_depth:negative = "downwards" ;
	double obs_Xgrid(datum) ;
		obs_Xgrid:long_name = "observation fractional x-grid location" ;
	double obs_Ygrid(datum) ;
		obs_Ygrid:long_name = "observation fractional y-grid location" ;
	double obs_Zgrid(datum) ;
		obs_Zgrid:long_name = "observation fractional z-grid location" ;
	double obs_error(datum) ;
		obs_error:long_name = "observation error covariance" ;
	double obs_value(datum) ;
		obs_value:long_name = "observation value" ;
	double obs_lon(datum) ;
		obs_lon:long_name = "observation longitude" ;
	double obs_lat(datum) ;
		obs_lat:long_name = "observation latitude" ;

// global attributes:
		:type = "ROMS observations" ;
		:title = "California Current System, 1/3 degree resolution (WC13)" ;
		:Conventions = "CF-1.4" ;
		:grd_file = "wc13_grd.nc" ;
		:state_variables = "\n",
			"1: free-surface (m) \n",
			"2: vertically integrated u-momentum component (m/s) \n",
			"3: vertically integrated v-momentum component (m/s) \n",
			"4: u-momentum component (m/s) \n",
			"5: v-momentum component (m/s) \n",
			"6: potential temperature (Celsius) \n",
			"7: salinity (nondimensional)" ;
		:obs_provenance = "\n",
			" 1: gridded AVISO sea level anomaly \n",
			" 2: blended satellite SST \n",
			" 3: XBT temperature from Met Office \n",
			" 4: CTD temperature from Met Office \n",
			" 5: CTD salinity from Met Office \n",
			" 6: ARGO floats temperature from Met Office \n",
			" 7: ARGO floats salinity from Met Office \n",
			" 8: CTD temperature from CalCOFI \n",
			" 9: CTD salinity from CalCOFI \n",
			"10: CTD temperature from GLOBEC \n",
			"11: CTD salinity from GLOBEC " ;
		:variance_units = "squared state variable units" ;
		:obs_sources = "\n",
			"http://opendap.aviso.oceanobs.com/thredds/dodsC \n",
			"http://hadobs.metoffice.com/en3" ;
		:history = "4D-Var observations, Monday - June 21, 2010 - 11:00:00 AM" ;
		:grid_Lm_Mm_N = 54, 53, 30 ;
data:

 spherical = 1 ;

 Nobs = 1246, 38, 40, 1246, 46, 46, 1258, 27, 14, 18, 1236, 30, 1570 ;

 survey_time = 13008.5, 13008.5979166667, 13009.34375, 13009.5, 
    13009.8034722222, 13010.0548611111, 13010.5, 13010.9763888889, 
    13011.0388888889, 13011.28125, 13011.5, 13011.875, 13012 ;

 obs_variance = 0.0004, 1e-08, 1e-08, 0.01, 0.01, 0.16, 0.0001 ;

 obs_type = 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 7, 7, 7, 7, 7, 
    7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 
    7, 7, 7, 7, 7, 7, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 
    7, 7, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 7, 7, 7, 7, 
    7, 7, 7, 6, 6, 6, 6, 6, 6, 6, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    7, 7, 7, 7, 7, 7, 7, 7, 7, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 obs_provenance = 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 7, 7, 7, 
    7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 
    7, 7, 7, 7, 7, 7, 7, 7, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 
    7, 7, 7, 7, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 
    7, 7, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 
    3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 4, 4, 4, 4, 4, 4, 4, 5, 5, 
    5, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 5, 5, 5, 5, 5, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 4, 4, 4, 4, 4, 4, 4, 
    4, 4, 5, 5, 5, 5, 5, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 
    4, 4, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1 ;

 obs_time = 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5979166667, 13008.5979166667, 13008.5979166667, 13008.5979166667, 
    13008.5979166667, 13008.5979166667, 13008.5979166667, 13008.5979166667, 
    13008.5979166667, 13008.5979166667, 13008.5979166667, 13008.5979166667, 
    13008.5979166667, 13008.5979166667, 13008.5979166667, 13008.5979166667, 
    13008.5979166667, 13008.5979166667, 13008.5979166667, 13008.5979166667, 
    13008.5979166667, 13008.5979166667, 13008.5979166667, 13008.5979166667, 
    13008.5979166667, 13008.5979166667, 13008.5979166667, 13008.5979166667, 
    13008.5979166667, 13008.5979166667, 13008.5979166667, 13008.5979166667, 
    13008.5979166667, 13008.5979166667, 13008.5979166667, 13008.5979166667, 
    13008.5979166667, 13008.5979166667, 13009.34375, 13009.34375, 
    13009.34375, 13009.34375, 13009.34375, 13009.34375, 13009.34375, 
    13009.34375, 13009.34375, 13009.34375, 13009.34375, 13009.34375, 
    13009.34375, 13009.34375, 13009.34375, 13009.34375, 13009.34375, 
    13009.34375, 13009.34375, 13009.34375, 13009.34375, 13009.34375, 
    13009.34375, 13009.34375, 13009.34375, 13009.34375, 13009.34375, 
    13009.34375, 13009.34375, 13009.34375, 13009.34375, 13009.34375, 
    13009.34375, 13009.34375, 13009.34375, 13009.34375, 13009.34375, 
    13009.34375, 13009.34375, 13009.34375, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.8034722222, 13009.8034722222, 
    13009.8034722222, 13009.8034722222, 13009.8034722222, 13009.8034722222, 
    13009.8034722222, 13009.8034722222, 13009.8034722222, 13009.8034722222, 
    13009.8034722222, 13009.8034722222, 13009.8034722222, 13009.8034722222, 
    13009.8034722222, 13009.8034722222, 13009.8034722222, 13009.8034722222, 
    13009.8034722222, 13009.8034722222, 13009.8034722222, 13009.8034722222, 
    13009.8034722222, 13009.8034722222, 13009.8034722222, 13009.8034722222, 
    13009.8034722222, 13009.8034722222, 13009.8034722222, 13009.8034722222, 
    13009.8034722222, 13009.8034722222, 13009.8034722222, 13009.8034722222, 
    13009.8034722222, 13009.8034722222, 13009.8034722222, 13009.8034722222, 
    13009.8034722222, 13009.8034722222, 13009.8034722222, 13009.8034722222, 
    13009.8034722222, 13009.8034722222, 13009.8034722222, 13009.8034722222, 
    13010.0548611111, 13010.0548611111, 13010.0548611111, 13010.0548611111, 
    13010.0548611111, 13010.0548611111, 13010.0548611111, 13010.0548611111, 
    13010.0548611111, 13010.0548611111, 13010.0548611111, 13010.0548611111, 
    13010.0548611111, 13010.0548611111, 13010.0548611111, 13010.0548611111, 
    13010.0548611111, 13010.0548611111, 13010.0548611111, 13010.0548611111, 
    13010.0548611111, 13010.0548611111, 13010.0548611111, 13010.0548611111, 
    13010.0548611111, 13010.0548611111, 13010.0548611111, 13010.0548611111, 
    13010.0548611111, 13010.0548611111, 13010.0548611111, 13010.0548611111, 
    13010.0548611111, 13010.0548611111, 13010.0548611111, 13010.0548611111, 
    13010.0548611111, 13010.0548611111, 13010.0548611111, 13010.0548611111, 
    13010.0548611111, 13010.0548611111, 13010.0548611111, 13010.0548611111, 
    13010.0548611111, 13010.0548611111, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.9763888889, 
    13010.9763888889, 13010.9763888889, 13010.9763888889, 13010.9763888889, 
    13010.9763888889, 13010.9763888889, 13010.9763888889, 13010.9763888889, 
    13010.9763888889, 13010.9763888889, 13010.9763888889, 13010.9763888889, 
    13010.9763888889, 13010.9763888889, 13010.9763888889, 13010.9763888889, 
    13010.9763888889, 13010.9763888889, 13010.9763888889, 13010.9763888889, 
    13010.9763888889, 13010.9763888889, 13010.9763888889, 13010.9763888889, 
    13010.9763888889, 13010.9763888889, 13011.0388888889, 13011.0388888889, 
    13011.0388888889, 13011.0388888889, 13011.0388888889, 13011.0388888889, 
    13011.0388888889, 13011.0388888889, 13011.0388888889, 13011.0388888889, 
    13011.0388888889, 13011.0388888889, 13011.0388888889, 13011.0388888889, 
    13011.28125, 13011.28125, 13011.28125, 13011.28125, 13011.28125, 
    13011.28125, 13011.28125, 13011.28125, 13011.28125, 13011.28125, 
    13011.28125, 13011.28125, 13011.28125, 13011.28125, 13011.28125, 
    13011.28125, 13011.28125, 13011.28125, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.875, 13011.875, 13011.875, 13011.875, 13011.875, 
    13011.875, 13011.875, 13011.875, 13011.875, 13011.875, 13011.875, 
    13011.875, 13011.875, 13011.875, 13011.875, 13011.875, 13011.875, 
    13011.875, 13011.875, 13011.875, 13011.875, 13011.875, 13011.875, 
    13011.875, 13011.875, 13011.875, 13011.875, 13011.875, 13011.875, 
    13011.875, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012 ;

 obs_depth = 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 29.2668575128976, 28.2931106880205, 
    27.4265565482546, 26.5039098414807, 24.423812685455, 23.3385752962144, 
    22.4948155714326, 21.4820027503705, 19.5909409766348, 18.5006832413942, 
    17.5652301596557, 16.5915422979033, 15.5603081578148, 14.5668286869143, 
    13.5724111828824, 12.5531948612262, 11.623666106713, 25.5704522143069, 
    20.66053580274, 29.2668575128976, 28.2931106880205, 27.4265565482546, 
    26.5039098414807, 24.423812685455, 23.3385752962144, 22.4948155714326, 
    21.4820027503705, 19.5909409766348, 18.5006832413942, 17.5652301596557, 
    16.5915422979033, 15.5603081578148, 14.5668286869143, 13.5724111828824, 
    12.5531948612262, 11.623666106713, 25.5704522143069, 20.66053580274, 
    29.1765930075953, 28.2006231286159, 27.3146042719267, 26.3481835357321, 
    25.4044519671984, 24.2381525822845, 23.1385108926005, 22.2941270709058, 
    21.5922015041614, 20.7078648990055, 19.5771362306175, 18.6068110796689, 
    17.6085979442171, 16.5775260280661, 15.4903276058566, 14.4401065754562, 
    13.5199418220692, 12.5752364248567, 11.4483834094807, 10.7162619835978, 
    29.1765930075953, 28.2006231286159, 27.3146042719267, 26.3481835357321, 
    25.4044519671984, 24.2381525822845, 23.1385108926005, 22.2941270709058, 
    21.5922015041614, 20.7078648990055, 19.5771362306175, 18.6068110796689, 
    17.6085979442171, 16.5775260280661, 15.4903276058566, 14.4401065754562, 
    13.5199418220692, 12.5752364248567, 11.4483834094807, 10.7162619835978, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 28.497942925279, 26.8672133975361, 25.7129072256134, 
    24.4366222221351, 23.4392429305181, 22.6538281968931, 21.6140740635757, 
    20.478584858072, 19.4404560056958, 18.4761277049908, 17.452493216506, 
    16.4583249953704, 15.607440036457, 14.7026758073398, 13.5822394262558, 
    12.4266717533476, 11.622671244914, 10.7970234065745, 9.50682217279063, 
    8.223448811319, 7.42083701055481, 6.6473812181214, 5.92611469679479, 
    28.497942925279, 26.8672133975361, 25.7129072256134, 24.4366222221351, 
    23.4392429305181, 22.6538281968931, 21.6140740635757, 20.478584858072, 
    19.4404560056958, 18.4761277049908, 17.452493216506, 16.4583249953704, 
    15.607440036457, 14.7026758073398, 13.5822394262558, 12.4266717533476, 
    11.622671244914, 10.7970234065745, 9.50682217279063, 8.223448811319, 
    7.42083701055481, 6.6473812181214, 5.92611469679479, 29.5194516493063, 
    28.5582946049245, 27.4108598597076, 26.4988476150163, 25.7405626789316, 
    24.7425589011678, 23.542568637073, 22.4113051531266, 21.5287880368751, 
    20.4720596262526, 19.6083439038047, 18.4643809131208, 17.4508813552931, 
    16.5446768113607, 15.5292117520068, 14.5494420567707, 13.5711432106657, 
    12.5626158316309, 11.5145888879628, 10.4180809638348, 9.48128195320091, 
    8.55472553700606, 7.83020373649257, 29.5194516493063, 28.5582946049245, 
    27.4108598597076, 26.4988476150163, 25.7405626789316, 24.7425589011678, 
    23.542568637073, 22.4113051531266, 21.5287880368751, 20.4720596262526, 
    19.6083439038047, 18.4643809131208, 17.4508813552931, 16.5446768113607, 
    15.5292117520068, 14.5494420567707, 13.5711432106657, 12.5626158316309, 
    11.5145888879628, 10.4180809638348, 9.48128195320091, 8.55472553700606, 
    7.83020373649257, 14.2689979780551, 9.80039242473299, 5.43671013393478, 
    27.4934257345086, 25.0633778892587, 23.2306492782743, 21.942642182963, 
    20.959151070739, 19.6070869399149, 18.071523939678, 16.3763420228374, 
    12.1315549015429, 7.45892315102195, 3.79940525580201, 2.5300881915662, 
    1.87581273183135, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 18.4689380153097, 26.8995934164539, 24.2643706312457, 
    22.3152597273092, 20.9584439536121, 19.9255863779856, 16.7701234354496, 
    14.742514807653, 8.82349156434568, 3.73425553800546, 11.9312521281224, 
    5.93909991295722, 2.03862534607762, 12.5203876949826, 6.80019426494749, 
    2.73974882827024, 15.135895876409, 9.64929540266797, 4.50509399197809, 
    1.35111636950138, 27.0242568463261, 24.4545506234755, 22.5262260215658, 
    21.1910920075557, 20.1661447299387, 17.0699949113717, 18.7247264689812, 
    28.7161612298962, 23.6721469892783, 20.9510541403711, 17.9068920995421, 
    15.601300155688, 13.5326890324778, 11.2924797492445, 28.7161612298962, 
    23.6721469892783, 20.9510541403711, 17.9068920995421, 15.601300155688, 
    13.5326890324778, 11.2924797492445, 27.6410529895551, 22.2708069912956, 
    19.3702405519766, 17.3850930789866, 15.7910968375277, 14.2732865119821, 
    11.8926434596387, 7.25410636362123, 2.64189350702765, 27.6410529895551, 
    22.2708069912956, 19.3702405519766, 17.3850930789866, 15.7910968375277, 
    14.2732865119821, 11.8926434596387, 7.25410636362123, 2.64189350702765, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 28.7735790246829, 
    23.0855182855433, 20.506091871842, 18.7392589766159, 17.3460545527911, 
    15.0037141121633, 12.1390236056492, 7.7703533271696, 2.05406206156723, 
    28.7735790246829, 23.0855182855433, 20.506091871842, 18.7392589766159, 
    17.3460545527911, 15.0037141121633, 12.1390236056492, 7.7703533271696, 
    2.05406206156723, 27.5892905279705, 23.8945051304732, 22.4844917818553, 
    21.3376579586492, 20.4633904430287, 19.3777085361571, 17.8264841802613, 
    16.088786419746, 13.8008164291014, 11.8528899502112, 9.97484218427245, 
    7.60465261531815, 5.17551143723144, 3.3097549891584, 1.48774566301297, 
    27.5892905279705, 23.8945051304732, 22.4844917818553, 21.3376579586492, 
    20.4633904430287, 19.3777085361571, 17.8264841802613, 16.088786419746, 
    13.8008164291014, 11.8528899502112, 9.97484218427245, 7.60465261531815, 
    5.17551143723144, 3.3097549891584, 1.48774566301297, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30 ;

 obs_Xgrid = 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.8999938964843, 12.8999938964843, 12.8999938964843, 12.8999938964843, 
    12.8999938964843, 12.8999938964843, 12.8999938964843, 12.8999938964843, 
    12.8999938964843, 12.8999938964843, 12.8999938964843, 12.8999938964843, 
    12.8999938964843, 12.8999938964843, 12.8999938964843, 12.8999938964843, 
    12.8999938964843, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 14.1000061035157, 
    14.1000061035157, 14.1000061035157, 14.1000061035157, 14.1000061035157, 
    14.1000061035157, 14.1000061035157, 14.1000061035157, 14.1000061035157, 
    14.1000061035157, 14.1000061035157, 14.1000061035157, 14.1000061035157, 
    14.1000061035157, 14.1000061035157, 14.1000061035157, 14.1000061035157, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 15, 15, 15, 15, 15, 15, 15, 15, 15, 
    15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 
    15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 
    15, 15, 15, 15, 15, 15, 15.8999938964843, 15.8999938964843, 
    15.8999938964843, 15.8999938964843, 15.8999938964843, 15.8999938964843, 
    15.8999938964843, 15.8999938964843, 15.8999938964843, 15.8999938964843, 
    15.8999938964843, 15.8999938964843, 15.8999938964843, 15.8999938964843, 
    15.8999938964843, 15.8999938964843, 15.8999938964843, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 17.1000061035157, 17.1000061035157, 17.1000061035157, 
    17.1000061035157, 17.1000061035157, 17.1000061035157, 17.1000061035157, 
    17.1000061035157, 17.1000061035157, 17.1000061035157, 17.1000061035157, 
    17.1000061035157, 17.1000061035157, 17.1000061035157, 17.1000061035157, 
    17.1000061035157, 17.1000061035157, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 
    18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 
    18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 
    18.8999938964844, 18.8999938964844, 18.8999938964844, 18.8999938964844, 
    18.8999938964844, 18.8999938964844, 18.8999938964844, 18.8999938964844, 
    18.8999938964844, 18.8999938964844, 18.8999938964844, 18.8999938964844, 
    18.8999938964844, 18.8999938964844, 18.8999938964844, 18.8999938964844, 
    18.8999938964844, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 20.1000061035156, 
    20.1000061035156, 20.1000061035156, 20.1000061035156, 20.1000061035156, 
    20.1000061035156, 20.1000061035156, 20.1000061035156, 20.1000061035156, 
    20.1000061035156, 20.1000061035156, 20.1000061035156, 20.1000061035156, 
    20.1000061035156, 20.1000061035156, 20.1000061035156, 20.1000061035156, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 21, 21, 21, 21, 21, 21, 21, 21, 21, 
    21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 
    21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 
    21, 21, 21, 21, 21, 21, 21.8999938964844, 21.8999938964844, 
    21.8999938964844, 21.8999938964844, 21.8999938964844, 21.8999938964844, 
    21.8999938964844, 21.8999938964844, 21.8999938964844, 21.8999938964844, 
    21.8999938964844, 21.8999938964844, 21.8999938964844, 21.8999938964844, 
    21.8999938964844, 21.8999938964844, 21.8999938964844, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 23.1000061035156, 23.1000061035156, 23.1000061035156, 
    23.1000061035156, 23.1000061035156, 23.1000061035156, 23.1000061035156, 
    23.1000061035156, 23.1000061035156, 23.1000061035156, 23.1000061035156, 
    23.1000061035156, 23.1000061035156, 23.1000061035156, 23.1000061035156, 
    23.1000061035156, 23.1000061035156, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 
    24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 
    24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 
    24.8999938964844, 24.8999938964844, 24.8999938964844, 24.8999938964844, 
    24.8999938964844, 24.8999938964844, 24.8999938964844, 24.8999938964844, 
    24.8999938964844, 24.8999938964844, 24.8999938964844, 24.8999938964844, 
    24.8999938964844, 24.8999938964844, 24.8999938964844, 24.8999938964844, 
    24.8999938964844, 25.0499954223633, 25.0499954223633, 25.0499954223633, 
    25.0499954223633, 25.0499954223633, 25.0499954223633, 25.0499954223633, 
    25.0499954223633, 25.0499954223633, 25.0499954223633, 25.0499954223633, 
    25.0499954223633, 25.0499954223633, 25.0499954223633, 25.0499954223633, 
    25.0499954223633, 25.0499954223633, 25.0363603071733, 25.0499954223633, 
    25.1571350097656, 25.5, 25.1142817905971, 25.1399963378906, 
    25.1624965667725, 25.0499954223633, 24.75, 24.8571428571429, 
    25.0499954223633, 24.9899963378906, 25.0499954223633, 25.0363603071733, 
    25.0363603071733, 25.0090859153054, 25.0499954223633, 26.1000061035156, 
    26.1000061035156, 26.1000061035156, 26.1000061035156, 26.1000061035156, 
    26.1000061035156, 26.1000061035156, 26.1000061035156, 26.1000061035156, 
    26.1000061035156, 26.1000061035156, 26.1000061035156, 26.1000061035156, 
    26.1000061035156, 26.1000061035156, 26.1000061035156, 26.1000061035156, 
    25.9500045776367, 25.9500045776367, 25.9500045776367, 25.9500045776367, 
    25.9500045776367, 25.9500045776367, 25.9500045776367, 25.9500045776367, 
    25.9500045776367, 25.9500045776367, 25.9500045776367, 25.9500045776367, 
    25.9500045776367, 25.9500045776367, 25.9500045776367, 25.9500045776367, 
    25.9636396928267, 25.9500045776367, 25.9500045776367, 25.8600036621094, 
    26.057144165039, 25.9800064086914, 25.6000061035156, 25.7500076293945, 
    25.7625045776367, 25.9500045776367, 25.8000052315848, 26.0100036621094, 
    25.9500045776367, 25.9500045776367, 25.5750045776367, 26.040005493164, 
    27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 
    27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 26.8999938964844, 
    27, 27, 26.9499969482422, 27.0857195172991, 26.9249954223633, 
    26.7999877929688, 27.3000183105469, 27.0500030517578, 26.6999816894531, 
    27.1500091552734, 27.0600036621094, 27.1000061035156, 27, 27, 27, 
    27.0375022888184, 27, 27, 27.8999938964844, 27.8999938964844, 
    27.8999938964844, 27.8999938964844, 27.8999938964844, 27.8999938964844, 
    27.8999938964844, 27.8999938964844, 27.8999938964844, 27.8999938964844, 
    27.8999938964844, 27.8999938964844, 27.8999938964844, 27.8999938964844, 
    27.8999938964844, 27.8999938964844, 27.8999938964844, 28.0499954223633, 
    28.0499954223633, 28.0499954223633, 28.0499954223633, 28.0499954223633, 
    28.0499954223633, 28.0499954223633, 28.0499954223633, 28.0499954223633, 
    28.0499954223633, 28.0499954223633, 28.0499954223633, 28.0499954223633, 
    28.0333302815755, 28.0499954223633, 28.2, 28.0090859153054, 
    28.0333302815755, 28.1142817905971, 27.8571363176618, 27.5999908447266, 
    27.75, 28.1999931335449, 27.999994913737, 28.0999959309896, 
    28.0499954223633, 28.0499954223633, 28.0499954223633, 28.0499954223633, 
    28.0499954223633, 28.0499954223633, 29.1000061035156, 29.1000061035156, 
    29.1000061035156, 29.1000061035156, 29.1000061035156, 29.1000061035156, 
    29.1000061035156, 29.1000061035156, 29.1000061035156, 29.1000061035156, 
    29.1000061035156, 29.1000061035156, 29.1000061035156, 29.1000061035156, 
    29.1000061035156, 29.1000061035156, 29.1000061035156, 28.9500045776367, 
    28.9500045776367, 28.9500045776367, 28.9500045776367, 28.9500045776367, 
    28.9500045776367, 28.9500045776367, 28.9500045776367, 28.9500045776367, 
    28.9500045776367, 28.9500045776367, 28.9500045776367, 28.7400054931641, 
    28.8000030517578, 28.9090950705788, 28.8000052315848, 28.7571454729352, 
    29.0999908447265, 28.6000061035156, 28.8750057220459, 28.9090950705788, 
    28.9500045776367, 28.9500045776367, 28.9500045776367, 28.9500045776367, 
    28.9090950705788, 28.7625045776367, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 29.8799926757813, 29.8499908447266, 29.8499908447266, 
    29.6999816894531, 30.8999938964844, 30.8999938964844, 30.8999938964844, 
    30.8999938964844, 30.8999938964844, 30.8999938964844, 30.8999938964844, 
    30.8999938964844, 30.8999938964844, 30.8999938964844, 30.8999938964844, 
    30.8999938964844, 30.8999938964844, 30.8999938964844, 30.8999938964844, 
    30.8999938964844, 30.8999938964844, 31.0499954223633, 31.0499954223633, 
    31.0499954223633, 31.0499954223633, 31.0499954223633, 31.0499954223633, 
    31.0499954223633, 31.0090859153054, 32.1000061035156, 32.1000061035156, 
    32.1000061035156, 32.1000061035156, 32.1000061035156, 32.1000061035156, 
    32.1000061035156, 32.1000061035156, 32.1000061035156, 32.1000061035156, 
    32.1000061035156, 32.1000061035156, 32.1000061035156, 32.1000061035156, 
    32.1000061035156, 32.1000061035156, 32.1000061035156, 31.9500045776367, 
    31.9500045776367, 31.9500045776367, 31.9500045776367, 31.9500045776367, 
    31.9500045776367, 31.9500045776367, 33, 33, 33, 33, 33, 33, 33, 33, 33, 
    33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33.8999938964844, 
    33.8999938964844, 33.8999938964844, 33.8999938964844, 33.8999938964844, 
    33.8999938964844, 33.8999938964844, 33.8999938964844, 33.8999938964844, 
    33.8999938964844, 33.8999938964844, 33.8999938964844, 33.8999938964844, 
    33.8999938964844, 33.8999938964844, 33.8999938964844, 33.8999938964844, 
    34.0499954223633, 34.0499954223633, 34.0499954223633, 34.0499954223633, 
    33.959994506836, 35.1000061035156, 35.1000061035156, 35.1000061035156, 
    35.1000061035156, 35.1000061035156, 35.1000061035156, 35.1000061035156, 
    35.1000061035156, 35.1000061035156, 35.1000061035156, 35.1000061035156, 
    35.1000061035156, 35.1000061035156, 35.1000061035156, 35.1000061035156, 
    35.1000061035156, 35.1000061035156, 34.9500045776367, 34.9500045776367, 
    34.9090950705788, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 
    36, 36, 36, 35.9624977111816, 35.9624977111816, 36.8999938964844, 
    36.8999938964844, 36.8999938964844, 36.8999938964844, 36.8999938964844, 
    36.8999938964844, 36.8999938964844, 36.8999938964844, 36.8999938964844, 
    36.8999938964844, 36.8999938964844, 36.8999938964844, 36.8999938964844, 
    36.8999938964844, 36.8999938964844, 36.8999938964844, 36.8624954223633, 
    38.1000061035156, 38.1000061035156, 38.1000061035156, 38.1000061035156, 
    38.1000061035156, 38.1000061035156, 38.1000061035156, 38.1000061035156, 
    38.1000061035156, 38.1000061035156, 38.1000061035156, 38.1000061035156, 
    38.1000061035156, 38.1000061035156, 38.1000061035156, 37.9800109863281, 
    39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 
    39.8999938964844, 39.8999938964844, 39.8999938964844, 39.8999938964844, 
    39.8999938964844, 39.8999938964844, 39.8999938964844, 39.8999938964844, 
    39.8999938964844, 39.8999938964844, 39.8999938964844, 39.8999938964844, 
    39.75, 39.75, 41.1000061035156, 41.1000061035156, 41.1000061035156, 
    41.1000061035156, 41.1000061035156, 41.1000061035156, 41.1000061035156, 
    41.1000061035156, 41.1000061035156, 41.1000061035156, 41.0625057220459, 
    41.1000061035156, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 
    42.0375022888184, 42, 42.8999938964844, 42.8999938964844, 
    42.8999938964844, 42.8999938964844, 42.8999938964844, 42.8999938964844, 
    42.8999938964844, 42.8999938964844, 42.8999938964844, 42.8999938964844, 
    42.8999938964844, 42.8999938964844, 44.1000061035156, 44.1000061035156, 
    44.1000061035156, 44.1000061035156, 44.1000061035156, 44.1000061035156, 
    44.1000061035156, 44.1000061035156, 44.1000061035156, 44.1000061035156, 
    44.1000061035156, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 
    45.8999938964844, 45.8999938964844, 45.8999938964844, 45.8999938964844, 
    45.8999938964844, 45.8999938964844, 45.8999938964844, 45.8999938964844, 
    45.8999938964844, 45.8999938964844, 45.8999938964844, 47.1000061035156, 
    47.1000061035156, 47.1000061035156, 47.1000061035156, 47.1000061035156, 
    47.1000061035156, 47.1000061035156, 47.1000061035156, 47.1375045776367, 
    47.1000061035156, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48.8999938964844, 
    48.8999938964844, 48.8999938964844, 48.8999938964844, 48.8999938964844, 
    48.8999938964844, 48.8999938964844, 48.8999938964844, 48.8624954223633, 
    50.1000061035156, 50.1000061035156, 50.1000061035156, 50.1000061035156, 
    50.1000061035156, 50.1000061035156, 50.0142909458706, 49.9200073242188, 
    51, 51, 51, 51, 51, 51.8999938964844, 51.8999938964844, 51.8999938964844, 
    51.75, 17.1239776611328, 17.1239776611328, 17.1239776611328, 
    17.1239776611328, 17.1239776611328, 17.1239776611328, 17.1239776611328, 
    17.1239776611328, 17.1239776611328, 17.1239776611328, 17.1239776611328, 
    17.1239776611328, 17.1239776611328, 17.1239776611328, 17.1239776611328, 
    17.1239776611328, 17.1239776611328, 17.1239776611328, 17.1239776611328, 
    17.1239776611328, 17.1239776611328, 17.1239776611328, 17.1239776611328, 
    17.1239776611328, 17.1239776611328, 17.1239776611328, 17.1239776611328, 
    17.1239776611328, 17.1239776611328, 17.1239776611328, 17.1239776611328, 
    17.1239776611328, 17.1239776611328, 17.1239776611328, 17.1239776611328, 
    17.1239776611328, 17.1239776611328, 17.1239776611328, 20.4299926757812, 
    20.4299926757812, 20.4299926757812, 20.4299926757812, 20.4299926757812, 
    20.4299926757812, 20.4299926757812, 20.4299926757812, 20.4299926757812, 
    20.4299926757812, 20.4299926757812, 20.4299926757812, 20.4299926757812, 
    20.4299926757812, 20.4299926757812, 20.4299926757812, 20.4299926757812, 
    20.4299926757812, 20.4299926757812, 20.4299926757812, 20.4299926757812, 
    20.4299926757812, 20.4299926757812, 20.4299926757812, 20.4299926757812, 
    20.4299926757812, 20.4299926757812, 20.4299926757812, 20.4299926757812, 
    20.4299926757812, 20.4299926757812, 20.4299926757812, 20.4299926757812, 
    20.4299926757812, 20.4299926757812, 20.4299926757812, 20.4299926757812, 
    20.4299926757812, 20.4299926757812, 20.4299926757812, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.8999938964843, 12.8999938964843, 
    12.8999938964843, 12.8999938964843, 12.8999938964843, 12.8999938964843, 
    12.8999938964843, 12.8999938964843, 12.8999938964843, 12.8999938964843, 
    12.8999938964843, 12.8999938964843, 12.8999938964843, 12.8999938964843, 
    12.8999938964843, 12.8999938964843, 12.8999938964843, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 14.1000061035157, 14.1000061035157, 14.1000061035157, 
    14.1000061035157, 14.1000061035157, 14.1000061035157, 14.1000061035157, 
    14.1000061035157, 14.1000061035157, 14.1000061035157, 14.1000061035157, 
    14.1000061035157, 14.1000061035157, 14.1000061035157, 14.1000061035157, 
    14.1000061035157, 14.1000061035157, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 
    15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 
    15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 
    15.8999938964843, 15.8999938964843, 15.8999938964843, 15.8999938964843, 
    15.8999938964843, 15.8999938964843, 15.8999938964843, 15.8999938964843, 
    15.8999938964843, 15.8999938964843, 15.8999938964843, 15.8999938964843, 
    15.8999938964843, 15.8999938964843, 15.8999938964843, 15.8999938964843, 
    15.8999938964843, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 17.1000061035157, 
    17.1000061035157, 17.1000061035157, 17.1000061035157, 17.1000061035157, 
    17.1000061035157, 17.1000061035157, 17.1000061035157, 17.1000061035157, 
    17.1000061035157, 17.1000061035157, 17.1000061035157, 17.1000061035157, 
    17.1000061035157, 17.1000061035157, 17.1000061035157, 17.1000061035157, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 18, 18, 18, 18, 18, 18, 18, 18, 18, 
    18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 
    18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 
    18, 18, 18, 18, 18, 18, 18.8999938964844, 18.8999938964844, 
    18.8999938964844, 18.8999938964844, 18.8999938964844, 18.8999938964844, 
    18.8999938964844, 18.8999938964844, 18.8999938964844, 18.8999938964844, 
    18.8999938964844, 18.8999938964844, 18.8999938964844, 18.8999938964844, 
    18.8999938964844, 18.8999938964844, 18.8999938964844, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 20.1000061035156, 20.1000061035156, 20.1000061035156, 
    20.1000061035156, 20.1000061035156, 20.1000061035156, 20.1000061035156, 
    20.1000061035156, 20.1000061035156, 20.1000061035156, 20.1000061035156, 
    20.1000061035156, 20.1000061035156, 20.1000061035156, 20.1000061035156, 
    20.1000061035156, 20.1000061035156, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 
    21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 
    21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 
    21.8999938964844, 21.8999938964844, 21.8999938964844, 21.8999938964844, 
    21.8999938964844, 21.8999938964844, 21.8999938964844, 21.8999938964844, 
    21.8999938964844, 21.8999938964844, 21.8999938964844, 21.8999938964844, 
    21.8999938964844, 21.8999938964844, 21.8999938964844, 21.8999938964844, 
    21.8999938964844, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 23.1000061035156, 
    23.1000061035156, 23.1000061035156, 23.1000061035156, 23.1000061035156, 
    23.1000061035156, 23.1000061035156, 23.1000061035156, 23.1000061035156, 
    23.1000061035156, 23.1000061035156, 23.1000061035156, 23.1000061035156, 
    23.1000061035156, 23.1000061035156, 23.1000061035156, 23.1000061035156, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 24, 24, 24, 24, 24, 24, 24, 24, 24, 
    24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 
    24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 
    24, 24, 24, 24, 24, 24, 24.8999938964844, 24.8999938964844, 
    24.8999938964844, 24.8999938964844, 24.8999938964844, 24.8999938964844, 
    24.8999938964844, 24.8999938964844, 24.8999938964844, 24.8999938964844, 
    24.8999938964844, 24.8999938964844, 24.8999938964844, 24.8999938964844, 
    24.8999938964844, 24.8999938964844, 24.8999938964844, 25.0499954223633, 
    25.0499954223633, 25.0499954223633, 25.0499954223633, 25.0499954223633, 
    25.0499954223633, 25.0499954223633, 25.0499954223633, 25.0499954223633, 
    25.0499954223633, 25.0499954223633, 25.0499954223633, 25.0499954223633, 
    25.0499954223633, 25.0499954223633, 25.0499954223633, 25.0499954223633, 
    25.0363603071733, 25.0499954223633, 25.1571350097656, 25.5, 25.125, 
    25.1399963378906, 25.1624965667725, 25.0499954223633, 24.75, 
    24.8571428571429, 25.0499954223633, 24.9899963378906, 25.0499954223633, 
    25.0363603071733, 24.9899963378906, 25.0090859153054, 25.0499954223633, 
    26.1000061035156, 26.1000061035156, 26.1000061035156, 26.1000061035156, 
    26.1000061035156, 26.1000061035156, 26.1000061035156, 26.1000061035156, 
    26.1000061035156, 26.1000061035156, 26.1000061035156, 26.1000061035156, 
    26.1000061035156, 26.1000061035156, 26.1000061035156, 26.1000061035156, 
    26.1000061035156, 25.9500045776367, 25.9500045776367, 25.9500045776367, 
    25.9500045776367, 25.9500045776367, 25.9500045776367, 25.9500045776367, 
    25.9500045776367, 25.9500045776367, 25.9500045776367, 25.9500045776367, 
    25.9500045776367, 25.9500045776367, 25.9500045776367, 25.9500045776367, 
    25.9500045776367, 25.9636396928267, 25.9500045776367, 25.9500045776367, 
    25.8600036621094, 26.057144165039, 25.9800064086914, 25.6000061035156, 
    25.7500076293945, 25.7625045776367, 25.9500045776367, 25.8000052315848, 
    26.0100036621094, 25.9500045776367, 25.9500045776367, 25.6000061035156, 
    26.040005493164, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 
    27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 
    26.8799926757813, 27, 27, 26.9499969482422, 27.0857195172991, 
    26.9249954223633, 26.7999877929688, 27.3000183105469, 27.0500030517578, 
    26.6999816894531, 27.1500091552734, 27.0600036621094, 27.1000061035156, 
    27, 27, 27, 27.0375022888184, 27, 27, 27.8999938964844, 27.8999938964844, 
    27.8999938964844, 27.8999938964844, 27.8999938964844, 27.8999938964844, 
    27.8999938964844, 27.8999938964844, 27.8999938964844, 27.8999938964844, 
    27.8999938964844, 27.8999938964844, 27.8999938964844, 27.8999938964844, 
    27.8999938964844, 27.8999938964844, 27.8999938964844, 28.0499954223633, 
    28.0499954223633, 28.0499954223633, 28.0499954223633, 28.0499954223633, 
    28.0499954223633, 28.0499954223633, 28.0499954223633, 28.0499954223633, 
    28.0499954223633, 28.0499954223633, 28.0499954223633, 28.0499954223633, 
    28.0333302815755, 28.0499954223633, 28.2, 28.0090859153054, 
    28.0333302815755, 28.1142817905971, 27.8571363176618, 27.5999908447266, 
    27.75, 28.1999931335449, 27.999994913737, 28.0999959309896, 
    28.0499954223633, 28.0499954223633, 28.0499954223633, 28.0499954223633, 
    28.0499954223633, 28.0499954223633, 29.1000061035156, 29.1000061035156, 
    29.1000061035156, 29.1000061035156, 29.1000061035156, 29.1000061035156, 
    29.1000061035156, 29.1000061035156, 29.1000061035156, 29.1000061035156, 
    29.1000061035156, 29.1000061035156, 29.1000061035156, 29.1000061035156, 
    29.1000061035156, 29.1000061035156, 29.1000061035156, 28.9500045776367, 
    28.9500045776367, 28.9500045776367, 28.9500045776367, 28.9500045776367, 
    28.9500045776367, 28.9500045776367, 28.9500045776367, 28.9500045776367, 
    28.9500045776367, 28.9500045776367, 28.9500045776367, 28.7400054931641, 
    28.8000011444092, 28.9090950705788, 28.8000052315848, 28.7571454729352, 
    29.0999908447265, 28.6000061035156, 28.8750057220459, 28.9090950705788, 
    28.9500045776367, 28.9500045776367, 28.9500045776367, 28.9500045776367, 
    28.9090950705788, 28.7625045776367, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 29.8799926757813, 29.8499908447266, 29.8499908447266, 
    29.6999816894531, 30.8999938964844, 30.8999938964844, 30.8999938964844, 
    30.8999938964844, 30.8999938964844, 30.8999938964844, 30.8999938964844, 
    30.8999938964844, 30.8999938964844, 30.8999938964844, 30.8999938964844, 
    30.8999938964844, 30.8999938964844, 30.8999938964844, 30.8999938964844, 
    30.8999938964844, 30.8999938964844, 31.0499954223633, 31.0499954223633, 
    31.0499954223633, 31.0499954223633, 31.0499954223633, 31.0499954223633, 
    31.0499954223633, 31.0090859153054, 32.1000061035156, 32.1000061035156, 
    32.1000061035156, 32.1000061035156, 32.1000061035156, 32.1000061035156, 
    32.1000061035156, 32.1000061035156, 32.1000061035156, 32.1000061035156, 
    32.1000061035156, 32.1000061035156, 32.1000061035156, 32.1000061035156, 
    32.1000061035156, 32.1000061035156, 32.1000061035156, 31.9500045776367, 
    31.9500045776367, 31.9500045776367, 31.9500045776367, 31.9500045776367, 
    31.9500045776367, 31.9500045776367, 33, 33, 33, 33, 33, 33, 33, 33, 33, 
    33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33.8999938964844, 
    33.8999938964844, 33.8999938964844, 33.8999938964844, 33.8999938964844, 
    33.8999938964844, 33.8999938964844, 33.8999938964844, 33.8999938964844, 
    33.8999938964844, 33.8999938964844, 33.8999938964844, 33.8999938964844, 
    33.8999938964844, 33.8999938964844, 33.8999938964844, 33.8999938964844, 
    34.0499954223633, 34.0499954223633, 34.0499954223633, 34.0499954223633, 
    33.959994506836, 35.1000061035156, 35.1000061035156, 35.1000061035156, 
    35.1000061035156, 35.1000061035156, 35.1000061035156, 35.1000061035156, 
    35.1000061035156, 35.1000061035156, 35.1000061035156, 35.1000061035156, 
    35.1000061035156, 35.1000061035156, 35.1000061035156, 35.1000061035156, 
    35.1000061035156, 35.1000061035156, 34.9500045776367, 34.9500045776367, 
    34.9090950705788, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 
    36, 36, 36, 35.9624977111816, 35.9624977111816, 36.8999938964844, 
    36.8999938964844, 36.8999938964844, 36.8999938964844, 36.8999938964844, 
    36.8999938964844, 36.8999938964844, 36.8999938964844, 36.8999938964844, 
    36.8999938964844, 36.8999938964844, 36.8999938964844, 36.8999938964844, 
    36.8999938964844, 36.8999938964844, 36.8999938964844, 36.8624954223633, 
    38.1000061035156, 38.1000061035156, 38.1000061035156, 38.1000061035156, 
    38.1000061035156, 38.1000061035156, 38.1000061035156, 38.1000061035156, 
    38.1000061035156, 38.1000061035156, 38.1000061035156, 38.1000061035156, 
    38.1000061035156, 38.1000061035156, 38.1000061035156, 37.9800109863281, 
    39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 
    39.8999938964844, 39.8999938964844, 39.8999938964844, 39.8999938964844, 
    39.8999938964844, 39.8999938964844, 39.8999938964844, 39.8999938964844, 
    39.8999938964844, 39.8999938964844, 39.8999938964844, 39.8999938964844, 
    39.75, 39.75, 41.1000061035156, 41.1000061035156, 41.1000061035156, 
    41.1000061035156, 41.1000061035156, 41.1000061035156, 41.1000061035156, 
    41.1000061035156, 41.1000061035156, 41.1000061035156, 41.0625057220459, 
    41.1000061035156, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 
    42.0375022888184, 42, 42.8999938964844, 42.8999938964844, 
    42.8999938964844, 42.8999938964844, 42.8999938964844, 42.8999938964844, 
    42.8999938964844, 42.8999938964844, 42.8999938964844, 42.8999938964844, 
    42.8999938964844, 42.8999938964844, 44.1000061035156, 44.1000061035156, 
    44.1000061035156, 44.1000061035156, 44.1000061035156, 44.1000061035156, 
    44.1000061035156, 44.1000061035156, 44.1000061035156, 44.1000061035156, 
    44.1000061035156, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 
    45.8999938964844, 45.8999938964844, 45.8999938964844, 45.8999938964844, 
    45.8999938964844, 45.8999938964844, 45.8999938964844, 45.8999938964844, 
    45.8999938964844, 45.8999938964844, 45.8999938964844, 47.1000061035156, 
    47.1000061035156, 47.1000061035156, 47.1000061035156, 47.1000061035156, 
    47.1000061035156, 47.1000061035156, 47.1000061035156, 47.1375045776367, 
    47.1000061035156, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48.8999938964844, 
    48.8999938964844, 48.8999938964844, 48.8999938964844, 48.8999938964844, 
    48.8999938964844, 48.8999938964844, 48.8999938964844, 48.8624954223633, 
    50.1000061035156, 50.1000061035156, 50.1000061035156, 50.1000061035156, 
    50.1000061035156, 50.1000061035156, 50.0142909458706, 49.9200073242188, 
    51, 51, 51, 51, 51, 51.8999938964844, 51.8999938964844, 51.8999938964844, 
    51.75, 36.1259994506836, 36.1259994506836, 36.1259994506836, 
    36.1259994506836, 36.1259994506836, 36.1259994506836, 36.1259994506836, 
    36.1259994506836, 36.1259994506836, 36.1259994506836, 36.1259994506836, 
    36.1259994506836, 36.1259994506836, 36.1259994506836, 36.1259994506836, 
    36.1259994506836, 36.1259994506836, 36.1259994506836, 36.1259994506836, 
    36.1259994506836, 36.1259994506836, 36.1259994506836, 36.1259994506836, 
    36.1259994506836, 36.1259994506836, 36.1259994506836, 36.1259994506836, 
    36.1259994506836, 36.1259994506836, 36.1259994506836, 36.1259994506836, 
    36.1259994506836, 36.1259994506836, 36.1259994506836, 36.1259994506836, 
    36.1259994506836, 36.1259994506836, 36.1259994506836, 36.1259994506836, 
    36.1259994506836, 36.1259994506836, 36.1259994506836, 36.1259994506836, 
    36.1259994506836, 36.1259994506836, 36.1259994506836, 5.97898864746094, 
    5.97898864746094, 5.97898864746094, 5.97898864746094, 5.97898864746094, 
    5.97898864746094, 5.97898864746094, 5.97898864746094, 5.97898864746094, 
    5.97898864746094, 5.97898864746094, 5.97898864746094, 5.97898864746094, 
    5.97898864746094, 5.97898864746094, 5.97898864746094, 5.97898864746094, 
    5.97898864746094, 5.97898864746094, 5.97898864746094, 5.97898864746094, 
    5.97898864746094, 5.97898864746094, 5.97898864746094, 5.97898864746094, 
    5.97898864746094, 5.97898864746094, 5.97898864746094, 5.97898864746094, 
    5.97898864746094, 5.97898864746094, 5.97898864746094, 5.97898864746094, 
    5.97898864746094, 5.97898864746094, 5.97898864746094, 5.97898864746094, 
    5.97898864746094, 5.97898864746094, 5.97898864746094, 5.97898864746094, 
    5.97898864746094, 5.97898864746094, 5.97898864746094, 5.97898864746094, 
    5.97898864746094, 26.4090042114258, 26.4090042114258, 26.4090042114258, 
    26.4090042114258, 26.4090042114258, 26.4090042114258, 26.4090042114258, 
    26.4090042114258, 26.4090042114258, 26.4090042114258, 26.4090042114258, 
    26.4090042114258, 26.4090042114258, 26.4090042114258, 26.4090042114258, 
    26.4090042114258, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.8999938964843, 12.8999938964843, 12.8999938964843, 12.8999938964843, 
    12.8999938964843, 12.8999938964843, 12.8999938964843, 12.8999938964843, 
    12.8999938964843, 12.8999938964843, 12.8999938964843, 12.8999938964843, 
    12.8999938964843, 12.8999938964843, 12.8999938964843, 12.8999938964843, 
    12.8999938964843, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 14.1000061035157, 
    14.1000061035157, 14.1000061035157, 14.1000061035157, 14.1000061035157, 
    14.1000061035157, 14.1000061035157, 14.1000061035157, 14.1000061035157, 
    14.1000061035157, 14.1000061035157, 14.1000061035157, 14.1000061035157, 
    14.1000061035157, 14.1000061035157, 14.1000061035157, 14.1000061035157, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 15, 15, 15, 15, 15, 15, 15, 15, 15, 
    15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 
    15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 
    15, 15, 15, 15, 15, 15, 15.8999938964843, 15.8999938964843, 
    15.8999938964843, 15.8999938964843, 15.8999938964843, 15.8999938964843, 
    15.8999938964843, 15.8999938964843, 15.8999938964843, 15.8999938964843, 
    15.8999938964843, 15.8999938964843, 15.8999938964843, 15.8999938964843, 
    15.8999938964843, 15.8999938964843, 15.8999938964843, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 17.1000061035157, 17.1000061035157, 17.1000061035157, 
    17.1000061035157, 17.1000061035157, 17.1000061035157, 17.1000061035157, 
    17.1000061035157, 17.1000061035157, 17.1000061035157, 17.1000061035157, 
    17.1000061035157, 17.1000061035157, 17.1000061035157, 17.1000061035157, 
    17.1000061035157, 17.1000061035157, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 
    18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 
    18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 
    18.8999938964844, 18.8999938964844, 18.8999938964844, 18.8999938964844, 
    18.8999938964844, 18.8999938964844, 18.8999938964844, 18.8999938964844, 
    18.8999938964844, 18.8999938964844, 18.8999938964844, 18.8999938964844, 
    18.8999938964844, 18.8999938964844, 18.8999938964844, 18.8999938964844, 
    18.8999938964844, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 20.1000061035156, 
    20.1000061035156, 20.1000061035156, 20.1000061035156, 20.1000061035156, 
    20.1000061035156, 20.1000061035156, 20.1000061035156, 20.1000061035156, 
    20.1000061035156, 20.1000061035156, 20.1000061035156, 20.1000061035156, 
    20.1000061035156, 20.1000061035156, 20.1000061035156, 20.1000061035156, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 21, 21, 21, 21, 21, 21, 21, 21, 21, 
    21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 
    21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 
    21, 21, 21, 21, 21, 21, 21.8999938964844, 21.8999938964844, 
    21.8999938964844, 21.8999938964844, 21.8999938964844, 21.8999938964844, 
    21.8999938964844, 21.8999938964844, 21.8999938964844, 21.8999938964844, 
    21.8999938964844, 21.8999938964844, 21.8999938964844, 21.8999938964844, 
    21.8999938964844, 21.8999938964844, 21.8999938964844, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 23.1000061035156, 23.1000061035156, 23.1000061035156, 
    23.1000061035156, 23.1000061035156, 23.1000061035156, 23.1000061035156, 
    23.1000061035156, 23.1000061035156, 23.1000061035156, 23.1000061035156, 
    23.1000061035156, 23.1000061035156, 23.1000061035156, 23.1000061035156, 
    23.1000061035156, 23.1000061035156, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 
    24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 
    24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 
    24.8999938964844, 24.8999938964844, 24.8999938964844, 24.8999938964844, 
    24.8999938964844, 24.8999938964844, 24.8999938964844, 24.8999938964844, 
    24.8999938964844, 24.8999938964844, 24.8999938964844, 24.8999938964844, 
    24.8999938964844, 24.8999938964844, 24.8999938964844, 24.8999938964844, 
    24.8999938964844, 25.0499954223633, 25.0499954223633, 25.0499954223633, 
    25.0499954223633, 25.0499954223633, 25.0499954223633, 25.0499954223633, 
    25.0499954223633, 25.0499954223633, 25.0499954223633, 25.0499954223633, 
    25.0499954223633, 25.0499954223633, 25.0499954223633, 25.0499954223633, 
    25.0499954223633, 25.0499954223633, 24.9333292643229, 25.0499954223633, 
    25.1999931335449, 25.125, 25.3499908447266, 25.1142817905971, 
    25.0499954223633, 24.75, 24.8571428571429, 24.9899963378906, 
    25.0090859153054, 25.0499954223633, 25.0363603071733, 24.9899963378906, 
    25.0090859153054, 25.0499954223633, 26.1000061035156, 26.1000061035156, 
    26.1000061035156, 26.1000061035156, 26.1000061035156, 26.1000061035156, 
    26.1000061035156, 26.1000061035156, 26.1000061035156, 26.1000061035156, 
    26.1000061035156, 26.1000061035156, 26.1000061035156, 26.1000061035156, 
    26.1000061035156, 26.1000061035156, 26.1000061035156, 25.9500045776367, 
    25.9500045776367, 25.9500045776367, 25.9500045776367, 25.9500045776367, 
    25.9500045776367, 25.9500045776367, 25.9500045776367, 25.9500045776367, 
    25.9500045776367, 25.9500045776367, 25.9500045776367, 25.9500045776367, 
    25.9500045776367, 25.9500045776367, 25.9500045776367, 25.9636396928267, 
    26.0666707356771, 25.9500045776367, 25.8600036621094, 26.1500015258789, 
    25.9800064086914, 25.5, 25.5, 25.7625045776367, 25.6500091552734, 
    25.8500061035156, 26.0100036621094, 25.9500045776367, 25.9500045776367, 
    25.6000061035156, 26.040005493164, 27, 27, 27, 27, 27, 27, 27, 27, 27, 
    27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 
    27, 27, 27, 27, 27, 26.7749862670898, 26.6999816894531, 26.9499969482422, 
    27.1000061035156, 27.0857195172991, 26.9249954223633, 26.7999877929688, 
    27.3000183105469, 27, 26.6999816894531, 27.1500091552734, 27, 
    27.1000061035156, 27, 27, 27, 27, 27, 27, 27.8999938964844, 
    27.8999938964844, 27.8999938964844, 27.8999938964844, 27.8999938964844, 
    27.8999938964844, 27.8999938964844, 27.8999938964844, 27.8999938964844, 
    27.8999938964844, 27.8999938964844, 27.8999938964844, 27.8999938964844, 
    27.8999938964844, 27.8999938964844, 27.8999938964844, 27.8999938964844, 
    28.0499954223633, 28.0499954223633, 28.0499954223633, 28.0499954223633, 
    28.0499954223633, 28.0499954223633, 28.0499954223633, 28.0499954223633, 
    28.0499954223633, 28.0499954223633, 28.0499954223633, 28.0499954223633, 
    28.0636305375533, 28.0333302815755, 28.079997253418, 28.5, 
    27.959994506836, 27.8999938964844, 27.8249931335449, 27.5999908447266, 
    27.75, 28.0499954223633, 28.0499954223633, 28.0999959309896, 
    28.0499954223633, 28.0499954223633, 28.0499954223633, 28.0499954223633, 
    28.0499954223633, 28.0499954223633, 29.1000061035156, 29.1000061035156, 
    29.1000061035156, 29.1000061035156, 29.1000061035156, 29.1000061035156, 
    29.1000061035156, 29.1000061035156, 29.1000061035156, 29.1000061035156, 
    29.1000061035156, 29.1000061035156, 29.1000061035156, 29.1000061035156, 
    29.1000061035156, 29.1000061035156, 29.1000061035156, 28.9500045776367, 
    28.9500045776367, 28.9500045776367, 28.9500045776367, 28.9500045776367, 
    28.9500045776367, 28.9500045776367, 28.9500045776367, 28.9500045776367, 
    28.9500045776367, 28.9500045776367, 28.9500045776367, 28.7400054931641, 
    28.8000011444092, 29.000005086263, 28.9500045776367, 28.6500091552734, 
    28.8750057220459, 28.9090950705788, 28.9500045776367, 28.9500045776367, 
    28.9500045776367, 28.9500045776367, 28.9090950705788, 28.7625045776367, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 29.8799926757813, 
    29.8499908447266, 29.8499908447266, 29.6999816894531, 30.8999938964844, 
    30.8999938964844, 30.8999938964844, 30.8999938964844, 30.8999938964844, 
    30.8999938964844, 30.8999938964844, 30.8999938964844, 30.8999938964844, 
    30.8999938964844, 30.8999938964844, 30.8999938964844, 30.8999938964844, 
    30.8999938964844, 30.8999938964844, 30.8999938964844, 30.8999938964844, 
    31.0499954223633, 31.0499954223633, 31.0499954223633, 31.0499954223633, 
    31.0499954223633, 31.0499954223633, 31.0499954223633, 31.0090859153054, 
    32.1000061035156, 32.1000061035156, 32.1000061035156, 32.1000061035156, 
    32.1000061035156, 32.1000061035156, 32.1000061035156, 32.1000061035156, 
    32.1000061035156, 32.1000061035156, 32.1000061035156, 32.1000061035156, 
    32.1000061035156, 32.1000061035156, 32.1000061035156, 32.1000061035156, 
    32.1000061035156, 31.9500045776367, 31.9500045776367, 31.9500045776367, 
    31.9500045776367, 31.9500045776367, 31.9500045776367, 31.9500045776367, 
    33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 
    33, 33, 33, 33, 33.8999938964844, 33.8999938964844, 33.8999938964844, 
    33.8999938964844, 33.8999938964844, 33.8999938964844, 33.8999938964844, 
    33.8999938964844, 33.8999938964844, 33.8999938964844, 33.8999938964844, 
    33.8999938964844, 33.8999938964844, 33.8999938964844, 33.8999938964844, 
    33.8999938964844, 33.8999938964844, 34.0499954223633, 34.0499954223633, 
    34.0499954223633, 34.0499954223633, 33.959994506836, 35.1000061035156, 
    35.1000061035156, 35.1000061035156, 35.1000061035156, 35.1000061035156, 
    35.1000061035156, 35.1000061035156, 35.1000061035156, 35.1000061035156, 
    35.1000061035156, 35.1000061035156, 35.1000061035156, 35.1000061035156, 
    35.1000061035156, 35.1000061035156, 35.1000061035156, 35.1000061035156, 
    34.9500045776367, 34.9500045776367, 34.9090950705788, 36, 36, 36, 36, 36, 
    36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 35.9624977111816, 
    35.9624977111816, 36.8999938964844, 36.8999938964844, 36.8999938964844, 
    36.8999938964844, 36.8999938964844, 36.8999938964844, 36.8999938964844, 
    36.8999938964844, 36.8999938964844, 36.8999938964844, 36.8999938964844, 
    36.8999938964844, 36.8999938964844, 36.8999938964844, 36.8999938964844, 
    36.8999938964844, 36.8624954223633, 38.1000061035156, 38.1000061035156, 
    38.1000061035156, 38.1000061035156, 38.1000061035156, 38.1000061035156, 
    38.1000061035156, 38.1000061035156, 38.1000061035156, 38.1000061035156, 
    38.1000061035156, 38.1000061035156, 38.1000061035156, 38.1000061035156, 
    38.1000061035156, 37.9800109863281, 39, 39, 39, 39, 39, 39, 39, 39, 39, 
    39, 39, 39, 39, 39, 39, 39.8999938964844, 39.8999938964844, 
    39.8999938964844, 39.8999938964844, 39.8999938964844, 39.8999938964844, 
    39.8999938964844, 39.8999938964844, 39.8999938964844, 39.8999938964844, 
    39.8999938964844, 39.8999938964844, 39.75, 39.75, 41.1000061035156, 
    41.1000061035156, 41.1000061035156, 41.1000061035156, 41.1000061035156, 
    41.1000061035156, 41.1000061035156, 41.1000061035156, 41.1000061035156, 
    41.1000061035156, 41.0625057220459, 41.1000061035156, 42, 42, 42, 42, 42, 
    42, 42, 42, 42, 42, 42.0375022888184, 42, 42.8999938964844, 
    42.8999938964844, 42.8999938964844, 42.8999938964844, 42.8999938964844, 
    42.8999938964844, 42.8999938964844, 42.8999938964844, 42.8999938964844, 
    42.8999938964844, 42.8999938964844, 42.8999938964844, 44.1000061035156, 
    44.1000061035156, 44.1000061035156, 44.1000061035156, 44.1000061035156, 
    44.1000061035156, 44.1000061035156, 44.1000061035156, 44.1000061035156, 
    44.1000061035156, 44.1000061035156, 45, 45, 45, 45, 45, 45, 45, 45, 45, 
    45, 45, 45.8999938964844, 45.8999938964844, 45.8999938964844, 
    45.8999938964844, 45.8999938964844, 45.8999938964844, 45.8999938964844, 
    45.8999938964844, 45.8999938964844, 45.8999938964844, 45.8999938964844, 
    47.1000061035156, 47.1000061035156, 47.1000061035156, 47.1000061035156, 
    47.1000061035156, 47.1000061035156, 47.1000061035156, 47.1000061035156, 
    47.1375045776367, 47.1000061035156, 48, 48, 48, 48, 48, 48, 48, 48, 48, 
    48.8999938964844, 48.8999938964844, 48.8999938964844, 48.8999938964844, 
    48.8999938964844, 48.8999938964844, 48.8999938964844, 48.8999938964844, 
    48.8624954223633, 50.1000061035156, 50.1000061035156, 50.1000061035156, 
    50.1000061035156, 50.1000061035156, 50.1000061035156, 50.0142909458706, 
    49.9200073242188, 51, 51, 51, 51, 51, 51.8999938964844, 51.8999938964844, 
    51.8999938964844, 51.75, 27.5969924926758, 27.5969924926758, 
    27.5969924926758, 27.5969924926758, 27.5969924926758, 27.5969924926758, 
    27.5969924926758, 27.5969924926758, 27.5969924926758, 27.5969924926758, 
    27.5969924926758, 27.5969924926758, 27.5969924926758, 27.7830047607422, 
    27.7830047607422, 27.7830047607422, 27.7830047607422, 27.7830047607422, 
    27.7830047607422, 27.7830047607422, 27.7830047607422, 27.7830047607422, 
    27.7830047607422, 27.7830047607422, 27.7830047607422, 27.7830047607422, 
    27.7830047607422, 50.0909957885742, 50.0909957885742, 50.0909957885742, 
    50.0909957885742, 50.0909957885742, 50.0909957885742, 50.0909957885742, 
    50.0909957885742, 50.0909957885742, 50.0909957885742, 50.0909957885742, 
    50.0909957885742, 50.0909957885742, 50.0909957885742, 49.754997253418, 
    49.754997253418, 49.754997253418, 49.754997253418, 49.754997253418, 
    49.754997253418, 49.754997253418, 49.754997253418, 49.754997253418, 
    49.754997253418, 49.754997253418, 49.754997253418, 49.754997253418, 
    49.754997253418, 49.754997253418, 49.754997253418, 49.754997253418, 
    49.754997253418, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.8999938964843, 12.8999938964843, 12.8999938964843, 12.8999938964843, 
    12.8999938964843, 12.8999938964843, 12.8999938964843, 12.8999938964843, 
    12.8999938964843, 12.8999938964843, 12.8999938964843, 12.8999938964843, 
    12.8999938964843, 12.8999938964843, 12.8999938964843, 12.8999938964843, 
    12.8999938964843, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 14.1000061035157, 
    14.1000061035157, 14.1000061035157, 14.1000061035157, 14.1000061035157, 
    14.1000061035157, 14.1000061035157, 14.1000061035157, 14.1000061035157, 
    14.1000061035157, 14.1000061035157, 14.1000061035157, 14.1000061035157, 
    14.1000061035157, 14.1000061035157, 14.1000061035157, 14.1000061035157, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 15, 15, 15, 15, 15, 15, 15, 15, 15, 
    15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 
    15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 
    15, 15, 15, 15, 15, 15, 15.8999938964843, 15.8999938964843, 
    15.8999938964843, 15.8999938964843, 15.8999938964843, 15.8999938964843, 
    15.8999938964843, 15.8999938964843, 15.8999938964843, 15.8999938964843, 
    15.8999938964843, 15.8999938964843, 15.8999938964843, 15.8999938964843, 
    15.8999938964843, 15.8999938964843, 15.8999938964843, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 17.1000061035157, 17.1000061035157, 17.1000061035157, 
    17.1000061035157, 17.1000061035157, 17.1000061035157, 17.1000061035157, 
    17.1000061035157, 17.1000061035157, 17.1000061035157, 17.1000061035157, 
    17.1000061035157, 17.1000061035157, 17.1000061035157, 17.1000061035157, 
    17.1000061035157, 17.1000061035157, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 
    18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 
    18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 
    18.8999938964844, 18.8999938964844, 18.8999938964844, 18.8999938964844, 
    18.8999938964844, 18.8999938964844, 18.8999938964844, 18.8999938964844, 
    18.8999938964844, 18.8999938964844, 18.8999938964844, 18.8999938964844, 
    18.8999938964844, 18.8999938964844, 18.8999938964844, 18.8999938964844, 
    18.8999938964844, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 20.1000061035156, 
    20.1000061035156, 20.1000061035156, 20.1000061035156, 20.1000061035156, 
    20.1000061035156, 20.1000061035156, 20.1000061035156, 20.1000061035156, 
    20.1000061035156, 20.1000061035156, 20.1000061035156, 20.1000061035156, 
    20.1000061035156, 20.1000061035156, 20.1000061035156, 20.1000061035156, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 21, 21, 21, 21, 21, 21, 21, 21, 21, 
    21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 
    21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 
    21, 21, 21, 21, 21, 21, 21.8999938964844, 21.8999938964844, 
    21.8999938964844, 21.8999938964844, 21.8999938964844, 21.8999938964844, 
    21.8999938964844, 21.8999938964844, 21.8999938964844, 21.8999938964844, 
    21.8999938964844, 21.8999938964844, 21.8999938964844, 21.8999938964844, 
    21.8999938964844, 21.8999938964844, 21.8999938964844, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 23.1000061035156, 23.1000061035156, 23.1000061035156, 
    23.1000061035156, 23.1000061035156, 23.1000061035156, 23.1000061035156, 
    23.1000061035156, 23.1000061035156, 23.1000061035156, 23.1000061035156, 
    23.1000061035156, 23.1000061035156, 23.1000061035156, 23.1000061035156, 
    23.1000061035156, 23.1000061035156, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 
    24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 
    24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 
    24.8999938964844, 24.8999938964844, 24.8999938964844, 24.8999938964844, 
    24.8999938964844, 24.8999938964844, 24.8999938964844, 24.8999938964844, 
    24.8999938964844, 24.8999938964844, 24.8999938964844, 24.8999938964844, 
    24.8999938964844, 24.8999938964844, 24.8999938964844, 24.8999938964844, 
    24.8999938964844, 25.0499954223633, 25.0499954223633, 25.0499954223633, 
    25.0499954223633, 25.0499954223633, 25.0499954223633, 25.0499954223633, 
    25.0499954223633, 25.0499954223633, 25.0499954223633, 25.0363603071733, 
    25.0499954223633, 25.0363603071733, 25.0499954223633, 25.0090859153054, 
    25.0499954223633, 25.0363603071733, 24.942855834961, 25.0499954223633, 
    25.5, 24.75, 24.959994506836, 24.8999977111817, 24.9333292643229, 
    25.0363603071733, 25.0499954223633, 25.0499954223633, 25.0499954223633, 
    25.0499954223633, 25.0499954223633, 26.1000061035156, 26.1000061035156, 
    26.1000061035156, 26.1000061035156, 26.1000061035156, 26.1000061035156, 
    26.1000061035156, 26.1000061035156, 26.1000061035156, 26.1000061035156, 
    26.1000061035156, 26.1000061035156, 26.1000061035156, 26.1000061035156, 
    26.1000061035156, 26.1000061035156, 26.1000061035156, 25.9500045776367, 
    25.9500045776367, 25.9500045776367, 25.9500045776367, 25.9500045776367, 
    25.9500045776367, 25.9500045776367, 25.9500045776367, 25.9500045776367, 
    25.9500045776367, 25.9090950705788, 25.9500045776367, 25.9500045776367, 
    25.9636396928267, 25.8, 25.8000052315848, 25.9125022888183, 
    25.7000122070312, 25.9666697184245, 25.6500091552734, 25.8000068664551, 
    25.9500045776367, 26.0250091552734, 25.9800018310547, 25.9500045776367, 
    25.9500045776367, 25.9500045776367, 25.9500045776367, 25.9500045776367, 
    27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 
    27, 27, 27, 27, 27, 27, 27, 27, 27, 26.9624977111816, 27, 
    26.9142804827009, 26.8799926757813, 26.6999816894531, 26.6999816894531, 
    27, 27.1000061035156, 27, 27, 27, 27, 27, 26.9624977111816, 
    27.8999938964844, 27.8999938964844, 27.8999938964844, 27.8999938964844, 
    27.8999938964844, 27.8999938964844, 27.8999938964844, 27.8999938964844, 
    27.8999938964844, 27.8999938964844, 27.8999938964844, 27.8999938964844, 
    27.8999938964844, 27.8999938964844, 27.8999938964844, 27.8999938964844, 
    27.8999938964844, 28.0499954223633, 28.0499954223633, 28.0499954223633, 
    28.0499954223633, 28.0499954223633, 28.0499954223633, 28.0499954223633, 
    28.0499954223633, 28.0499954223633, 28.0499954223633, 28.0909049294212, 
    28.0090859153054, 28.0874977111817, 28.079997253418, 28.5, 
    27.5999908447266, 28.0499954223633, 28.109994506836, 28.0499954223633, 
    28.0499954223633, 28.0499954223633, 28.0499954223633, 28.0499954223633, 
    28.0499954223633, 29.1000061035156, 29.1000061035156, 29.1000061035156, 
    29.1000061035156, 29.1000061035156, 29.1000061035156, 29.1000061035156, 
    29.1000061035156, 29.1000061035156, 29.1000061035156, 29.1000061035156, 
    29.1000061035156, 29.1000061035156, 29.1000061035156, 29.1000061035156, 
    29.1000061035156, 29.1000061035156, 28.9500045776367, 28.9500045776367, 
    28.9500045776367, 28.9500045776367, 28.9500045776367, 28.9500045776367, 
    28.9500045776367, 28.9500045776367, 28.9500045776367, 28.9500045776367, 
    28.9500045776367, 28.8857182094029, 28.7400054931641, 28.7000045776367, 
    28.5, 28.8750057220459, 28.9090950705788, 28.9500045776367, 
    28.9500045776367, 28.9500045776367, 28.9500045776367, 28.9090950705788, 
    28.7625045776367, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 29.8799926757813, 
    29.8499908447266, 29.8499908447266, 29.6999816894531, 30.8999938964844, 
    30.8999938964844, 30.8999938964844, 30.8999938964844, 30.8999938964844, 
    30.8999938964844, 30.8999938964844, 30.8999938964844, 30.8999938964844, 
    30.8999938964844, 30.8999938964844, 30.8999938964844, 30.8999938964844, 
    30.8999938964844, 30.8999938964844, 30.8999938964844, 30.8999938964844, 
    31.0499954223633, 31.0499954223633, 31.0499954223633, 31.0499954223633, 
    31.0499954223633, 31.0499954223633, 31.0499954223633, 31.0090859153054, 
    32.1000061035156, 32.1000061035156, 32.1000061035156, 32.1000061035156, 
    32.1000061035156, 32.1000061035156, 32.1000061035156, 32.1000061035156, 
    32.1000061035156, 32.1000061035156, 32.1000061035156, 32.1000061035156, 
    32.1000061035156, 32.1000061035156, 32.1000061035156, 32.1000061035156, 
    32.1000061035156, 31.9500045776367, 31.9500045776367, 31.9500045776367, 
    31.9500045776367, 31.9500045776367, 31.9500045776367, 31.9500045776367, 
    33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 
    33, 33, 33, 33, 33.8999938964844, 33.8999938964844, 33.8999938964844, 
    33.8999938964844, 33.8999938964844, 33.8999938964844, 33.8999938964844, 
    33.8999938964844, 33.8999938964844, 33.8999938964844, 33.8999938964844, 
    33.8999938964844, 33.8999938964844, 33.8999938964844, 33.8999938964844, 
    33.8999938964844, 33.8999938964844, 34.0499954223633, 34.0499954223633, 
    34.0499954223633, 34.0499954223633, 33.8999938964844, 35.1000061035156, 
    35.1000061035156, 35.1000061035156, 35.1000061035156, 35.1000061035156, 
    35.1000061035156, 35.1000061035156, 35.1000061035156, 35.1000061035156, 
    35.1000061035156, 35.1000061035156, 35.1000061035156, 35.1000061035156, 
    35.1000061035156, 35.1000061035156, 35.1000061035156, 35.1000061035156, 
    34.9500045776367, 34.9500045776367, 34.9090950705788, 36, 36, 36, 36, 36, 
    36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 35.9624977111816, 
    35.9624977111816, 36.8999938964844, 36.8999938964844, 36.8999938964844, 
    36.8999938964844, 36.8999938964844, 36.8999938964844, 36.8999938964844, 
    36.8999938964844, 36.8999938964844, 36.8999938964844, 36.8999938964844, 
    36.8999938964844, 36.8999938964844, 36.8999938964844, 36.8999938964844, 
    36.8999938964844, 36.8624954223633, 38.1000061035156, 38.1000061035156, 
    38.1000061035156, 38.1000061035156, 38.1000061035156, 38.1000061035156, 
    38.1000061035156, 38.1000061035156, 38.1000061035156, 38.1000061035156, 
    38.1000061035156, 38.1000061035156, 38.1000061035156, 38.1000061035156, 
    38.1000061035156, 37.9800109863281, 39, 39, 39, 39, 39, 39, 39, 39, 39, 
    39, 39, 39, 39, 39, 39, 39.8999938964844, 39.8999938964844, 
    39.8999938964844, 39.8999938964844, 39.8999938964844, 39.8999938964844, 
    39.8999938964844, 39.8999938964844, 39.8999938964844, 39.8999938964844, 
    39.8999938964844, 39.8999938964844, 39.75, 39.75, 41.1000061035156, 
    41.1000061035156, 41.1000061035156, 41.1000061035156, 41.1000061035156, 
    41.1000061035156, 41.1000061035156, 41.1000061035156, 41.1000061035156, 
    41.1000061035156, 41.0625057220459, 41.1000061035156, 42, 42, 42, 42, 42, 
    42, 42, 42, 42, 42, 42.0375022888184, 42, 42.8999938964844, 
    42.8999938964844, 42.8999938964844, 42.8999938964844, 42.8999938964844, 
    42.8999938964844, 42.8999938964844, 42.8999938964844, 42.8999938964844, 
    42.8999938964844, 42.8999938964844, 42.8999938964844, 44.1000061035156, 
    44.1000061035156, 44.1000061035156, 44.1000061035156, 44.1000061035156, 
    44.1000061035156, 44.1000061035156, 44.1000061035156, 44.1000061035156, 
    44.1000061035156, 44.1000061035156, 45, 45, 45, 45, 45, 45, 45, 45, 45, 
    45, 45, 45.8999938964844, 45.8999938964844, 45.8999938964844, 
    45.8999938964844, 45.8999938964844, 45.8999938964844, 45.8999938964844, 
    45.8999938964844, 45.8999938964844, 45.8999938964844, 45.8999938964844, 
    47.1000061035156, 47.1000061035156, 47.1000061035156, 47.1000061035156, 
    47.1000061035156, 47.1000061035156, 47.1000061035156, 47.1000061035156, 
    47.1375045776367, 47.1000061035156, 48, 48, 48, 48, 48, 48, 48, 48, 48, 
    48.8999938964844, 48.8999938964844, 48.8999938964844, 48.8999938964844, 
    48.8999938964844, 48.8999938964844, 48.8999938964844, 48.8999938964844, 
    48.8624954223633, 50.1000061035156, 50.1000061035156, 50.1000061035156, 
    50.1000061035156, 50.1000061035156, 50.1000061035156, 50.0142909458706, 
    49.9200073242188, 51, 51, 51, 51, 51, 51.8999938964844, 51.8999938964844, 
    51.8999938964844, 51.75, 48.375, 48.375, 48.375, 48.375, 48.375, 48.375, 
    48.375, 48.375, 48.375, 48.375, 48.375, 48.375, 48.375, 48.375, 48.375, 
    48.375, 48.375, 48.375, 46.343994140625, 46.343994140625, 
    46.343994140625, 46.343994140625, 46.343994140625, 46.343994140625, 
    46.343994140625, 46.343994140625, 46.343994140625, 46.343994140625, 
    46.343994140625, 46.343994140625, 46.343994140625, 46.343994140625, 
    46.343994140625, 46.343994140625, 46.343994140625, 46.343994140625, 
    46.343994140625, 46.343994140625, 46.343994140625, 46.343994140625, 
    46.343994140625, 46.343994140625, 46.343994140625, 46.343994140625, 
    46.343994140625, 46.343994140625, 46.343994140625, 46.343994140625, 
    2.99999999993187, 3.99999999993179, 2.99999999993187, 4.9999999999317, 
    3.99999999993179, 5.99999999993162, 4.9999999999317, 6.99999999993145, 
    5.99999999993162, 2.99999999993187, 7.99999999993145, 6.99999999993145, 
    3.99999999993179, 8.99999999993127, 2.99999999993187, 7.99999999993145, 
    4.9999999999317, 9.99999999993119, 3.99999999993179, 8.99999999993128, 
    5.99999999993162, 2.99999999993187, 10.9999999999311, 4.9999999999317, 
    9.99999999993119, 6.99999999993145, 3.99999999993179, 11.999999999931, 
    5.99999999993162, 2.99999999993187, 10.9999999999311, 7.99999999993145, 
    4.9999999999317, 12.9999999999308, 6.99999999993145, 3.99999999993179, 
    11.999999999931, 8.99999999993128, 5.99999999993162, 13.9999999999308, 
    2.99999999993187, 7.99999999993145, 4.9999999999317, 12.9999999999308, 
    9.99999999993119, 6.99999999993145, 14.9999999999307, 3.99999999993179, 
    8.99999999993128, 5.99999999993162, 13.9999999999308, 2.99999999993187, 
    10.9999999999311, 7.99999999993145, 15.9999999999306, 4.9999999999317, 
    9.99999999993119, 6.99999999993145, 14.9999999999307, 3.99999999993179, 
    11.999999999931, 8.99999999993128, 16.9999999999305, 5.99999999993162, 
    2.99999999993187, 10.9999999999311, 7.99999999993145, 15.9999999999306, 
    4.9999999999317, 12.9999999999309, 9.99999999993119, 17.9999999999304, 
    6.99999999993145, 3.99999999993179, 11.999999999931, 8.99999999993128, 
    16.9999999999305, 5.99999999993162, 13.9999999999308, 2.99999999993187, 
    10.9999999999311, 18.9999999999303, 7.99999999993145, 4.9999999999317, 
    12.9999999999308, 9.99999999993119, 17.9999999999304, 6.99999999993145, 
    14.9999999999307, 3.99999999993179, 11.999999999931, 19.9999999999302, 
    8.99999999993128, 5.99999999993162, 13.9999999999308, 2.99999999993187, 
    10.9999999999311, 18.9999999999303, 7.99999999993145, 15.9999999999306, 
    4.9999999999317, 12.9999999999308, 20.9999999999301, 9.99999999993119, 
    6.99999999993145, 14.9999999999307, 3.99999999993179, 11.999999999931, 
    19.9999999999302, 8.99999999993127, 16.9999999999305, 5.99999999993162, 
    13.9999999999308, 21.99999999993, 2.99999999993187, 10.9999999999311, 
    7.99999999993145, 15.9999999999306, 4.9999999999317, 12.9999999999308, 
    20.9999999999301, 9.99999999993119, 17.9999999999304, 6.99999999993145, 
    14.9999999999307, 22.9999999999299, 3.99999999993179, 11.999999999931, 
    8.99999999993128, 16.9999999999305, 5.99999999993162, 13.9999999999308, 
    21.99999999993, 2.99999999993187, 10.9999999999311, 18.9999999999303, 
    7.99999999993145, 15.9999999999306, 23.9999999999298, 4.9999999999317, 
    12.9999999999308, 9.99999999993119, 17.9999999999304, 6.99999999993145, 
    14.9999999999307, 22.9999999999299, 3.99999999993179, 11.999999999931, 
    19.9999999999302, 8.99999999993127, 16.9999999999305, 24.9999999999297, 
    5.99999999993162, 13.9999999999308, 2.99999999993187, 10.9999999999311, 
    18.9999999999303, 7.99999999993145, 15.9999999999306, 23.9999999999298, 
    4.9999999999317, 12.9999999999308, 20.9999999999301, 9.99999999993119, 
    17.9999999999304, 25.9999999999296, 6.99999999993145, 14.9999999999307, 
    3.99999999993179, 11.999999999931, 19.9999999999302, 8.99999999993128, 
    16.9999999999305, 24.9999999999297, 5.99999999993162, 13.9999999999308, 
    21.99999999993, 2.99999999993187, 10.9999999999311, 18.9999999999303, 
    26.9999999999295, 7.99999999993145, 15.9999999999306, 4.9999999999317, 
    12.9999999999308, 20.9999999999301, 9.99999999993119, 17.9999999999304, 
    25.9999999999296, 6.99999999993145, 14.9999999999307, 22.9999999999299, 
    3.99999999993179, 11.999999999931, 19.9999999999302, 27.9999999999294, 
    8.99999999993128, 16.9999999999305, 5.99999999993162, 13.9999999999309, 
    21.99999999993, 2.99999999993187, 10.9999999999311, 18.9999999999303, 
    26.9999999999295, 7.99999999993145, 15.9999999999306, 23.9999999999298, 
    4.9999999999317, 12.9999999999308, 20.9999999999301, 28.9999999999293, 
    9.99999999993119, 17.9999999999304, 6.99999999993145, 14.9999999999307, 
    22.9999999999299, 3.99999999993179, 11.999999999931, 19.9999999999302, 
    27.9999999999294, 8.99999999993128, 16.9999999999305, 24.9999999999297, 
    5.99999999993162, 13.9999999999308, 21.99999999993, 2.99999999993187, 
    29.9999999999292, 10.9999999999311, 18.9999999999303, 7.99999999993145, 
    15.9999999999306, 23.9999999999298, 4.9999999999317, 12.9999999999308, 
    20.9999999999301, 28.9999999999293, 9.99999999993119, 17.9999999999304, 
    25.9999999999296, 6.99999999993145, 14.9999999999307, 22.9999999999299, 
    3.99999999993179, 30.9999999999291, 11.999999999931, 19.9999999999302, 
    8.99999999993128, 16.9999999999305, 24.9999999999297, 5.99999999993162, 
    13.9999999999308, 21.99999999993, 2.99999999993187, 29.9999999999292, 
    10.9999999999311, 18.9999999999303, 26.9999999999295, 7.99999999993145, 
    15.9999999999306, 23.9999999999298, 4.9999999999317, 31.999999999929, 
    12.9999999999308, 20.9999999999301, 9.99999999993119, 17.9999999999304, 
    25.9999999999296, 6.99999999993145, 14.9999999999307, 22.9999999999299, 
    3.99999999993179, 30.9999999999291, 11.999999999931, 19.9999999999302, 
    27.9999999999294, 8.99999999993128, 16.9999999999305, 24.9999999999297, 
    5.99999999993162, 32.9999999999289, 13.9999999999308, 21.99999999993, 
    2.99999999993187, 10.9999999999311, 18.9999999999303, 26.9999999999295, 
    7.99999999993145, 15.9999999999306, 23.9999999999298, 4.9999999999317, 
    31.999999999929, 12.9999999999309, 20.9999999999301, 28.9999999999293, 
    9.99999999993119, 17.9999999999304, 25.9999999999296, 6.99999999993145, 
    33.9999999999288, 14.9999999999307, 22.9999999999299, 3.99999999993179, 
    11.999999999931, 19.9999999999302, 27.9999999999294, 8.99999999993128, 
    16.9999999999305, 24.9999999999297, 5.99999999993162, 32.9999999999289, 
    13.9999999999308, 21.99999999993, 2.99999999993187, 29.9999999999292, 
    10.9999999999311, 18.9999999999303, 26.9999999999295, 7.99999999993145, 
    34.9999999999287, 15.9999999999306, 23.9999999999298, 4.9999999999317, 
    12.9999999999308, 20.9999999999301, 28.9999999999293, 9.99999999993119, 
    17.9999999999304, 25.9999999999296, 6.99999999993145, 33.9999999999288, 
    14.9999999999307, 22.9999999999299, 3.99999999993179, 30.9999999999291, 
    11.999999999931, 19.9999999999302, 27.9999999999294, 8.99999999993128, 
    35.9999999999286, 16.9999999999305, 24.9999999999297, 5.99999999993162, 
    13.9999999999308, 21.99999999993, 2.99999999993187, 29.9999999999292, 
    10.9999999999311, 18.9999999999303, 26.9999999999295, 7.99999999993145, 
    34.9999999999287, 15.9999999999306, 23.9999999999298, 4.9999999999317, 
    31.999999999929, 12.9999999999308, 20.9999999999301, 28.9999999999293, 
    9.99999999993119, 36.9999999999285, 17.9999999999304, 25.9999999999296, 
    6.99999999993145, 14.9999999999307, 22.9999999999299, 3.99999999993179, 
    30.9999999999291, 11.999999999931, 19.9999999999302, 27.9999999999294, 
    8.99999999993127, 35.9999999999286, 16.9999999999305, 24.9999999999297, 
    5.99999999993162, 32.9999999999289, 13.9999999999308, 21.99999999993, 
    2.99999999993187, 29.9999999999292, 10.9999999999311, 37.9999999999284, 
    18.9999999999303, 26.9999999999295, 7.99999999993145, 15.9999999999306, 
    23.9999999999298, 4.9999999999317, 31.999999999929, 12.9999999999308, 
    20.9999999999301, 28.9999999999293, 9.99999999993119, 36.9999999999285, 
    17.9999999999304, 25.9999999999296, 6.99999999993145, 33.9999999999288, 
    14.9999999999307, 22.9999999999299, 3.99999999993179, 30.9999999999291, 
    11.999999999931, 38.9999999999283, 19.9999999999302, 27.9999999999294, 
    8.99999999993128, 16.9999999999305, 24.9999999999297, 5.99999999993162, 
    32.9999999999289, 13.9999999999308, 21.99999999993, 2.99999999993187, 
    29.9999999999292, 10.9999999999311, 37.9999999999284, 18.9999999999303, 
    26.9999999999295, 7.99999999993145, 34.9999999999287, 15.9999999999306, 
    23.9999999999298, 4.9999999999317, 31.999999999929, 12.9999999999309, 
    39.9999999999283, 20.9999999999301, 28.9999999999293, 9.99999999993119, 
    17.9999999999304, 25.9999999999296, 6.99999999993145, 33.9999999999288, 
    14.9999999999307, 22.9999999999299, 3.99999999993179, 30.9999999999291, 
    11.999999999931, 38.9999999999283, 19.9999999999302, 27.9999999999294, 
    8.99999999993128, 35.9999999999286, 16.9999999999305, 24.9999999999297, 
    5.99999999993162, 32.9999999999289, 13.9999999999309, 40.9999999999281, 
    21.99999999993, 2.99999999993187, 29.9999999999292, 10.9999999999311, 
    18.9999999999303, 26.9999999999295, 7.99999999993145, 34.9999999999287, 
    15.9999999999306, 23.9999999999298, 4.9999999999317, 31.999999999929, 
    12.9999999999308, 39.9999999999282, 20.9999999999301, 28.9999999999293, 
    9.99999999993119, 36.9999999999285, 17.9999999999304, 25.9999999999296, 
    6.99999999993145, 33.9999999999288, 14.9999999999307, 41.999999999928, 
    22.9999999999299, 3.99999999993179, 30.9999999999291, 11.999999999931, 
    19.9999999999302, 27.9999999999294, 8.99999999993128, 35.9999999999286, 
    16.9999999999305, 24.9999999999297, 5.99999999993162, 32.9999999999289, 
    13.9999999999309, 40.9999999999281, 21.99999999993, 2.99999999993187, 
    29.9999999999292, 10.9999999999311, 37.9999999999284, 18.9999999999303, 
    26.9999999999295, 7.99999999993145, 34.9999999999287, 15.9999999999306, 
    42.9999999999279, 23.9999999999298, 4.9999999999317, 31.999999999929, 
    12.9999999999308, 20.9999999999301, 28.9999999999293, 9.99999999993119, 
    36.9999999999285, 17.9999999999304, 25.9999999999296, 6.99999999993145, 
    33.9999999999288, 14.9999999999307, 41.999999999928, 22.9999999999299, 
    3.99999999993179, 30.9999999999291, 11.999999999931, 38.9999999999283, 
    19.9999999999302, 27.9999999999294, 8.99999999993128, 35.9999999999286, 
    16.9999999999305, 43.9999999999278, 24.9999999999297, 5.99999999993162, 
    32.9999999999289, 13.9999999999308, 21.99999999993, 2.99999999993187, 
    29.9999999999292, 10.9999999999311, 37.9999999999284, 18.9999999999303, 
    26.9999999999295, 7.99999999993145, 34.9999999999287, 15.9999999999306, 
    42.9999999999279, 23.9999999999298, 4.9999999999317, 31.999999999929, 
    12.9999999999308, 39.9999999999282, 20.9999999999301, 28.9999999999293, 
    9.99999999993119, 36.9999999999285, 17.9999999999304, 44.9999999999277, 
    25.9999999999296, 6.99999999993145, 33.9999999999288, 14.9999999999307, 
    22.9999999999299, 3.99999999993179, 30.9999999999291, 11.999999999931, 
    38.9999999999283, 19.9999999999302, 27.9999999999294, 8.99999999993127, 
    35.9999999999286, 16.9999999999305, 43.9999999999278, 24.9999999999297, 
    5.99999999993162, 32.9999999999289, 13.9999999999308, 40.9999999999281, 
    21.99999999993, 2.99999999993187, 29.9999999999292, 10.9999999999311, 
    37.9999999999284, 18.9999999999303, 45.9999999999277, 26.9999999999295, 
    7.99999999993145, 34.9999999999287, 15.9999999999306, 23.9999999999298, 
    4.9999999999317, 31.999999999929, 12.9999999999308, 39.9999999999282, 
    20.9999999999301, 28.9999999999293, 9.99999999993119, 36.9999999999285, 
    17.9999999999304, 44.9999999999277, 25.9999999999296, 6.99999999993145, 
    33.9999999999288, 14.9999999999307, 41.999999999928, 22.9999999999299, 
    3.99999999993179, 30.9999999999291, 11.999999999931, 38.9999999999283, 
    19.9999999999302, 46.9999999999275, 27.9999999999294, 8.99999999993128, 
    35.9999999999286, 16.9999999999305, 24.9999999999297, 5.99999999993162, 
    32.9999999999289, 13.9999999999308, 40.9999999999281, 21.99999999993, 
    2.99999999993187, 29.9999999999292, 10.9999999999311, 37.9999999999284, 
    18.9999999999303, 45.9999999999277, 26.9999999999295, 7.99999999993145, 
    34.9999999999287, 15.9999999999306, 42.9999999999279, 23.9999999999298, 
    4.9999999999317, 31.999999999929, 12.9999999999308, 39.9999999999282, 
    20.9999999999301, 47.9999999999274, 28.9999999999293, 9.99999999993119, 
    36.9999999999285, 17.9999999999304, 25.9999999999296, 6.99999999993145, 
    33.9999999999288, 14.9999999999307, 41.999999999928, 22.9999999999299, 
    3.99999999993179, 30.9999999999291, 11.999999999931, 38.9999999999283, 
    19.9999999999302, 46.9999999999275, 27.9999999999294, 8.99999999993128, 
    35.9999999999286, 16.9999999999305, 43.9999999999278, 24.9999999999297, 
    5.99999999993162, 32.9999999999289, 13.9999999999308, 40.9999999999281, 
    21.99999999993, 2.99999999993187, 48.9999999999273, 29.9999999999292, 
    10.9999999999311, 37.9999999999284, 18.9999999999303, 26.9999999999295, 
    7.99999999993145, 34.9999999999287, 15.9999999999306, 42.9999999999279, 
    23.9999999999298, 4.9999999999317, 31.999999999929, 12.9999999999308, 
    39.9999999999282, 20.9999999999301, 47.9999999999274, 28.9999999999293, 
    9.99999999993119, 36.9999999999285, 17.9999999999304, 44.9999999999277, 
    25.9999999999296, 6.99999999993145, 33.9999999999288, 14.9999999999307, 
    41.999999999928, 22.9999999999299, 3.99999999993179, 49.9999999999273, 
    30.9999999999291, 11.999999999931, 38.9999999999283, 19.9999999999302, 
    27.9999999999294, 8.99999999993128, 35.9999999999286, 16.9999999999305, 
    43.9999999999278, 24.9999999999297, 5.99999999993162, 32.9999999999289, 
    13.9999999999308, 40.9999999999281, 21.99999999993, 2.99999999993187, 
    48.9999999999273, 29.9999999999292, 10.9999999999311, 37.9999999999284, 
    18.9999999999303, 45.9999999999277, 26.9999999999295, 7.99999999993145, 
    34.9999999999287, 15.9999999999306, 42.9999999999279, 23.9999999999298, 
    4.9999999999317, 50.9999999999271, 31.999999999929, 12.9999999999308, 
    39.9999999999282, 20.9999999999301, 28.9999999999293, 9.99999999993119, 
    36.9999999999285, 17.9999999999304, 44.9999999999277, 25.9999999999296, 
    6.99999999993145, 33.9999999999288, 14.9999999999307, 41.999999999928, 
    22.9999999999299, 3.99999999993179, 49.9999999999273, 30.9999999999291, 
    11.999999999931, 38.9999999999283, 19.9999999999302, 46.9999999999275, 
    27.9999999999294, 8.99999999993128, 35.9999999999286, 16.9999999999305, 
    43.9999999999278, 24.9999999999297, 5.99999999993162, 51.9999999999271, 
    32.9999999999289, 13.9999999999309, 40.9999999999281, 21.99999999993, 
    2.99999999993187, 29.9999999999292, 10.9999999999311, 37.9999999999284, 
    18.9999999999303, 45.9999999999277, 26.9999999999295, 7.99999999993145, 
    34.9999999999287, 15.9999999999306, 42.9999999999279, 23.9999999999298, 
    4.9999999999317, 50.9999999999271, 31.999999999929, 12.9999999999308, 
    39.9999999999282, 20.9999999999301, 47.9999999999274, 28.9999999999293, 
    9.99999999993119, 36.9999999999285, 17.9999999999304, 44.9999999999277, 
    25.9999999999296, 6.99999999993145, 33.9999999999288, 14.9999999999307, 
    41.999999999928, 22.9999999999299, 3.99999999993179, 30.9999999999291, 
    11.999999999931, 38.9999999999283, 19.9999999999302, 46.9999999999275, 
    27.9999999999294, 8.99999999993128, 35.9999999999286, 16.9999999999305, 
    43.9999999999278, 24.9999999999297, 5.99999999993162, 51.9999999999271, 
    32.9999999999289, 13.9999999999309, 40.9999999999281, 21.99999999993, 
    2.99999999993187, 48.9999999999273, 29.9999999999292, 10.9999999999311, 
    37.9999999999284, 18.9999999999303, 45.9999999999277, 26.9999999999295, 
    7.99999999993145, 34.9999999999287, 15.9999999999306, 42.9999999999279, 
    23.9999999999298, 4.9999999999317, 31.999999999929, 12.9999999999308, 
    39.9999999999282, 20.9999999999301, 47.9999999999274, 28.9999999999293, 
    9.99999999993119, 36.9999999999285, 17.9999999999304, 44.9999999999277, 
    25.9999999999296, 6.99999999993145, 33.9999999999288, 14.9999999999307, 
    41.999999999928, 22.9999999999299, 3.99999999993179, 49.9999999999273, 
    30.9999999999291, 11.999999999931, 38.9999999999283, 19.9999999999302, 
    46.9999999999275, 27.9999999999294, 8.99999999993128, 35.9999999999286, 
    16.9999999999305, 43.9999999999278, 24.9999999999297, 5.99999999993162, 
    32.9999999999289, 13.9999999999308, 40.9999999999281, 21.99999999993, 
    2.99999999993187, 48.9999999999273, 29.9999999999292, 10.9999999999311, 
    37.9999999999284, 18.9999999999303, 45.9999999999277, 26.9999999999295, 
    7.99999999993145, 34.9999999999287, 15.9999999999306, 42.9999999999279, 
    23.9999999999298, 4.9999999999317, 50.9999999999271, 31.999999999929, 
    12.9999999999308, 39.9999999999282, 20.9999999999301, 47.9999999999274, 
    28.9999999999293, 9.99999999993119, 36.9999999999285, 17.9999999999304, 
    44.9999999999277, 25.9999999999296, 6.99999999993145, 33.9999999999288, 
    14.9999999999307, 41.999999999928, 22.9999999999299, 3.99999999993179, 
    49.9999999999273, 30.9999999999291, 11.999999999931, 38.9999999999283, 
    19.9999999999302, 46.9999999999275, 27.9999999999294, 8.99999999993128, 
    35.9999999999286, 16.9999999999305, 43.9999999999278, 24.9999999999297, 
    5.99999999993162, 32.9999999999289, 13.9999999999308, 40.9999999999281, 
    21.99999999993, 2.99999999993187, 48.9999999999273, 29.9999999999292, 
    10.9999999999311, 37.9999999999284, 18.9999999999303, 45.9999999999277, 
    26.9999999999295, 7.99999999993145, 34.9999999999287, 15.9999999999306, 
    42.9999999999279, 23.9999999999298, 4.9999999999317, 31.999999999929, 
    12.9999999999308, 39.9999999999282, 20.9999999999301, 28.9999999999293, 
    9.99999999993119, 36.9999999999285, 17.9999999999304, 44.9999999999277, 
    25.9999999999296, 6.99999999993145, 33.9999999999288, 14.9999999999307, 
    41.999999999928, 22.9999999999299, 3.99999999993179, 49.9999999999273, 
    30.9999999999291, 11.999999999931, 38.9999999999283, 19.9999999999302, 
    46.9999999999275, 27.9999999999294, 8.99999999993128, 35.9999999999286, 
    16.9999999999305, 24.9999999999297, 5.99999999993162, 32.9999999999289, 
    13.9999999999308, 21.99999999993, 2.99999999993187, 29.9999999999292, 
    10.9999999999311, 37.9999999999284, 18.9999999999303, 45.9999999999276, 
    26.9999999999295, 7.99999999993145, 34.9999999999287, 15.9999999999306, 
    42.9999999999279, 23.9999999999298, 4.9999999999317, 31.999999999929, 
    12.9999999999309, 39.9999999999282, 20.9999999999301, 28.9999999999293, 
    9.99999999993119, 36.9999999999285, 17.9999999999304, 25.9999999999296, 
    6.99999999993145, 33.9999999999288, 14.9999999999307, 22.9999999999299, 
    3.99999999993179, 30.9999999999291, 11.999999999931, 38.9999999999283, 
    19.9999999999302, 46.9999999999275, 27.9999999999294, 8.99999999993128, 
    35.9999999999286, 16.9999999999305, 24.9999999999297, 5.99999999993162, 
    32.9999999999289, 13.9999999999309, 21.99999999993, 2.99999999993187, 
    29.9999999999292, 10.9999999999311, 37.9999999999284, 18.9999999999303, 
    26.9999999999295, 7.99999999993145, 34.9999999999287, 15.9999999999306, 
    23.9999999999298, 4.9999999999317, 31.999999999929, 12.9999999999308, 
    20.9999999999301, 28.9999999999293, 9.99999999993119, 36.9999999999285, 
    17.9999999999304, 25.9999999999296, 6.99999999993145, 33.9999999999288, 
    14.9999999999307, 22.9999999999299, 3.99999999993179, 30.9999999999291, 
    11.999999999931, 19.9999999999302, 27.9999999999294, 8.99999999993128, 
    35.9999999999286, 16.9999999999305, 24.9999999999297, 5.99999999993162, 
    32.9999999999289, 13.9999999999308, 21.99999999993, 2.99999999993187, 
    29.9999999999292, 10.9999999999311, 18.9999999999303, 26.9999999999295, 
    7.99999999993145, 34.9999999999287, 15.9999999999306, 23.9999999999298, 
    4.9999999999317, 31.999999999929, 12.9999999999308, 20.9999999999301, 
    28.9999999999293, 9.99999999993119, 17.9999999999304, 25.9999999999296, 
    6.99999999993145, 33.9999999999288, 14.9999999999307, 22.9999999999299, 
    3.99999999993179, 30.9999999999291, 11.999999999931, 19.9999999999302, 
    27.9999999999294, 8.99999999993128, 35.9999999999286, 16.9999999999305, 
    24.9999999999297, 5.99999999993162, 32.9999999999289, 13.9999999999309, 
    21.99999999993, 2.99999999993187, 29.9999999999292, 10.9999999999311, 
    18.9999999999303, 26.9999999999295, 7.99999999993145, 34.9999999999287, 
    15.9999999999306, 23.9999999999298, 4.9999999999317, 31.999999999929, 
    12.9999999999308, 20.9999999999301, 28.9999999999293, 9.99999999993119, 
    17.9999999999304, 25.9999999999296, 6.99999999993145, 33.9999999999288, 
    14.9999999999307, 22.9999999999299, 3.99999999993179, 30.9999999999291, 
    11.999999999931, 19.9999999999302, 27.9999999999294, 8.99999999993128, 
    16.9999999999305, 24.9999999999297, 5.99999999993162, 32.9999999999289, 
    13.9999999999308, 21.99999999993, 2.99999999993187, 29.9999999999292, 
    10.9999999999311, 18.9999999999303, 26.9999999999295, 7.99999999993145, 
    15.9999999999306, 23.9999999999298, 4.9999999999317, 31.999999999929, 
    12.9999999999308, 20.9999999999301, 28.9999999999293, 9.99999999993119, 
    17.9999999999304, 25.9999999999296, 6.99999999993145, 33.9999999999288, 
    14.9999999999307, 22.9999999999299, 3.99999999993179, 30.9999999999291, 
    11.999999999931, 19.9999999999302, 27.9999999999294, 8.99999999993128, 
    16.9999999999305, 24.9999999999297, 5.99999999993162, 13.9999999999308, 
    21.99999999993, 2.99999999993187, 29.9999999999292, 10.9999999999311, 
    18.9999999999303, 26.9999999999295, 7.99999999993145, 15.9999999999306, 
    23.9999999999298, 4.9999999999317, 12.9999999999308, 20.9999999999301, 
    28.9999999999293, 9.99999999993119, 17.9999999999304, 25.9999999999296, 
    6.99999999993145, 14.9999999999307, 22.9999999999299, 3.99999999993179, 
    30.9999999999291, 11.999999999931, 19.9999999999302, 27.9999999999294, 
    8.99999999993128, 16.9999999999305, 24.9999999999297, 5.99999999993162, 
    13.9999999999308, 21.99999999993, 2.99999999993187, 29.9999999999292, 
    10.9999999999311, 18.9999999999303, 26.9999999999295, 7.99999999993145, 
    15.9999999999306, 23.9999999999298, 4.9999999999317, 12.9999999999308, 
    20.9999999999301, 28.9999999999293, 9.99999999993119, 17.9999999999304, 
    25.9999999999296, 6.99999999993145, 14.9999999999307, 22.9999999999299, 
    3.99999999993179, 11.999999999931, 19.9999999999302, 27.9999999999294, 
    8.99999999993128, 16.9999999999305, 24.9999999999297, 5.99999999993162, 
    13.9999999999308, 21.99999999993, 2.99999999993187, 29.9999999999292, 
    10.9999999999311, 18.9999999999303, 26.9999999999295, 7.99999999993145, 
    15.9999999999306, 23.9999999999298, 4.9999999999317, 12.9999999999308, 
    20.9999999999301, 28.9999999999293, 9.99999999993119, 17.9999999999304, 
    25.9999999999296, 6.99999999993145, 14.9999999999307, 22.9999999999299, 
    3.99999999993179, 11.999999999931, 19.9999999999302, 27.9999999999294, 
    8.99999999993127, 16.9999999999305, 24.9999999999297, 5.99999999993162, 
    13.9999999999308, 21.99999999993, 2.99999999993187, 29.9999999999292, 
    10.9999999999311, 18.9999999999303, 26.9999999999295, 7.99999999993145, 
    15.9999999999306, 23.9999999999298, 4.9999999999317, 12.9999999999308, 
    20.9999999999301, 28.9999999999293, 9.99999999993119, 17.9999999999304, 
    25.9999999999296, 6.99999999993145, 14.9999999999307, 22.9999999999299, 
    3.99999999993179, 11.999999999931, 19.9999999999302, 27.9999999999294, 
    8.99999999993128, 16.9999999999305, 24.9999999999297, 5.99999999993162, 
    13.9999999999309, 21.99999999993, 2.99999999993187, 10.9999999999311, 
    18.9999999999303, 26.9999999999295, 7.99999999993145, 15.9999999999306, 
    23.9999999999298, 4.9999999999317, 12.9999999999308, 20.9999999999301, 
    9.99999999993119, 17.9999999999304, 25.9999999999296, 6.99999999993145, 
    14.9999999999307, 22.9999999999299, 3.99999999993179, 11.999999999931, 
    19.9999999999302, 27.9999999999294, 8.99999999993128, 16.9999999999305, 
    24.9999999999297, 5.99999999993162, 13.9999999999308, 21.99999999993, 
    2.99999999993187, 10.9999999999311, 18.9999999999303, 26.9999999999295, 
    7.99999999993145, 15.9999999999306, 23.9999999999298, 4.9999999999317, 
    12.9999999999308, 20.9999999999301, 28.9999999999293, 9.99999999993119, 
    17.9999999999304, 25.9999999999296, 6.99999999993145, 14.9999999999307, 
    22.9999999999299, 3.99999999993179, 11.999999999931, 19.9999999999302, 
    27.9999999999294, 8.99999999993128, 16.9999999999305, 24.9999999999297, 
    5.99999999993162, 13.9999999999308, 21.99999999993, 2.99999999993187, 
    10.9999999999311, 18.9999999999303, 26.9999999999295, 7.99999999993145, 
    15.9999999999306, 23.9999999999298, 4.9999999999317, 12.9999999999308, 
    20.9999999999301, 28.9999999999293, 9.99999999993119, 17.9999999999304, 
    25.9999999999296, 6.99999999993145, 14.9999999999307, 22.9999999999299, 
    3.99999999993179, 11.999999999931, 19.9999999999302, 8.99999999993128, 
    16.9999999999305, 24.9999999999297, 5.99999999993162, 13.9999999999308, 
    21.99999999993, 2.99999999993187, 10.9999999999311, 18.9999999999303, 
    26.9999999999295, 7.99999999993145, 15.9999999999306, 23.9999999999298, 
    4.9999999999317, 12.9999999999308, 20.9999999999301, 9.99999999993119, 
    17.9999999999304, 25.9999999999296, 6.99999999993145, 14.9999999999307, 
    22.9999999999299, 3.99999999993179, 11.999999999931, 19.9999999999302, 
    8.99999999993128, 16.9999999999305, 24.9999999999297, 5.99999999993162, 
    13.9999999999308, 21.99999999993, 2.99999999993187, 10.9999999999311, 
    18.9999999999303, 26.9999999999295, 7.99999999993145, 15.9999999999306, 
    23.9999999999298, 4.9999999999317, 12.9999999999308, 20.9999999999301, 
    9.99999999993119, 17.9999999999304, 25.9999999999296, 6.99999999993145, 
    14.9999999999307, 22.9999999999299, 3.99999999993179, 11.999999999931, 
    19.9999999999302, 8.99999999993128, 16.9999999999305, 24.9999999999297, 
    5.99999999993162, 13.9999999999308, 21.99999999993, 10.9999999999311, 
    18.9999999999303, 26.9999999999295, 7.99999999993145, 15.9999999999306, 
    23.9999999999298, 4.9999999999317, 12.9999999999308, 20.9999999999301, 
    9.99999999993119, 17.9999999999304, 25.9999999999296, 6.99999999993145, 
    14.9999999999307, 22.9999999999299, 11.999999999931, 19.9999999999302, 
    27.9999999999294, 8.99999999993127, 16.9999999999305, 24.9999999999297, 
    5.99999999993162, 13.9999999999309, 21.99999999993, 10.9999999999311, 
    18.9999999999303, 26.9999999999295, 7.99999999993145, 15.9999999999306, 
    23.9999999999298, 12.9999999999308, 20.9999999999301, 9.99999999993119, 
    17.9999999999304, 25.9999999999296, 6.99999999993145, 14.9999999999307, 
    22.9999999999299, 11.999999999931, 19.9999999999302, 27.9999999999294, 
    8.99999999993128, 16.9999999999305, 24.9999999999297, 13.9999999999308, 
    21.99999999993, 10.9999999999311, 18.9999999999303, 26.9999999999295, 
    7.99999999993145, 15.9999999999306, 23.9999999999298, 12.9999999999309, 
    20.9999999999301, 9.99999999993119, 17.9999999999304, 25.9999999999296, 
    14.9999999999307, 22.9999999999299, 11.999999999931, 19.9999999999302, 
    27.9999999999294, 8.99999999993128, 16.9999999999305, 24.9999999999297, 
    13.9999999999308, 21.99999999993, 10.9999999999311, 18.9999999999303, 
    26.9999999999295, 15.9999999999306, 23.9999999999298, 12.9999999999308, 
    20.9999999999301, 9.99999999993119, 17.9999999999304, 25.9999999999296, 
    14.9999999999307, 22.9999999999299, 11.999999999931, 19.9999999999302, 
    27.9999999999294, 16.9999999999305, 24.9999999999297, 13.9999999999309, 
    21.99999999993, 10.9999999999311, 18.9999999999303, 26.9999999999295, 
    15.9999999999306, 23.9999999999298, 12.9999999999309, 20.9999999999301, 
    17.9999999999304, 25.9999999999296, 14.9999999999307, 22.9999999999299, 
    11.999999999931, 19.9999999999302, 27.9999999999294, 16.9999999999305, 
    24.9999999999297, 13.9999999999308, 21.99999999993, 18.9999999999303, 
    26.9999999999295, 15.9999999999306, 23.9999999999298, 12.9999999999308, 
    20.9999999999301, 28.9999999999293, 17.9999999999304, 25.9999999999296, 
    14.9999999999307, 22.9999999999299, 19.9999999999302, 27.9999999999294, 
    16.9999999999305, 24.9999999999297, 13.9999999999308, 21.99999999993, 
    18.9999999999303, 26.9999999999295, 15.9999999999306, 23.9999999999298, 
    20.9999999999301, 28.9999999999293, 17.9999999999304, 25.9999999999296, 
    14.9999999999307, 22.9999999999299, 19.9999999999302, 27.9999999999294, 
    16.9999999999305, 24.9999999999297, 21.99999999993, 18.9999999999303, 
    26.9999999999295, 15.9999999999306, 23.9999999999298, 20.9999999999301, 
    28.9999999999293, 17.9999999999304, 25.9999999999296, 22.9999999999299, 
    19.9999999999302, 27.9999999999294, 16.9999999999305, 24.9999999999297, 
    21.99999999993, 18.9999999999303, 26.9999999999295, 23.9999999999298, 
    20.9999999999301, 28.9999999999293, 17.9999999999304, 25.9999999999296, 
    22.9999999999299, 19.9999999999302, 27.9999999999294, 24.9999999999297, 
    21.99999999993, 18.9999999999303, 26.9999999999295, 23.9999999999298, 
    20.9999999999301, 28.9999999999293, 25.9999999999296, 22.9999999999299, 
    19.9999999999302, 27.9999999999294, 24.9999999999297, 21.99999999993, 
    26.9999999999295, 23.9999999999298, 20.9999999999301, 28.9999999999293, 
    25.9999999999296, 22.9999999999299, 27.9999999999294, 24.9999999999297, 
    21.99999999993, 29.9999999999292, 26.9999999999295, 23.9999999999298, 
    28.9999999999293, 25.9999999999296, 22.9999999999299, 27.9999999999294, 
    24.9999999999297, 29.9999999999292, 26.9999999999295, 23.9999999999298, 
    28.9999999999293, 25.9999999999296, 27.9999999999294, 24.9999999999297, 
    29.9999999999292, 26.9999999999295, 28.9999999999293, 25.9999999999296, 
    27.9999999999294, 26.9999999999295, 28.9999999999293, 27.9999999999294, 
    29.9999999999292, 28.9999999999293 ;

 obs_Ygrid = 2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36.0272723111239, 36.9000015258789, 38.0571408952985, 
    38.7000045776367, 39.9857155936105, 41.0999977111816, 41.8875017166138, 
    42.9000015258789, 44.0999984741211, 45.042856488909, 45.9000015258789, 
    47.0699981689453, 48, 48.9000018726696, 50.1272714788263, 51, 
    51.9000015258789, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0727258162065, 36, 
    36.9000015258789, 38.0999977111816, 38.9142870221819, 39.9000011444092, 
    41.1999969482422, 42.0999984741211, 42.8625011444092, 45.2999954223633, 
    45.9000026157924, 47.0999977111816, 48, 48.9000015258789, 
    50.0999994277954, 51, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.8000011444092, 38.1428555079869, 38.7750034332275, 40.1000022888183, 
    40.9499988555908, 42.0999984741211, 42.75, 43.7999954223633, 
    45.0599990844727, 46.0000038146972, 47.0999984741211, 48, 
    48.9000015258789, 50.1374988555908, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.1666653951009, 33, 34.020002746582, 35.0727258162065, 
    35.9333343505859, 36.9857155936105, 38.1857136317662, 38.7000045776367, 
    40.9499988555908, 41.9250011444092, 45.0999984741211, 45.9000027974446, 
    47.0999984741211, 48, 48.9000015258789, 50.0999984741211, 51, 
    51.9000015258789, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 32.2799995422363, 33, 
    33.9272741837935, 35.0142844063895, 35.9142870221819, 40.9499988555908, 
    42, 45.1124982833862, 45.9272741837935, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 50.9727276888761, 51.8625011444092, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 45.960001373291, 47.0999984741211, 
    48, 50.0999984741211, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0727258162065, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.1299983978271, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 
    20.9727276888761, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.8625011444092, 20.1374988555908, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 17.9625005722046, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    16.979997253418, 2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 
    11.8500022888184, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 11.8500022888184, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.86250114440917, 10.9499988555908, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.86250114440917, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.05714089529856, 8.94000091552734, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 2.10000038146972, 
    3, 3.89999961853028, 5.10000038146972, 23.7539978027344, 
    23.7539978027344, 23.7539978027344, 23.7539978027344, 23.7539978027344, 
    23.7539978027344, 23.7539978027344, 23.7539978027344, 23.7539978027344, 
    23.7539978027344, 23.7539978027344, 23.7539978027344, 23.7539978027344, 
    23.7539978027344, 23.7539978027344, 23.7539978027344, 23.7539978027344, 
    23.7539978027344, 23.7539978027344, 23.7539978027344, 23.7539978027344, 
    23.7539978027344, 23.7539978027344, 23.7539978027344, 23.7539978027344, 
    23.7539978027344, 23.7539978027344, 23.7539978027344, 23.7539978027344, 
    23.7539978027344, 23.7539978027344, 23.7539978027344, 23.7539978027344, 
    23.7539978027344, 23.7539978027344, 23.7539978027344, 23.7539978027344, 
    23.7539978027344, 26.3579978942871, 26.3579978942871, 26.3579978942871, 
    26.3579978942871, 26.3579978942871, 26.3579978942871, 26.3579978942871, 
    26.3579978942871, 26.3579978942871, 26.3579978942871, 26.3579978942871, 
    26.3579978942871, 26.3579978942871, 26.3579978942871, 26.3579978942871, 
    26.3579978942871, 26.3579978942871, 26.3579978942871, 26.3579978942871, 
    26.3579978942871, 26.3579978942871, 26.3579978942871, 26.3579978942871, 
    26.3579978942871, 26.3579978942871, 26.3579978942871, 26.3579978942871, 
    26.3579978942871, 26.3579978942871, 26.3579978942871, 26.3579978942871, 
    26.3579978942871, 26.3579978942871, 26.3579978942871, 26.3579978942871, 
    26.3579978942871, 26.3579978942871, 26.3579978942871, 26.3579978942871, 
    26.3579978942871, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36.0272723111239, 36.9000015258789, 38.0571408952985, 
    38.7000045776367, 39.9000005722046, 41.0999977111816, 41.8875017166138, 
    42.9000015258789, 44.0999984741211, 45.042856488909, 45.9000015258789, 
    47.0699981689453, 48, 48.9000018726696, 50.1599990844726, 51, 
    51.9000015258789, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0727258162065, 36, 
    36.9000015258789, 38.0999977111816, 38.9142870221819, 39.9000011444092, 
    41.1999969482422, 42.0999984741211, 42.8625011444092, 45.2999954223633, 
    45.9000026157924, 47.0999977111816, 48, 48.9000015258789, 
    50.2000007629394, 51, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000022888184, 35.0999984741211, 36, 
    36.8000011444092, 38.1428555079869, 38.7750034332275, 40.1000022888183, 
    40.9499988555908, 42.0999984741211, 42.75, 43.7999954223633, 
    45.0599990844727, 46.0000038146972, 47.0999984741211, 48, 
    48.9000015258789, 50.1374988555908, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.1666653951009, 33, 34.020002746582, 35.0727258162065, 
    35.9333343505859, 36.9857155936105, 38.1857136317662, 38.7000045776367, 
    40.9499988555908, 41.9250011444092, 45.0999984741211, 45.9000027974446, 
    47.0999984741211, 48, 48.9000015258789, 50.0999984741211, 51, 
    51.9000015258789, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 32.2799995422363, 
    33.0374994277954, 33.9272741837935, 35.0142844063895, 35.9142870221819, 
    40.9499988555908, 42, 45.1124982833862, 45.9272741837935, 
    47.0999984741211, 48, 48.9000015258789, 50.0999984741211, 
    50.9727276888761, 51.8625011444092, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 
    45.960001373291, 47.0999984741211, 48, 50.0999984741211, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0727258162065, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.1299983978271, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 
    20.9727276888761, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.8625011444092, 20.1374988555908, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 17.9625005722046, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    16.979997253418, 2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 
    11.8500022888184, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 11.8500022888184, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.86250114440917, 10.9499988555908, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.86250114440917, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.05714089529856, 8.94000091552734, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 2.10000038146972, 
    3, 3.89999961853028, 5.10000038146972, 13.3680038452148, 
    13.3680038452148, 13.3680038452148, 13.3680038452148, 13.3680038452148, 
    13.3680038452148, 13.3680038452148, 13.3680038452148, 13.3680038452148, 
    13.3680038452148, 13.3680038452148, 13.3680038452148, 13.3680038452148, 
    13.3680038452148, 13.3680038452148, 13.3680038452148, 13.3680038452148, 
    13.3680038452148, 13.3680038452148, 13.3680038452148, 13.3680038452148, 
    13.3680038452148, 13.3680038452148, 13.3680038452148, 13.3680038452148, 
    13.3680038452148, 13.3680038452148, 13.3680038452148, 13.3680038452148, 
    13.3680038452148, 13.3680038452148, 13.3680038452148, 13.3680038452148, 
    13.3680038452148, 13.3680038452148, 13.3680038452148, 13.3680038452148, 
    13.3680038452148, 13.3680038452148, 13.3680038452148, 13.3680038452148, 
    13.3680038452148, 13.3680038452148, 13.3680038452148, 13.3680038452148, 
    13.3680038452148, 37.7250022888184, 37.7250022888184, 37.7250022888184, 
    37.7250022888184, 37.7250022888184, 37.7250022888184, 37.7250022888184, 
    37.7250022888184, 37.7250022888184, 37.7250022888184, 37.7250022888184, 
    37.7250022888184, 37.7250022888184, 37.7250022888184, 37.7250022888184, 
    37.7250022888184, 37.7250022888184, 37.7250022888184, 37.7250022888184, 
    37.7250022888184, 37.7250022888184, 37.7250022888184, 37.7250022888184, 
    37.7250022888184, 37.7250022888184, 37.7250022888184, 37.7250022888184, 
    37.7250022888184, 37.7250022888184, 37.7250022888184, 37.7250022888184, 
    37.7250022888184, 37.7250022888184, 37.7250022888184, 37.7250022888184, 
    37.7250022888184, 37.7250022888184, 37.7250022888184, 37.7250022888184, 
    37.7250022888184, 37.7250022888184, 37.7250022888184, 37.7250022888184, 
    37.7250022888184, 37.7250022888184, 37.7250022888184, 45.6870002746582, 
    45.6870002746582, 45.6870002746582, 45.6870002746582, 45.6870002746582, 
    45.6870002746582, 45.6870002746582, 45.6870002746582, 45.6870002746582, 
    45.6870002746582, 45.6870002746582, 45.6870002746582, 45.6870002746582, 
    45.6870002746582, 45.6870002746582, 45.6870002746582, 2.10000038146972, 
    3, 3.89999961853028, 5.10000038146972, 5.99999809265136, 
    6.90000152587891, 8.09999847412109, 9, 9.90000152587891, 
    11.0999984741211, 12, 12.9000015258789, 14.0999984741211, 15, 
    15.9000015258789, 17.0999984741211, 18, 18.9000015258789, 
    20.0999984741211, 21, 21.9000015258789, 23.0999984741211, 24, 
    24.9000015258789, 26.0999984741211, 27, 27.9000015258789, 
    29.0999984741211, 30, 30.9000015258789, 32.0999984741211, 33, 
    33.9000015258789, 35.0999984741211, 36, 36.9000015258789, 
    38.0999984741211, 39, 39.9000015258789, 41.0999984741211, 42, 
    42.9000015258789, 44.0999984741211, 45, 45.9000015258789, 
    47.0999984741211, 48, 48.9000015258789, 50.0999984741211, 51, 
    51.9000015258789, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 
    36.0666656494141, 36.9000015258789, 37.874997138977, 39.9000005722046, 
    40.7999954223633, 41.8285740443638, 42.9000015258789, 44.0999984741211, 
    45.042856488909, 45.9000022888184, 47.0999981273304, 48, 
    48.9000018726696, 50.1599990844726, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0727258162065, 
    36.033332824707, 36.9000015258789, 38.0999977111816, 38.9500007629395, 
    39.9000011444092, 40.7999954223633, 41.8500022888184, 42.8625011444092, 
    45.2999954223633, 45.9000034332275, 47.0999977111816, 48, 
    48.9000015258789, 50.2000007629394, 51, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.8250017166138, 
    35.0999965667724, 36.0999984741211, 36.7000007629395, 38.1428555079869, 
    38.7750034332275, 40.1000022888183, 41.1000022888183, 42.0599990844727, 
    42.75, 43.7999954223633, 45.2999954223633, 46.0000038146972, 
    47.0999984741211, 48, 48.9000015258789, 50.0999984741211, 51, 
    51.9000015258789, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.8727285211736, 
    32.1666653951009, 32.9700004577637, 33.6000022888184, 35.0399963378906, 
    35.7000045776367, 38.1750011444092, 38.7000045776367, 40.9499988555908, 
    42.1499977111816, 45.1499977111816, 45.9000027974446, 47.0999984741211, 
    48, 48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 32.2799995422363, 
    33.0374994277954, 33.9000015258789, 36, 42.1499977111816, 
    45.1124982833862, 45.9272741837935, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 50.9727276888761, 51.8625011444092, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 45.960001373291, 47.0999984741211, 
    48, 50.0999984741211, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0727258162065, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.1299983978271, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 
    20.9727276888761, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.8625011444092, 20.1374988555908, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 17.9625005722046, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    16.979997253418, 2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 
    11.8500022888184, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 11.8500022888184, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.86250114440917, 10.9499988555908, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.86250114440917, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.05714089529856, 8.94000091552734, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 2.10000038146972, 
    3, 3.89999961853028, 5.10000038146972, 34.7880020141601, 
    34.7880020141601, 34.7880020141601, 34.7880020141601, 34.7880020141601, 
    34.7880020141601, 34.7880020141601, 34.7880020141601, 34.7880020141601, 
    34.7880020141601, 34.7880020141601, 34.7880020141601, 34.7880020141601, 
    33.6509971618652, 33.6509971618652, 33.6509971618652, 33.6509971618652, 
    33.6509971618652, 33.6509971618652, 33.6509971618652, 33.6509971618652, 
    33.6509971618652, 33.6509971618652, 33.6509971618652, 33.6509971618652, 
    33.6509971618652, 33.6509971618652, 8.8440055847168, 8.8440055847168, 
    8.8440055847168, 8.8440055847168, 8.8440055847168, 8.8440055847168, 
    8.8440055847168, 8.8440055847168, 8.8440055847168, 8.8440055847168, 
    8.8440055847168, 8.8440055847168, 8.8440055847168, 8.8440055847168, 
    8.7509994506836, 8.7509994506836, 8.7509994506836, 8.7509994506836, 
    8.7509994506836, 8.7509994506836, 8.7509994506836, 8.7509994506836, 
    8.7509994506836, 8.7509994506836, 8.7509994506836, 8.7509994506836, 
    8.7509994506836, 8.7509994506836, 8.7509994506836, 8.7509994506836, 
    8.7509994506836, 8.7509994506836, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999981273304, 30, 
    30.8727285211736, 32.0999984741211, 33, 33.9000015258789, 
    35.0727258162065, 36.042856488909, 36.8625011444092, 38.1000022888183, 
    42.9000015258789, 44.0999988555908, 45.0374994277954, 45.8666687011719, 
    47.0999981273304, 48, 48.9000015258789, 50.0999984741211, 51, 
    51.9000015258789, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999981273304, 30, 30.9000015258789, 
    32.0999981273304, 32.8800018310547, 34.0285737173898, 34.9874982833862, 
    36.0999984741211, 36.8000005086263, 37.9499988555908, 44.1750011444092, 
    45.1499977111816, 45.7500028610229, 47.1299983978271, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.8625011444092, 29.0624985694885, 30, 30.8571444920131, 
    31.979997253418, 34.7999954223633, 36.2999954223633, 45.1499977111816, 
    46.0000019073486, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.8625011444092, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0727258162065, 
    29.9727276888761, 32.2124991416931, 32.9700004577637, 33.6000022888184, 
    38.7000045776367, 45.1499977111816, 45.9000022888184, 47.0999984741211, 
    48, 48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 29.9142870221819, 32.2799995422363, 
    33, 33.6000022888184, 45.1124982833862, 45.9272741837935, 
    47.0999984741211, 48, 48.9000015258789, 50.0999984741211, 
    50.9727276888761, 51.8625011444092, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 
    45.960001373291, 47.0999984741211, 48, 50.0999984741211, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0727258162065, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 
    20.9727276888761, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.8625011444092, 20.1374988555908, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 17.9625005722046, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    16.979997253418, 2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 
    11.8500022888184, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 11.8500022888184, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.86250114440917, 10.9499988555908, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.86250114440917, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.05714089529856, 8.94000091552734, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 2.10000038146972, 
    3, 3.89999961853028, 5.10000038146972, 8.04899597167969, 
    8.04899597167969, 8.04899597167969, 8.04899597167969, 8.04899597167969, 
    8.04899597167969, 8.04899597167969, 8.04899597167969, 8.04899597167969, 
    8.04899597167969, 8.04899597167969, 8.04899597167969, 8.04899597167969, 
    8.04899597167969, 8.04899597167969, 8.04899597167969, 8.04899597167969, 
    8.04899597167969, 7.04100036621093, 7.04100036621093, 7.04100036621093, 
    7.04100036621093, 7.04100036621093, 7.04100036621093, 7.04100036621093, 
    7.04100036621093, 7.04100036621093, 7.04100036621093, 7.04100036621093, 
    7.04100036621093, 7.04100036621093, 7.04100036621093, 7.04100036621093, 
    7.04100036621093, 7.04100036621093, 7.04100036621093, 7.04100036621093, 
    7.04100036621093, 7.04100036621093, 7.04100036621093, 7.04100036621093, 
    7.04100036621093, 7.04100036621093, 7.04100036621093, 7.04100036621093, 
    7.04100036621093, 7.04100036621093, 7.04100036621093, 2.8511893712683, 
    2.8511893712683, 3.70751696511747, 2.8511893712683, 3.70751696511747, 
    2.8511893712683, 3.70751696511747, 2.8511893712683, 3.70751696511747, 
    6.26097000315193, 2.8511893712683, 3.70751696511747, 6.26097000315193, 
    2.8511893712683, 7.10690132310917, 3.70751696511747, 6.26097000315193, 
    2.8511893712683, 7.10690132310917, 3.70751696511747, 6.26097000315193, 
    7.95020197539848, 2.8511893712683, 7.10690132310917, 3.70751696511747, 
    6.26097000315193, 7.95020197539848, 2.8511893712683, 7.10690132310917, 
    8.79085990591997, 3.70751696511747, 6.26097000315193, 7.95020197539848, 
    2.8511893712683, 7.10690132310917, 8.79085990591997, 3.70751696511747, 
    6.26097000315193, 7.95020197539848, 2.8511893712683, 9.62886335158985, 
    7.10690132310916, 8.79085990591997, 3.70751696511747, 6.26097000315193, 
    7.95020197539848, 2.8511893712683, 9.62886335158985, 7.10690132310917, 
    8.79085990591997, 3.70751696511747, 11.296861184434, 6.26097000315193, 
    7.95020197539848, 2.8511893712683, 9.62886335158985, 7.10690132310917, 
    8.79085990591997, 3.70751696511747, 11.296861184434, 6.26097000315193, 
    7.95020197539848, 2.8511893712683, 9.62886335158985, 12.126833490299, 
    7.10690132310916, 8.79085990591997, 3.70751696511747, 11.296861184434, 
    6.26097000315193, 7.95020197539848, 2.8511893712683, 9.62886335158985, 
    12.126833490299, 7.10690132310917, 8.79085990591997, 3.70751696511747, 
    11.296861184434, 6.26097000315193, 12.9541071462105, 7.95020197539848, 
    2.8511893712683, 9.62886335158985, 12.126833490299, 7.10690132310916, 
    8.79085990591997, 3.70751696511747, 11.296861184434, 6.26097000315193, 
    12.9541071462105, 7.95020197539848, 2.8511893712683, 9.62886335158985, 
    12.126833490299, 7.10690132310916, 13.7786718264961, 8.79085990591997, 
    3.70751696511747, 11.296861184434, 6.26097000315193, 12.9541071462105, 
    7.95020197539848, 2.8511893712683, 9.62886335158985, 12.126833490299, 
    7.10690132310917, 13.7786718264961, 8.79085990591997, 3.70751696511747, 
    11.296861184434, 6.26097000315193, 12.9541071462105, 7.95020197539848, 
    2.8511893712683, 14.60051748906, 9.62886335158985, 12.126833490299, 
    7.10690132310916, 13.7786718264961, 8.79085990591997, 3.70751696511747, 
    11.296861184434, 6.26097000315193, 12.9541071462105, 7.95020197539848, 
    2.8511893712683, 14.60051748906, 9.62886335158985, 12.126833490299, 
    7.10690132310916, 13.7786718264961, 8.79085990591997, 3.70751696511747, 
    16.2360130019538, 11.296861184434, 6.26097000315193, 12.9541071462105, 
    7.95020197539848, 2.8511893712683, 14.60051748906, 9.62886335158985, 
    12.126833490299, 7.10690132310917, 13.7786718264961, 8.79085990591997, 
    3.70751696511747, 16.2360130019538, 11.296861184434, 6.26097000315193, 
    12.9541071462105, 7.95020197539848, 2.8511893712683, 14.60051748906, 
    9.62886335158985, 17.0496441729557, 12.126833490299, 7.10690132310917, 
    13.7786718264961, 8.79085990591997, 3.70751696511747, 16.2360130019538, 
    11.296861184434, 6.26097000315193, 12.9541071462105, 7.95020197539848, 
    2.8511893712683, 14.60051748906, 9.62886335158985, 17.0496441729557, 
    12.126833490299, 7.10690132310917, 13.7786718264961, 8.79085990591997, 
    3.70751696511747, 16.2360130019538, 11.296861184434, 6.26097000315193, 
    17.860518964504, 12.9541071462105, 7.95020197539848, 2.8511893712683, 
    14.60051748906, 9.62886335158985, 17.0496441729557, 12.126833490299, 
    7.10690132310916, 13.7786718264961, 8.79085990591997, 3.70751696511747, 
    16.2360130019538, 11.296861184434, 6.26097000315193, 17.860518964504, 
    12.9541071462105, 7.95020197539848, 2.8511893712683, 14.60051748906, 
    9.62886335158985, 17.0496441729557, 12.126833490299, 7.10690132310916, 
    18.6686287301423, 13.7786718264961, 8.79085990591997, 3.70751696511747, 
    16.2360130019538, 11.296861184434, 6.26097000315193, 17.860518964504, 
    12.9541071462105, 7.95020197539848, 2.8511893712683, 14.60051748906, 
    9.62886335158985, 17.0496441729557, 12.126833490299, 7.10690132310917, 
    18.6686287301423, 13.7786718264961, 8.79085990591997, 3.70751696511747, 
    16.2360130019538, 11.296861184434, 6.26097000315193, 17.860518964504, 
    12.9541071462105, 7.95020197539848, 20.2765199679718, 2.8511893712683, 
    14.60051748906, 9.62886335158985, 17.0496441729557, 12.126833490299, 
    7.10690132310916, 18.6686287301423, 13.7786718264961, 8.79085990591997, 
    3.70751696511747, 16.2360130019538, 11.296861184434, 6.26097000315193, 
    17.860518964504, 12.9541071462105, 7.95020197539848, 20.2765199679718, 
    2.8511893712683, 14.60051748906, 9.62886335158985, 17.0496441729557, 
    12.126833490299, 7.10690132310917, 18.6686287301423, 13.7786718264961, 
    8.79085990591997, 21.0762855122492, 3.70751696511747, 16.2360130019538, 
    11.296861184434, 6.26097000315193, 17.860518964504, 12.9541071462105, 
    7.95020197539848, 20.2765199679718, 2.8511893712683, 14.60051748906, 
    9.62886335158985, 17.0496441729557, 12.126833490299, 7.10690132310917, 
    18.6686287301423, 13.7786718264961, 8.79085990591997, 21.0762855122492, 
    3.70751696511747, 16.2360130019538, 11.296861184434, 6.26097000315193, 
    17.860518964504, 12.9541071462105, 7.95020197539848, 20.2765199679718, 
    2.8511893712683, 14.60051748906, 9.62886335158985, 21.8732541712884, 
    17.0496441729557, 12.126833490299, 7.10690132310916, 18.6686287301423, 
    13.7786718264961, 8.79085990591997, 21.0762855122492, 3.70751696511747, 
    16.2360130019538, 11.296861184434, 6.26097000315193, 17.860518964504, 
    12.9541071462105, 7.95020197539848, 20.2765199679718, 2.8511893712683, 
    14.60051748906, 9.62886335158985, 21.8732541712884, 17.0496441729557, 
    12.126833490299, 7.10690132310917, 18.6686287301423, 13.7786718264961, 
    8.79085990591997, 21.0762855122492, 3.70751696511747, 16.2360130019538, 
    11.296861184434, 22.6674186531335, 6.26097000315193, 17.860518964504, 
    12.9541071462105, 7.95020197539848, 20.2765199679718, 2.8511893712683, 
    14.60051748906, 9.62886335158985, 21.8732541712884, 17.0496441729557, 
    12.126833490299, 7.10690132310917, 18.6686287301423, 13.7786718264961, 
    8.79085990591997, 21.0762855122492, 3.70751696511747, 16.2360130019538, 
    11.296861184434, 22.6674186531335, 6.26097000315193, 17.860518964504, 
    12.9541071462105, 7.95020197539848, 20.2765199679718, 2.8511893712683, 
    14.60051748906, 9.62886335158985, 21.8732541712884, 17.0496441729557, 
    12.126833490299, 24.2473072431218, 7.10690132310916, 18.6686287301423, 
    13.7786718264961, 8.79085990591997, 21.0762855122492, 3.70751696511747, 
    16.2360130019538, 11.296861184434, 22.6674186531335, 6.26097000315193, 
    17.860518964504, 12.9541071462105, 7.95020197539848, 20.2765199679718, 
    2.8511893712683, 14.60051748906, 9.62886335158985, 21.8732541712884, 
    17.0496441729557, 12.126833490299, 24.2473072431218, 7.10690132310916, 
    18.6686287301423, 13.7786718264961, 8.79085990591997, 21.0762855122492, 
    3.70751696511747, 16.2360130019538, 11.296861184434, 22.6674186531335, 
    6.26097000315193, 17.860518964504, 12.9541071462105, 25.0330180873813, 
    7.95020197539848, 20.2765199679718, 2.8511893712683, 14.60051748906, 
    9.62886335158985, 21.8732541712884, 17.0496441729557, 12.126833490299, 
    24.2473072431218, 7.10690132310917, 18.6686287301423, 13.7786718264961, 
    8.79085990591997, 21.0762855122492, 3.70751696511747, 16.2360130019538, 
    11.296861184434, 22.6674186531335, 6.26097000315193, 17.860518964504, 
    12.9541071462105, 25.0330180873813, 7.95020197539848, 20.2765199679718, 
    2.8511893712683, 14.60051748906, 9.62886335158985, 21.8732541712884, 
    17.0496441729557, 12.126833490299, 24.2473072431218, 7.10690132310916, 
    18.6686287301423, 13.7786718264961, 25.8158982228162, 8.79085990591997, 
    21.0762855122492, 3.70751696511747, 16.2360130019538, 11.296861184434, 
    22.6674186531335, 6.26097000315193, 17.860518964504, 12.9541071462105, 
    25.0330180873813, 7.95020197539848, 20.2765199679718, 2.8511893712683, 
    14.60051748906, 9.62886335158985, 21.8732541712884, 17.0496441729557, 
    12.126833490299, 24.2473072431218, 7.10690132310916, 18.6686287301423, 
    13.7786718264961, 25.8158982228162, 8.79085990591997, 21.0762855122492, 
    3.70751696511747, 16.2360130019538, 11.296861184434, 22.6674186531335, 
    6.26097000315193, 17.860518964504, 12.9541071462105, 25.0330180873813, 
    7.95020197539848, 20.2765199679718, 2.8511893712683, 14.60051748906, 
    26.9845421774241, 9.62886335158985, 21.8732541712884, 17.0496441729557, 
    12.126833490299, 24.2473072431218, 7.10690132310916, 18.6686287301423, 
    13.7786718264961, 25.8158982228162, 8.79085990591997, 21.0762855122492, 
    3.70751696511747, 16.2360130019538, 11.296861184434, 22.6674186531335, 
    6.26097000315193, 17.860518964504, 12.9541071462105, 25.0330180873813, 
    7.95020197539848, 20.2765199679718, 2.8511893712683, 14.60051748906, 
    26.9845421774241, 9.62886335158985, 21.8732541712884, 17.0496441729557, 
    12.126833490299, 24.2473072431218, 7.10690132310916, 18.6686287301423, 
    13.7786718264961, 25.8158982228162, 8.79085990591997, 21.0762855122492, 
    3.70751696511747, 16.2360130019538, 28.147495817899, 11.296861184434, 
    22.6674186531335, 6.26097000315193, 17.860518964504, 12.9541071462105, 
    25.0330180873813, 7.95020197539848, 20.2765199679718, 2.8511893712683, 
    14.60051748906, 26.9845421774241, 9.62886335158985, 21.8732541712884, 
    17.0496441729557, 12.126833490299, 24.2473072431218, 7.10690132310916, 
    18.6686287301423, 13.7786718264961, 25.8158982228162, 8.79085990591997, 
    21.0762855122492, 3.70751696511747, 16.2360130019538, 28.147495817899, 
    11.296861184434, 22.6674186531335, 6.26097000315193, 17.860518964504, 
    12.9541071462105, 25.0330180873813, 7.95020197539848, 20.2765199679718, 
    2.8511893712683, 14.60051748906, 26.9845421774241, 9.62886335158985, 
    21.8732541712884, 17.0496441729557, 28.9189958304827, 12.126833490299, 
    24.2473072431218, 7.10690132310916, 18.6686287301423, 13.7786718264961, 
    25.8158982228162, 8.79085990591997, 21.0762855122492, 3.70751696511747, 
    16.2360130019538, 28.147495817899, 11.296861184434, 22.6674186531335, 
    6.26097000315193, 17.860518964504, 12.9541071462105, 25.0330180873813, 
    7.95020197539848, 20.2765199679718, 2.8511893712683, 14.60051748906, 
    26.9845421774241, 9.62886335158985, 21.8732541712884, 17.0496441729557, 
    28.9189958304827, 12.126833490299, 24.2473072431218, 7.10690132310917, 
    18.6686287301423, 13.7786718264961, 25.8158982228162, 8.79085990591997, 
    21.0762855122492, 3.70751696511747, 16.2360130019538, 28.147495817899, 
    11.296861184434, 22.6674186531335, 6.26097000315193, 17.860518964504, 
    29.6876377539464, 12.9541071462105, 25.0330180873813, 7.95020197539848, 
    20.2765199679718, 2.8511893712683, 14.60051748906, 26.9845421774241, 
    9.62886335158985, 21.8732541712884, 17.0496441729557, 28.9189958304827, 
    12.126833490299, 24.2473072431218, 7.10690132310916, 18.6686287301423, 
    13.7786718264961, 25.8158982228162, 8.79085990591997, 21.0762855122492, 
    3.70751696511747, 16.2360130019538, 28.147495817899, 11.296861184434, 
    22.6674186531335, 6.26097000315193, 17.860518964504, 29.6876377539464, 
    12.9541071462105, 25.0330180873813, 7.95020197539848, 20.2765199679718, 
    2.8511893712683, 14.60051748906, 26.9845421774241, 9.62886335158985, 
    21.8732541712884, 17.0496441729557, 28.9189958304827, 12.126833490299, 
    24.2473072431218, 7.10690132310916, 18.6686287301423, 31.2163286776756, 
    13.7786718264961, 25.8158982228162, 8.79085990591997, 21.0762855122492, 
    3.70751696511747, 16.2360130019538, 28.147495817899, 11.296861184434, 
    22.6674186531335, 6.26097000315193, 17.860518964504, 29.6876377539464, 
    12.9541071462105, 25.0330180873813, 7.95020197539848, 20.2765199679718, 
    2.8511893712683, 14.60051748906, 26.9845421774241, 9.62886335158985, 
    21.8732541712884, 17.0496441729557, 28.9189958304827, 12.126833490299, 
    24.2473072431218, 7.10690132310917, 18.6686287301423, 31.2163286776756, 
    13.7786718264961, 25.8158982228162, 8.79085990591997, 21.0762855122492, 
    3.70751696511747, 16.2360130019538, 28.147495817899, 11.296861184434, 
    22.6674186531335, 6.26097000315193, 17.860518964504, 29.6876377539464, 
    12.9541071462105, 25.0330180873813, 7.95020197539848, 20.2765199679718, 
    31.9763689611184, 2.8511893712683, 14.60051748906, 26.9845421774241, 
    9.62886335158985, 21.8732541712884, 17.0496441729557, 28.9189958304827, 
    12.126833490299, 24.2473072431218, 7.10690132310916, 18.6686287301423, 
    31.2163286776756, 13.7786718264961, 25.8158982228162, 8.79085990591997, 
    21.0762855122492, 3.70751696511747, 16.2360130019538, 28.147495817899, 
    11.296861184434, 22.6674186531335, 6.26097000315193, 17.860518964504, 
    29.6876377539464, 12.9541071462105, 25.0330180873813, 7.95020197539848, 
    20.2765199679718, 31.9763689611184, 2.8511893712683, 14.60051748906, 
    26.9845421774241, 9.62886335158985, 21.8732541712884, 17.0496441729557, 
    28.9189958304827, 12.126833490299, 24.2473072431218, 7.10690132310916, 
    18.6686287301423, 31.2163286776756, 13.7786718264961, 25.8158982228162, 
    8.79085990591997, 21.0762855122492, 32.7335337174312, 3.70751696511747, 
    16.2360130019538, 28.147495817899, 11.296861184434, 22.6674186531335, 
    6.26097000315193, 17.860518964504, 29.6876377539464, 12.9541071462105, 
    25.0330180873813, 7.95020197539848, 20.2765199679718, 31.9763689611184, 
    2.8511893712683, 14.60051748906, 26.9845421774241, 9.62886335158985, 
    21.8732541712884, 17.0496441729557, 28.9189958304827, 12.126833490299, 
    24.2473072431218, 7.10690132310916, 18.6686287301423, 31.2163286776756, 
    13.7786718264961, 25.8158982228162, 8.79085990591997, 21.0762855122492, 
    32.7335337174312, 3.70751696511747, 16.2360130019538, 28.147495817899, 
    11.296861184434, 22.6674186531335, 6.26097000315193, 17.860518964504, 
    29.6876377539464, 12.9541071462105, 25.0330180873813, 7.95020197539848, 
    20.2765199679718, 31.9763689611184, 2.8511893712683, 14.60051748906, 
    26.9845421774241, 9.62886335158985, 21.8732541712884, 34.2392218564619, 
    17.0496441729557, 28.9189958304827, 12.126833490299, 24.2473072431218, 
    7.10690132310916, 18.6686287301423, 31.2163286776756, 13.7786718264961, 
    25.8158982228162, 8.79085990591997, 21.0762855122492, 32.7335337174312, 
    3.70751696511747, 16.2360130019538, 28.147495817899, 11.296861184434, 
    22.6674186531335, 6.26097000315193, 17.860518964504, 29.6876377539464, 
    12.9541071462105, 25.0330180873813, 7.95020197539848, 20.2765199679718, 
    31.9763689611184, 14.60051748906, 26.9845421774241, 9.62886335158985, 
    21.8732541712884, 34.2392218564619, 17.0496441729557, 28.9189958304827, 
    12.126833490299, 24.2473072431218, 7.10690132310917, 18.6686287301423, 
    31.2163286776756, 13.7786718264961, 25.8158982228162, 8.79085990591997, 
    21.0762855122492, 32.7335337174312, 3.70751696511747, 16.2360130019538, 
    28.147495817899, 11.296861184434, 22.6674186531335, 34.9877384320501, 
    6.26097000315193, 17.860518964504, 29.6876377539464, 12.9541071462105, 
    25.0330180873813, 7.95020197539848, 20.2765199679718, 31.9763689611184, 
    14.60051748906, 26.9845421774241, 9.62886335158985, 21.8732541712884, 
    34.2392218564619, 17.0496441729557, 28.9189958304827, 12.126833490299, 
    24.2473072431218, 7.10690132310917, 18.6686287301423, 31.2163286776756, 
    13.7786718264961, 25.8158982228162, 8.79085990591997, 21.0762855122492, 
    32.7335337174312, 16.2360130019538, 28.147495817899, 11.296861184434, 
    22.6674186531335, 34.9877384320501, 6.26097000315193, 17.860518964504, 
    29.6876377539464, 12.9541071462105, 25.0330180873813, 7.95020197539848, 
    20.2765199679718, 31.9763689611184, 14.60051748906, 26.9845421774241, 
    9.62886335158985, 21.8732541712884, 34.2392218564619, 17.0496441729557, 
    28.9189958304827, 12.126833490299, 24.2473072431218, 35.7333658617202, 
    7.10690132310916, 18.6686287301423, 31.2163286776756, 13.7786718264961, 
    25.8158982228162, 8.79085990591997, 21.0762855122492, 32.7335337174312, 
    16.2360130019538, 28.147495817899, 11.296861184434, 22.6674186531335, 
    34.9877384320501, 6.26097000315193, 17.860518964504, 29.6876377539464, 
    12.9541071462105, 25.0330180873813, 7.95020197539848, 20.2765199679718, 
    31.9763689611184, 14.60051748906, 26.9845421774241, 9.62886335158985, 
    21.8732541712884, 34.2392218564619, 17.0496441729557, 28.9189958304827, 
    12.126833490299, 24.2473072431218, 35.7333658617202, 7.10690132310917, 
    18.6686287301423, 31.2163286776756, 13.7786718264961, 25.8158982228162, 
    8.79085990591997, 21.0762855122492, 32.7335337174312, 16.2360130019538, 
    28.147495817899, 11.296861184434, 22.6674186531335, 34.9877384320501, 
    17.860518964504, 29.6876377539464, 12.9541071462105, 25.0330180873813, 
    37.2159422114215, 7.95020197539848, 20.2765199679718, 31.9763689611184, 
    14.60051748906, 26.9845421774241, 9.62886335158985, 21.8732541712884, 
    34.2392218564619, 17.0496441729557, 28.9189958304827, 12.126833490299, 
    24.2473072431218, 35.7333658617202, 18.6686287301423, 31.2163286776756, 
    13.7786718264961, 25.8158982228162, 21.0762855122492, 32.7335337174312, 
    16.2360130019538, 28.147495817899, 11.296861184434, 22.6674186531335, 
    34.9877384320501, 17.860518964504, 29.6876377539464, 12.9541071462105, 
    25.0330180873813, 37.2159422114215, 7.95020197539848, 20.2765199679718, 
    31.9763689611184, 14.60051748906, 26.9845421774241, 9.62886335158985, 
    21.8732541712884, 34.2392218564619, 17.0496441729557, 28.9189958304827, 
    24.2473072431218, 35.7333658617202, 18.6686287301423, 31.2163286776756, 
    25.8158982228162, 37.9528861616004, 21.0762855122492, 32.7335337174312, 
    16.2360130019538, 28.147495817899, 11.296861184434, 22.6674186531335, 
    34.9877384320501, 17.860518964504, 29.6876377539464, 12.9541071462105, 
    25.0330180873813, 37.2159422114215, 20.2765199679718, 31.9763689611184, 
    14.60051748906, 26.9845421774241, 21.8732541712884, 34.2392218564619, 
    17.0496441729557, 28.9189958304827, 24.2473072431218, 35.7333658617202, 
    18.6686287301423, 31.2163286776756, 25.8158982228162, 37.9528861616004, 
    21.0762855122492, 32.7335337174312, 16.2360130019538, 28.147495817899, 
    11.296861184434, 22.6674186531335, 34.9877384320501, 17.860518964504, 
    29.6876377539464, 25.0330180873813, 37.2159422114215, 20.2765199679718, 
    31.9763689611184, 26.9845421774241, 38.6869310214985, 21.8732541712884, 
    34.2392218564619, 17.0496441729557, 28.9189958304827, 24.2473072431218, 
    35.7333658617202, 18.6686287301423, 31.2163286776756, 25.8158982228162, 
    37.9528861616004, 21.0762855122492, 32.7335337174312, 28.147495817899, 
    22.6674186531335, 34.9877384320501, 17.860518964504, 29.6876377539464, 
    25.0330180873813, 37.2159422114215, 20.2765199679718, 31.9763689611184, 
    26.9845421774241, 38.6869310214985, 21.8732541712884, 34.2392218564619, 
    28.9189958304827, 24.2473072431218, 35.7333658617202, 18.6686287301423, 
    31.2163286776756, 25.8158982228162, 37.9528861616004, 21.0762855122492, 
    32.7335337174312, 28.147495817899, 40.146315971085, 22.6674186531335, 
    34.9877384320501, 29.6876377539464, 25.0330180873813, 37.2159422114215, 
    20.2765199679718, 31.9763689611184, 26.9845421774241, 38.6869310214985, 
    21.8732541712884, 34.2392218564619, 28.9189958304827, 24.2473072431218, 
    35.7333658617202, 31.2163286776756, 25.8158982228162, 37.9528861616004, 
    21.0762855122492, 32.7335337174312, 28.147495817899, 40.146315971085, 
    22.6674186531335, 34.9877384320501, 29.6876377539464, 25.0330180873813, 
    37.2159422114215, 20.2765199679718, 31.9763689611184, 26.9845421774241, 
    38.6869310214985, 21.8732541712884, 34.2392218564619, 28.9189958304827, 
    40.8716528537064, 24.2473072431218, 35.7333658617202, 31.2163286776756, 
    25.8158982228162, 37.9528861616004, 21.0762855122492, 32.7335337174312, 
    28.147495817899, 40.146315971085, 22.6674186531335, 34.9877384320501, 
    29.6876377539464, 25.0330180873813, 37.2159422114215, 31.9763689611184, 
    26.9845421774241, 38.6869310214985, 21.8732541712884, 34.2392218564619, 
    28.9189958304827, 40.8716528537064, 24.2473072431218, 35.7333658617202, 
    31.2163286776756, 25.8158982228162, 37.9528861616004, 32.7335337174312, 
    28.147495817899, 40.146315971085, 22.6674186531335, 34.9877384320501, 
    29.6876377539464, 42.313609019804, 25.0330180873813, 37.2159422114215, 
    31.9763689611184, 26.9845421774241, 38.6869310214985, 34.2392218564619, 
    28.9189958304827, 40.8716528537064, 24.2473072431218, 35.7333658617202, 
    31.2163286776756, 25.8158982228162, 37.9528861616004, 32.7335337174312, 
    28.147495817899, 40.146315971085, 22.6674186531335, 34.9877384320501, 
    29.6876377539464, 42.313609019804, 25.0330180873813, 37.2159422114215, 
    31.9763689611184, 26.9845421774241, 38.6869310214985, 34.2392218564619, 
    28.9189958304827, 40.8716528537064, 35.7333658617202, 31.2163286776756, 
    43.0302263684599, 25.8158982228162, 37.9528861616004, 32.7335337174312, 
    28.147495817899, 40.146315971085, 34.9877384320501, 29.6876377539464, 
    42.313609019804, 37.2159422114215, 31.9763689611184, 26.9845421774241, 
    38.6869310214985, 34.2392218564619, 28.9189958304827, 40.8716528537064, 
    35.7333658617202, 31.2163286776756, 43.0302263684599, 25.8158982228162, 
    37.9528861616004, 32.7335337174312, 28.147495817899, 40.146315971085, 
    34.9877384320501, 29.6876377539464, 42.313609019804, 37.2159422114215, 
    31.9763689611184, 43.743935615978, 26.9845421774241, 38.6869310214985, 
    34.2392218564619, 28.9189958304827, 40.8716528537064, 35.7333658617202, 
    31.2163286776756, 43.0302263684599, 37.9528861616004, 32.7335337174312, 
    28.147495817899, 40.146315971085, 34.9877384320501, 29.6876377539464, 
    42.313609019804, 37.2159422114215, 31.9763689611184, 43.7439356159779, 
    38.6869310214985, 34.2392218564619, 28.9189958304827, 40.8716528537064, 
    35.7333658617202, 31.2163286776756, 43.0302263684599, 37.9528861616004, 
    32.7335337174312, 45.1626281947156, 28.147495817899, 40.146315971085, 
    34.9877384320501, 29.6876377539464, 42.313609019804, 37.2159422114215, 
    31.9763689611184, 43.7439356159779, 38.6869310214985, 34.2392218564619, 
    28.9189958304827, 40.8716528537064, 35.7333658617202, 31.2163286776756, 
    43.0302263684599, 37.9528861616004, 32.7335337174312, 45.1626281947156, 
    40.146315971085, 34.9877384320501, 29.6876377539464, 42.313609019804, 
    37.2159422114215, 31.9763689611184, 43.7439356159779, 38.6869310214985, 
    34.2392218564619, 45.8676112200792, 28.9189958304827, 40.8716528537064, 
    35.7333658617202, 31.2163286776756, 43.0302263684599, 37.9528861616004, 
    32.7335337174312, 45.1626281947156, 40.146315971085, 34.9877384320501, 
    29.6876377539464, 42.313609019804, 37.2159422114215, 31.9763689611184, 
    43.7439356159779, 38.6869310214985, 34.2392218564619, 45.8676112200792, 
    40.8716528537064, 35.7333658617202, 31.2163286776756, 43.0302263684599, 
    37.9528861616004, 32.7335337174312, 45.1626281947156, 40.146315971085, 
    34.9877384320501, 47.268851454425, 42.313609019804, 37.2159422114215, 
    31.9763689611184, 43.7439356159779, 38.6869310214985, 34.2392218564619, 
    45.8676112200792, 40.8716528537064, 35.7333658617202, 43.0302263684599, 
    37.9528861616004, 32.7335337174312, 45.1626281947156, 40.146315971085, 
    34.9877384320501, 47.268851454425, 42.313609019804, 37.2159422114215, 
    31.9763689611184, 43.7439356159779, 38.6869310214985, 34.2392218564619, 
    45.8676112200792, 40.8716528537064, 35.7333658617202, 47.965109528352, 
    43.0302263684599, 37.9528861616004, 32.7335337174312, 45.1626281947156, 
    40.146315971085, 34.9877384320501, 47.268851454425, 42.313609019804, 
    37.2159422114215, 31.9763689611184, 43.7439356159779, 38.6869310214985, 
    34.2392218564619, 45.8676112200792, 40.8716528537064, 35.7333658617202, 
    47.965109528352, 43.0302263684599, 37.9528861616004, 32.7335337174312, 
    45.1626281947156, 40.146315971085, 34.9877384320501, 47.268851454425, 
    42.313609019804, 37.2159422114215, 49.0036828201845, 43.7439356159779, 
    38.6869310214985, 34.2392218564619, 45.8676112200792, 40.8716528537064, 
    35.7333658617202, 47.965109528352, 43.0302263684599, 37.9528861616004, 
    32.7335337174312, 45.1626281947156, 40.146315971085, 34.9877384320501, 
    47.268851454425, 42.313609019804, 37.2159422114215, 49.0036828201845, 
    43.7439356159779, 38.6869310214985, 45.8676112200792, 40.8716528537064, 
    35.7333658617202, 47.965109528352, 43.0302263684599, 37.9528861616004, 
    50.0364447368152, 45.1626281947156, 40.146315971085, 34.9877384320501, 
    47.268851454425, 42.313609019804, 37.2159422114215, 49.0036828201845, 
    43.7439356159779, 38.6869310214985, 45.8676112200792, 40.8716528537064, 
    35.7333658617202, 47.965109528352, 43.0302263684599, 37.9528861616004, 
    50.0364447368153, 45.1626281947156, 40.146315971085, 47.268851454425, 
    42.313609019804, 37.2159422114215, 49.0036828201845, 43.7439356159779, 
    38.6869310214985, 51.0619470586162, 45.8676112200792, 40.8716528537064, 
    35.7333658617202, 47.965109528352, 43.0302263684599, 37.9528861616004, 
    50.0364447368152, 45.1626281947156, 40.146315971085, 47.268851454425, 
    42.313609019804, 37.2159422114215, 49.0036828201845, 43.7439356159779, 
    38.6869310214985, 51.0619470586162, 45.8676112200792, 40.8716528537064, 
    47.965109528352, 43.0302263684599, 37.9528861616004, 50.0364447368153, 
    45.1626281947156, 40.146315971085, 47.268851454425, 42.313609019804, 
    37.2159422114215, 49.0036828201845, 43.7439356159779, 38.6869310214985, 
    51.0619470586162, 45.8676112200792, 40.8716528537064, 47.965109528352, 
    43.0302263684599, 37.9528861616004, 50.0364447368152, 45.1626281947156, 
    40.146315971085, 47.268851454425, 42.313609019804, 37.2159422114215, 
    49.0036828201845, 43.743935615978, 38.6869310214985, 51.0619470586162, 
    45.8676112200792, 40.8716528537064, 47.965109528352, 43.0302263684599, 
    37.9528861616004, 50.0364447368152, 45.1626281947156, 40.146315971085, 
    47.268851454425, 42.313609019804, 49.0036828201845, 43.7439356159779, 
    38.6869310214985, 51.0619470586162, 45.8676112200792, 40.8716528537064, 
    47.965109528352, 43.0302263684599, 37.9528861616004, 50.0364447368152, 
    45.1626281947156, 40.1463159710849, 47.268851454425, 42.313609019804, 
    49.0036828201845, 43.7439356159779, 38.6869310214985, 51.0619470586162, 
    45.8676112200792, 40.8716528537064, 47.965109528352, 43.0302263684599, 
    50.0364447368152, 45.1626281947156, 40.146315971085, 47.268851454425, 
    42.313609019804, 49.0036828201845, 43.743935615978, 38.6869310214985, 
    51.0619470586162, 45.8676112200792, 40.8716528537064, 47.965109528352, 
    43.0302263684599, 50.0364447368152, 45.1626281947156, 40.1463159710849, 
    47.268851454425, 42.313609019804, 49.0036828201845, 43.743935615978, 
    51.0619470586162, 45.8676112200792, 40.8716528537064, 47.965109528352, 
    43.0302263684599, 50.0364447368153, 45.1626281947156, 40.146315971085, 
    47.268851454425, 42.313609019804, 49.0036828201845, 43.7439356159779, 
    51.0619470586162, 45.8676112200792, 40.8716528537064, 47.965109528352, 
    43.0302263684599, 50.0364447368153, 45.1626281947156, 47.268851454425, 
    42.313609019804, 49.0036828201845, 43.7439356159779, 51.0619470586162, 
    45.8676112200792, 40.8716528537064, 47.965109528352, 43.0302263684599, 
    50.0364447368152, 45.1626281947156, 47.268851454425, 42.313609019804, 
    49.0036828201845, 43.7439356159779, 51.0619470586162, 45.8676112200792, 
    40.8716528537064, 47.965109528352, 43.0302263684599, 50.0364447368152, 
    45.1626281947156, 47.268851454425, 42.313609019804, 49.0036828201845, 
    43.7439356159779, 51.0619470586162, 45.8676112200792, 47.965109528352, 
    43.0302263684599, 50.0364447368153, 45.1626281947156, 47.268851454425, 
    42.313609019804, 49.0036828201845, 43.7439356159779, 51.0619470586162, 
    45.8676112200792, 47.965109528352, 43.0302263684599, 50.0364447368152, 
    45.1626281947156, 47.268851454425, 49.0036828201845, 43.7439356159779, 
    51.0619470586162, 45.8676112200792, 47.965109528352, 43.0302263684599, 
    50.0364447368152, 45.1626281947156, 47.268851454425, 49.0036828201845, 
    43.743935615978, 51.0619470586162, 45.8676112200792, 47.965109528352, 
    50.0364447368152, 45.1626281947156, 47.268851454425, 49.0036828201845, 
    43.7439356159779, 51.0619470586162, 45.8676112200792, 47.965109528352, 
    50.0364447368153, 45.1626281947156, 47.268851454425, 49.0036828201845, 
    51.0619470586162, 45.8676112200792, 47.965109528352, 50.0364447368152, 
    45.1626281947156, 47.268851454425, 49.0036828201845, 51.0619470586162, 
    45.8676112200792, 47.965109528352, 50.0364447368152, 47.268851454425, 
    49.0036828201845, 51.0619470586162, 45.8676112200792, 47.965109528352, 
    50.0364447368152, 47.268851454425, 49.0036828201845, 51.0619470586162, 
    45.8676112200792, 47.965109528352, 50.0364447368153, 47.268851454425, 
    49.0036828201845, 51.0619470586162, 47.965109528352, 50.0364447368152, 
    47.268851454425, 49.0036828201845, 51.0619470586162, 47.965109528352, 
    50.0364447368152, 49.0036828201845, 51.0619470586162, 47.965109528352, 
    50.0364447368152, 49.0036828201845, 51.0619470586162, 50.0364447368153, 
    51.0619470586162, 50.0364447368152, 51.0619470586162, 50.0364447368152, 
    51.0619470586162 ;

 obs_Zgrid = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0 ;

 obs_error = 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.169206023673944, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.236255327678716, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.17556760861175, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.223196763845215, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.235533601422048, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.228712343216355, 
    0.235744558228311, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.171836779133628, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.162895037797164, 0.16, 0.16, 0.16, 0.16, 0.16, 0.308477104980401, 
    0.166997650688514, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.420906402871828, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.171623836939502, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.231263474606969, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.255906707668323, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.180739066770684, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.27305871365506, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.210282059700098, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.168947220181749, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.326175480240323, 0.182336397522704, 0.841617820109869, 
    0.366017024386714, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.623906398614281, 0.431207267386656, 0.16, 0.16, 0.16, 
    0.177744377255522, 0.18731242704398, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.344668699428943, 0.16, 0.16, 0.16, 0.1875, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.203616172396576, 
    0.182449070394366, 0.404810133831867, 0.16, 0.740713460286497, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.265203209058028, 0.302222301430447, 
    0.16, 0.16, 0.427500114441024, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.620789541319744, 0.311053361730535, 0.16, 0.225260973199566, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.426319582634096, 0.379140454928221, 
    0.223218806743733, 0.16, 1.12154779706686, 0.16, 1.14083316802983, 0.16, 
    0.16, 0.170368834762154, 0.16, 0.175736671657219, 0.567207416934328, 
    0.51060831967175, 0.203242975359103, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.181969531788809, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.173249823331889, 0.16, 0.196412271437081, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.258867296792914, 0.16, 0.01, 0.01, 0.01, 0.01, 
    0.324375324438734, 0.0121287765138732, 0.038382151443966, 
    0.0240197479604376, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    1.62889755259069, 0.0419550288354458, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0504894010198768, 0.0221785731046111, 0.00233577516773949, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.00138104300034077, 0.0001, 0.01, 0.01, 0.01, 0.01, 1.65763796959436, 
    0.189741286346634, 0.048849569938443, 0.01, 0.0358767342185502, 
    0.058099554037949, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.0001, 0.0001, 0.0001, 0.0001, 0.0017334126799445, 
    0.0272445019581937, 0.0356001375475898, 0.00522243865998462, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.170362611578033, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.231153241230707, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.236314026755609, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.168976922597216, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.236366940216031, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.17166405154689, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.165160361550926, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.425309012322209, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.180274257448211, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.252474126695068, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.259657617495375, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.341411981870082, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.425859563795815, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.189787504936653, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.190438281970163, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.306693419502507, 0.163760513292607, 0.736021128966869, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.623906398614281, 
    0.431207267386656, 0.16, 0.16, 0.16, 0.16, 0.173249955654228, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.317612613250406, 0.16, 
    0.16, 0.16, 0.1875, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.209003817931969, 0.182449070394366, 0.404810133831867, 0.16, 
    0.740713460286497, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.265203209058028, 0.302222301430447, 0.16, 0.16, 0.427500114441024, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.620789541319744, 
    0.311053361730535, 0.16, 0.225260973199566, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.426319582634096, 0.417856958934457, 0.223218806743733, 0.16, 
    1.12154779706686, 0.16, 1.14083316802983, 0.16, 0.16, 0.170368834762154, 
    0.16, 0.175736671657219, 0.556349767466951, 0.51060831967175, 
    0.203242975359103, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.188555043171618, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.173249823331889, 
    0.16, 0.196412271437081, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.17800923363263, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.17775111871942, 0.16, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.01, 
    0.01, 0.01, 0.01, 0.0156910209739181, 0.0438008630647649, 
    0.547292163201109, 0.01, 0.01, 0.0314631155523557, 0.0151807135847169, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.000624001098913141, 
    0.0338037966459524, 0.0263323568316991, 0.00419089860952226, 
    0.000151686307799537, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.01, 0.01, 
    0.0297230925192713, 0.01, 0.01, 0.01, 0.01, 0.24514808984577, 
    0.019256473790154, 0.01, 0.01, 0.01, 0.0154299090933584, 
    0.0226917920130563, 0.0147561568154877, 0.01, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.167758493312198, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.218476031769064, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.253970290586694, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.188556690375325, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.387052559211043, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.22082990681889, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.168922335643806, 0.16, 0.16, 0.16, 0.16, 0.268183449650678, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.262984531641855, 0.16, 0.16, 0.16, 
    0.16, 0.166218503489694, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.197824004295878, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.21219825571601, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.171913918265311, 
    0.175010843616946, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.178992779608507, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.164015345904828, 0.16, 0.16, 0.16, 0.16, 
    0.175879345169278, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.635867754907122, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.172933733402274, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.180385724258734, 
    0.266562116742534, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    1.85281286716463, 0.307151112715443, 0.16, 0.16, 0.16, 0.16, 
    0.173249955654228, 0.16, 0.16, 0.16, 0.16, 0.16, 0.236560948623365, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.433475232442288, 0.16, 0.16, 0.16, 0.1875, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.209003817931969, 0.215377181021369, 
    0.392152663601792, 0.16, 0.740713460286497, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.180353030772818, 
    0.16, 0.16, 0.194176510876754, 0.16, 0.365316369772144, 0.16, 
    0.468000037193633, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.620789541319744, 0.311053361730535, 0.16, 0.225260973199566, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.491905725717697, 0.417856958934457, 
    0.165017488267823, 0.28125, 1.36124937057502, 0.16, 0.16, 
    0.170368834762154, 0.16, 0.175736671657219, 0.556349767466951, 
    0.51060831967175, 0.203242975359103, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.193488433406502, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.173249823331889, 0.16, 0.196412271437081, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.175906727605004, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.164341237621102, 0.16, 0.16, 0.16, 0.240545853331848, 
    0.16, 0.16, 0.16, 0.25061127991992, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.229806806459753, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.0688564273720011, 0.0211968311302344, 0.0321866176903616, 
    0.0439302069940496, 0.0189343745927172, 0.0284255121212581, 
    0.0495865738129722, 0.0279395934441173, 0.0217164937494265, 
    0.113565808354486, 0.0328322511322492, 0.0464301975957755, 
    0.0277489334581181, 0.01, 0.01, 0.01, 0.01, 0.01, 0.0941105779414708, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.0548090222587234, 0.0316542262025905, 0.0148340101627582, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0040500137329218, 
    0.00884493024204858, 0.00414046389778378, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.161494834401866, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.181779190759471, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.204750810126136, 0.16, 0.214176758009671, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.172032629036425, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.234138924188629, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.164342905655177, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.170321954357658, 0.173788603214462, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.411187648673831, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.186857271570489, 0.16, 0.16, 0.16, 
    0.16, 0.280361056149205, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.216000270656145, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.179386209794233, 0.176948346328152, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.170538680574771, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.175471568958549, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.208095779020798, 0.18113227749968, 0.16, 0.16, 
    0.161913314600745, 0.330000085830718, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.255720028948417, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.178928526469723, 0.16, 0.20812522888203, 
    0.16, 0.16, 0.16, 0.619104246457482, 0.403072977860802, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.162498701384215, 0.16, 
    0.181687655925816, 0.16, 0.16, 0.243416638692361, 0.16, 0.16, 
    0.209003817931969, 0.215377181021369, 0.216501779556388, 0.16, 
    0.631827416931044, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.170457777174559, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.203557247767941, 0.16, 
    0.224656370163046, 0.278738629818106, 0.302562340736495, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.620789541319744, 0.311053361730535, 0.16, 
    0.203623897367992, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.247499814033563, 
    0.186749908447382, 0.16, 0.16, 0.16, 0.170368834762154, 0.16, 
    0.175736671657219, 0.556349767466951, 0.51060831967175, 
    0.203242975359103, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.237740099601852, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.173249823331889, 
    0.16, 0.196412271437081, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.170997930777528, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.190835307095182, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.446182357798484, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.170163644763279, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.220951519713526, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.172033131606693, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.181123597304602, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.01, 0.01, 0.01, 0.01, 0.01, 2.22978286072005, 0.01, 
    0.110309041844024, 0.0295305330382689, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.00360850169090554, 0.0001, 0.0438204756792402, 
    0.00819178906385787, 0.0341147000726778, 0.01, 0.01, 0.01, 0.01, 
    1.20238138122841, 0.01, 0.0131558080029208, 0.0694856064951637, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.00145784015330719, 0.0226847665107925, 0.0139444694214035, 
    0.0030419309696299, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.000732873089436909, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.00178545430973173, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.00222919926121832, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0017237827368197, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.000618576550867875, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.00146547146141529, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.00319360671211034, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.00344839172363281, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.00312514992430806, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.00306183930981205, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.00215113790524192, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.000772919896536042, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.000453614406473938, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.000614632743236143, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.000491725297656379, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004 ;

 obs_value = 17.8686498006185, 17.8131071726481, 17.8617830276489, 
    17.6225627263387, 17.1223834355672, 16.9473829269409, 16.7027254104614, 
    16.6388298670451, 16.740306854248, 16.4919951756795, 16.374140103658, 
    16.3761348724365, 16.0612738927205, 15.6583701769511, 15.605455716451, 
    14.8883198102315, 14.4206415812174, 14.3832081158956, 13.8395233154297, 
    13.6499096552531, 13.1701434453328, 13.2680602073669, 13.2600247065226, 
    13.4456125895182, 13.3635026613871, 13.4539214769999, 13.7342659632365, 
    13.0989408493042, 12.7016830444336, 12.7761775652568, 11.9570039113363, 
    11.7327136993408, 11.5222371419271, 11.249197324117, 10.9549608230591, 
    10.781909942627, 10.7043263117472, 10.7628067334493, 10.7439735730489, 
    11.2142833073934, 11.1918082237244, 10.9110434850057, 11.1261164347331, 
    10.8196873664856, 10.6027889251709, 10.2856755256653, 10.4315498669942, 
    9.87392600377401, 9.83848222096761, 9.58017428716024, 9.37397400538127, 
    17.902720981174, 17.7539225684272, 17.6760533650716, 17.5449314117432, 
    17.1177950965034, 16.8860143025716, 16.5799312591553, 16.5810521443685, 
    16.5950130886502, 16.4062904781765, 16.321013768514, 16.3073289659288, 
    16.1882004208035, 15.6307292514377, 15.5051152971056, 15.1281949149238, 
    14.4904933505588, 14.5163915952047, 14.2146603266398, 13.8862502574921, 
    13.6025365193685, 13.6202226479848, 13.5435059865316, 13.5756066640218, 
    13.5631836255391, 13.6322495142619, 13.5650587876638, 12.8016896247864, 
    12.4629538853963, 12.210329691569, 12.2411887645721, 11.8469492594401, 
    11.5793776512146, 11.5222968260447, 11.1392214298248, 10.9604073365529, 
    10.7619397640228, 10.9713776906331, 11.0695140361786, 11.1925318241119, 
    10.9902223745982, 11.0476109981537, 11.0335791905721, 10.7934989134471, 
    10.435835202535, 10.4300451278687, 10.1385598977407, 10.0796749591827, 
    9.62425168355306, 9.66027688980103, 9.58813381195068, 17.6685240003798, 
    17.5441362592909, 17.4093339708116, 17.3339163462321, 17.0588575998942, 
    16.579709370931, 16.4384117126465, 16.5931549072266, 16.5161732567681, 
    16.3779218461778, 16.3396731482612, 16.2868169148763, 16.3915076785617, 
    15.9734265009562, 15.6506340238783, 15.1115172704061, 14.8780102199978, 
    14.8882077534993, 14.7659137248993, 14.3006910483042, 14.0097931226095, 
    13.9310528437297, 13.9156708717346, 13.8826749324799, 13.5762342611949, 
    13.4387756983439, 13.2277731100718, 12.4343460400899, 12.3752910296122, 
    12.377716700236, 12.164178053538, 11.8559877872467, 11.7691961129506, 
    11.718638420105, 11.1890168190002, 11.1178963184357, 11.0474449793498, 
    11.1153093179067, 11.2982345422109, 11.3646145661672, 11.2251887321472, 
    11.0229583581289, 10.6965347131093, 10.7022506395976, 10.3992682298025, 
    10.0641298294067, 9.94975781440735, 9.72301204999288, 9.77265508969625, 
    9.88398782412211, 9.82052246729533, 17.8643211788601, 17.5660885704888, 
    17.3851555718316, 17.1644221411811, 16.8518784840902, 16.4433966742622, 
    16.2801149156358, 16.3657266828749, 16.4109128316243, 16.3826620313856, 
    16.2061865064833, 16.2727419535319, 16.276765399509, 16.0027279324002, 
    15.582453833686, 15.4504129621718, 15.1324907938639, 15.018320719401, 
    14.1425299114651, 13.5889497333103, 13.6990977393256, 14.0432945887248, 
    13.7892492082384, 13.6638476053874, 13.5874565972222, 13.256067276001, 
    12.8657422595554, 12.2033785714044, 12.1095161437988, 11.7979148228963, 
    11.6323902342055, 11.3136403825548, 11.4431229697333, 11.8368631998698, 
    11.263252682156, 11.4188646740384, 11.0170679092407, 11.4953223334418, 
    11.5026312934028, 10.899735238817, 11.153423945109, 10.9864328172472, 
    10.9134111404419, 10.4472222858005, 10.1945996814304, 9.97936598459879, 
    9.60224363538954, 9.62567117479112, 9.86019388834635, 9.98873117234972, 
    9.98170778486464, 18.0199442969428, 17.7590065002441, 17.2391632927789, 
    16.8445248074002, 16.6465733846029, 16.4957205454508, 16.0748896068997, 
    16.2683410644531, 16.3235003153483, 16.2869290245904, 16.1319358613756, 
    16.2453132205539, 16.1663838492499, 15.8937543233236, 15.710226588779, 
    15.5261217753092, 15.2293580373128, 14.3206237157186, 13.3676670392354, 
    13.1091509660085, 13.2072250048319, 13.5499849319458, 13.6086343129476, 
    13.6254851818085, 13.3893189430237, 12.8595005671183, 12.4759302934011, 
    12.338770866394, 11.7873073418935, 11.3035844167074, 11.2414281368256, 
    11.0850691000621, 11.0477206707001, 11.1969409783681, 11.3570636113485, 
    11.1844186782837, 10.8272945086161, 10.9952200253805, 11.0786762237549, 
    10.8792855739594, 10.9872721036275, 10.7128615379333, 10.6246434052785, 
    9.94160429636637, 9.72100361188253, 9.53459604581197, 9.4722912311554, 
    9.65840101242065, 9.6197235584259, 9.88399235407511, 9.98665579160055, 
    17.7009154425727, 17.5789824591743, 17.1332092285156, 16.9326489766439, 
    16.8175843556722, 16.5973731146918, 16.1374693976508, 16.3025512695312, 
    16.2559343973796, 16.1199090745714, 16.0837603674995, 16.0409804450141, 
    15.9943709903293, 15.673135333591, 15.5815919240316, 15.2156396441989, 
    14.5940988328722, 13.59010887146, 13.0655469894409, 12.9491009712219, 
    13.1538377602895, 13.4721104303996, 13.5177763303121, 13.6241952578227, 
    13.3411426544189, 12.5562081336975, 12.2922523021698, 11.9097426732381, 
    11.3092327912649, 11.2333728472392, 11.1744136810303, 11.2402401765188, 
    10.8076803684235, 11.0387280782064, 11.033539613088, 10.934552192688, 
    10.7047639687856, 10.7170461813609, 10.8562707901001, 10.8051074345907, 
    10.6753590901693, 10.5273989836375, 10.0264480908712, 9.84856613477071, 
    9.86593238512675, 9.51769963900248, 9.53892199198405, 9.62269139289856, 
    9.78984610239665, 9.69866625467936, 9.90589157740275, 17.6028116014269, 
    17.6113736894396, 17.3912599351671, 16.8856870863173, 16.8895681169298, 
    16.6807166205512, 16.1919623480903, 16.2148068745931, 16.0463875664605, 
    15.8665758768717, 15.8888018925985, 15.9329424964057, 15.6039623684353, 
    15.4220310846965, 15.4123918745253, 15.0238551033868, 13.74520556132, 
    13.0483843485514, 12.989968723721, 13.1687825520833, 13.3401367399428, 
    13.4320959515042, 13.5714970694648, 13.5118360519409, 13.2521700329251, 
    12.6334020826552, 11.8846242692735, 11.2785120010376, 11.1115425957574, 
    11.2083404329088, 11.1808550092909, 11.3472635481093, 11.0289876725939, 
    10.909107208252, 10.7710780037774, 10.6348027123345, 10.6212383906047, 
    10.7047668033176, 10.9113020367093, 10.8953300052219, 10.6949564615885, 
    10.3004207611084, 9.89880996280246, 10.0633770624797, 10.1181305779351, 
    9.88602574666341, 9.72119808197021, 9.7685522503323, 9.79260084364149, 
    9.20212512546115, 9.40839693281386, 17.7412052154541, 17.6021075778537, 
    17.3496534559462, 16.9679419199626, 16.8956127166748, 16.633267932468, 
    16.2120193905301, 16.1111454433865, 15.7553897433811, 15.7244053946601, 
    15.904599931505, 15.7626298268636, 15.6105767356025, 15.5001724031236, 
    15.0587934917874, 14.551583925883, 13.2095504336887, 12.9099601904551, 
    13.1324632962545, 13.3077109654744, 13.4097334543864, 13.3170934518178, 
    13.3796151479085, 13.2215209007263, 13.102506796519, 12.2115104198456, 
    11.4274423917135, 11.1176384290059, 11.1875011920929, 11.1681145826975, 
    11.2096800804138, 11.2104723453522, 11.1818552017212, 10.8214148680369, 
    10.6481671333313, 10.5365335146586, 10.7371890544891, 10.7612276871999, 
    10.7428054014842, 11.0097764333089, 10.8647513389587, 10.7389195760091, 
    10.3815069993337, 10.0843800703684, 10.2859400908152, 10.0456237792969, 
    9.72928563753764, 9.60072875022888, 9.27522460619609, 9.26683020591736, 
    9.84079869588216, 17.8264122009277, 17.6364163292779, 17.6271606021457, 
    17.259800169203, 16.9632778167725, 16.4979864756266, 16.230035993788, 
    16.0902796851264, 15.8471589618259, 15.8726453781128, 15.7299062940809, 
    14.9159389071994, 15.095788107978, 15.2666282653809, 15.0101013183594, 
    14.0720207426283, 13.042195532057, 12.7828991413116, 13.1682035923004, 
    13.4103170235952, 13.3750964005788, 13.30495540301, 13.3638764222463, 
    13.3633289337158, 12.8981987635295, 11.7944509188334, 11.2285717328389, 
    11.065572977066, 11.2689394950867, 11.3391540845235, 11.2757557233175, 
    11.1330415407817, 11.1177975336711, 10.8609031836192, 10.6383199691772, 
    10.8754473527273, 10.638486067454, 10.6567704677582, 10.6553152402242, 
    10.8320926030477, 10.9443678855896, 10.7345778942108, 10.4634408950806, 
    10.2523949146271, 10.250873486201, 10.0680010318756, 9.79902680714925, 
    9.32157532374064, 8.79749234517415, 9.53988711039225, 10.0852352778117, 
    17.8208457099067, 17.6720951928033, 17.5554358164469, 17.2240113152398, 
    16.7869582706028, 16.3353231218126, 16.3282324473063, 16.1936158074273, 
    16.0250906414456, 15.7660064697266, 15.0044167836507, 14.6308188968235, 
    14.6093427870009, 15.1613915761312, 15.0414596133762, 13.7811891767714, 
    13.0439778433906, 12.5793139139811, 13.0025089051988, 13.3656131956312, 
    13.309105237325, 13.2741913265652, 13.1729532877604, 13.0002508163452, 
    12.6922752592299, 11.6331615447998, 11.0862038930257, 11.0864955054389, 
    11.3518313301934, 11.4748825497097, 11.237471792433, 11.1656413608127, 
    11.1809567345513, 10.7635019090441, 10.631396929423, 10.5984117719862, 
    10.5454712973701, 10.4675868352254, 10.658835305108, 10.8727882173326, 
    11.0236953099569, 10.6267618603177, 10.433439678616, 10.5103601879544, 
    10.0601825714111, 10.017853418986, 10.0602272881402, 9.47212759653727, 
    9.24998537699381, 10.0335140228271, 10.028789308336, 17.806751675076, 
    17.5662708282471, 17.4335505167643, 17.3674023946126, 17.2081707848443, 
    16.6736867692735, 16.5820914374457, 16.3212912877401, 15.848478741116, 
    15.3983489142524, 14.7520723342896, 14.6551904678345, 14.3877025180393, 
    14.4336366653442, 14.5765027999878, 13.442386203342, 13.1544272104899, 
    12.6320009231567, 12.5607833862305, 12.9405498504639, 13.1890299320221, 
    13.1316666603088, 13.0223200321198, 12.882461309433, 12.6328237056732, 
    11.6320850849152, 11.1299397150675, 11.1505583922068, 11.3746054967244, 
    11.6599852244059, 11.3427301247915, 11.5044706662496, 11.2542022864024, 
    11.006786108017, 10.6719636122386, 10.6243744691213, 10.5895075798035, 
    10.4794416427612, 10.8959666093191, 10.7225592931112, 10.5128107070923, 
    10.4009798367818, 10.4326225916545, 10.3359718322754, 10.1406003634135, 
    10.0445350805918, 9.8684667746226, 9.6552050113678, 9.75360989570618, 
    10.2284070650736, 9.95206395785014, 17.4773616790771, 17.439728418986, 
    17.3446824815538, 17.4639818403456, 17.4404021369086, 17.1504692501492, 
    16.7966232299805, 16.2445588641697, 15.6625797483656, 15.131136364407, 
    14.5887150234646, 14.556719356113, 14.2977734671699, 14.0645848380195, 
    13.9321426815457, 13.2347113291423, 13.129828453064, 12.6229612827301, 
    12.5664873917898, 12.5571709473928, 13.017871538798, 12.937243382136, 
    12.8408591747284, 12.8055454889933, 12.4790213108063, 11.7397116820017, 
    11.2407761414846, 11.4613250096639, 11.9286359151204, 12.0463620821635, 
    11.2490148544312, 11.3920844395955, 11.3825311660767, 11.0961714585622, 
    10.8651951948802, 10.6444195906321, 10.7374013264974, 10.5873325665792, 
    10.8382159868876, 10.7148042519887, 10.5115649700165, 10.4034101963043, 
    10.412383556366, 10.3893005847931, 10.2036020755768, 10.0885475476583, 
    9.91014615694682, 9.42600893974304, 10.1750884056091, 10.3201859792074, 
    10.0052728652954, 17.1840029822456, 17.3383384280735, 17.2045665317112, 
    17.2749262915717, 17.3671120537652, 17.2288265228271, 16.6493184831407, 
    16.1576750013563, 15.6531579759386, 14.8095438215468, 14.5511629316542, 
    14.5960733625624, 14.2198066711426, 14.2272093031141, 14.0841466055976, 
    13.3366684383816, 13.1227495405409, 12.7298672993978, 12.9693313174778, 
    12.7153290642632, 12.726454310947, 12.8297713597616, 12.6739433076647, 
    12.6370987362332, 12.3672902848985, 12.1135889689128, 11.854240099589, 
    12.120166460673, 12.30351946089, 12.1950885984633, 11.1856772104899, 
    10.9993022282918, 11.1989393234253, 11.0322364171346, 11.0713130103217, 
    10.6779696146647, 11.0253166622586, 10.9325436486138, 11.0269550747342, 
    11.0111149681939, 10.6976925532023, 10.4212410185072, 10.4820054372152, 
    10.2026970121596, 9.98784690433078, 10.2526546054416, 10.2286703321669, 
    9.81193044450548, 10.3288114335802, 10.1794766320123, 9.80511336856418, 
    16.9263485802544, 17.2302186754015, 17.1730774773492, 17.3546373579237, 
    17.4236189524333, 17.1738957299127, 16.4787108103434, 16.2181760999892, 
    15.8224564658271, 14.8799469206068, 14.6637399461534, 14.6929047902425, 
    14.1821202172173, 14.2238669925266, 14.2059072918362, 13.545115047031, 
    13.1697787178887, 12.8228424390157, 13.2275823752085, 12.9264861742655, 
    12.5462508201599, 12.5235587755839, 12.5382173061371, 12.700515349706, 
    12.7435689767202, 12.7285847663879, 12.533770720164, 11.7227299213409, 
    11.72798426946, 11.5600167115529, 11.0773317813873, 10.9342215061188, 
    10.7637391885122, 10.9474337100983, 10.7288604216142, 10.6729708512624, 
    9.99999986376081, 10.1999998092651, 10.2910713468279, 10.533749961853, 
    10.428658246994, 10.3317415714264, 10.9522763888041, 10.4354976926531, 
    9.99507403373718, 9.85002794265747, 9.3729043006897, 9.74030009183017, 
    9.82614785974676, 9.86240369623358, 9.54256304105123, 16.7831810845269, 
    16.7887465159098, 16.8574470943875, 17.0785927242703, 17.2093717787001, 
    16.8833484649658, 16.4858462015788, 16.1154221428765, 15.9110057618883, 
    15.1512944963243, 14.5927799012926, 14.5875798331367, 14.2906640370687, 
    14.2880047692193, 14.302638053894, 13.6480691697862, 13.4153170055813, 
    12.960916519165, 13.2307871977488, 13.1495540142059, 12.5491460164388, 
    12.3106647332509, 12.3542804718018, 12.4939960638682, 12.8044987519582, 
    12.8055377006531, 12.1909607251485, 11.3653008937836, 11.3768981297811, 
    11.2964475154877, 11.2066859404246, 10.9633156458537, 10.8241041501363, 
    11.0431148355657, 10.6669385433197, 10.5407814184825, 10.1969999313354, 
    10.2910714830671, 10.178750038147, 10.375, 10.2679562568665, 
    10.2842186689377, 9.23125004768372, 9.44553579602923, 9.59716653823853, 
    9.36710691452026, 9.75086291631063, 9.14531254768372, 9.71999988555908, 
    16.8455515967475, 16.670398288303, 16.5924254523383, 16.7193902333577, 
    16.9921724531386, 17.0061558617486, 16.7068116929796, 16.2812455495199, 
    16.0771551132202, 15.2430523766412, 14.8340001636081, 14.5557398266262, 
    14.1941146850586, 14.3197728263007, 14.3050056033664, 13.815357208252, 
    13.453172577752, 13.2799819310506, 13.3244272867839, 13.2742685741848, 
    12.7056620915731, 12.4720680448744, 12.2622829013401, 12.4706433614095, 
    12.721126238505, 12.8023256725735, 11.7744862238566, 11.2716440624661, 
    11.5676364898682, 11.6010559929742, 11.4533996582031, 10.6454860899183, 
    10.9812501271566, 11.2478250927395, 10.8089843988419, 10.6052098274231, 
    10.3124081747872, 10.0362501144409, 11.0500001907349, 10.2791666984558, 
    10.3552083969116, 9.75, 10.1999998092651, 9.75749988555908, 
    9.70666631062826, 9.76518938276503, 9.79342608981662, 10.1500220828586, 
    9.88437521457672, 9.82392480638292, 9.77708339691162, 16.8266201019287, 
    16.6703048282199, 16.5996913909912, 16.5696125030518, 16.730989880032, 
    16.6187121073405, 16.3444904751248, 16.2734188503689, 16.3026496039497, 
    15.3992634879218, 14.9586522844103, 14.4224809010824, 14.101053237915, 
    14.3224902682834, 14.4494726392958, 14.1119792726305, 13.6111681196425, 
    13.430597225825, 13.433385848999, 13.249836842219, 12.7235169410706, 
    12.5479542414347, 12.3736299673716, 12.2824199994405, 12.4724773565928, 
    12.6209418773651, 11.5942851702372, 11.2586677869161, 11.7538615862528, 
    11.7440587679545, 11.3050923877292, 11.4008680184682, 11.0583333969116, 
    11.1414774114435, 10.8548458947076, 9.69999994550433, 9.99892861502511, 
    10.1999998092651, 10.3078126907349, 9.95000004768372, 9.61514854431152, 
    9.60738393995497, 9.91185609499613, 9.77400024731954, 9.18947919209798, 
    9.72964421908061, 9.82457224527995, 9.37186543146769, 16.8794000413683, 
    16.6359712812636, 16.5487177107069, 16.426879035102, 16.366141849094, 
    16.1442111333211, 16.1457302305434, 16.2361077202691, 16.4487692515055, 
    15.7744834687975, 15.3182440863715, 14.1497858895196, 13.9635717603895, 
    14.0594823625353, 13.9738202624851, 13.8740448421902, 13.7653101815118, 
    13.6771697998047, 13.4317735036214, 13.313229004542, 12.7764935493469, 
    12.4558240572611, 12.472663640976, 12.5351433753967, 12.6020941734314, 
    12.4170015652974, 11.7714300950368, 11.5159757932027, 11.6049584547679, 
    10.8580003738403, 11.5541666878594, 11.1625001213767, 10.8682735988072, 
    9.87142876216343, 9.09999990463257, 10.483333269755, 9.8746874332428, 
    9.73693171414462, 9.60545444488525, 9.44629796346029, 8.29400690396627, 
    8.48249777158101, 8.63380159031261, 8.3155323266983, 16.9477994706896, 
    16.7322296566433, 16.7102896372477, 16.4096588558621, 16.2166614532471, 
    16.132671462165, 15.9399919509888, 16.3124287923177, 16.0978140301175, 
    15.7933065626356, 15.2180204391479, 14.1952080196804, 13.8165542814467, 
    13.7741102642483, 13.6997520658705, 13.654659377204, 13.744639078776, 
    13.6563516192966, 13.0154858695136, 12.8971887164646, 12.8131279415554, 
    12.4989048639933, 12.3425937228733, 12.2767884996202, 11.9908799065484, 
    11.9892830318875, 11.7684735192193, 11.604575475057, 8.24499979019165, 
    8.83703136444092, 8.65571673711141, 8.13243993123372, 16.9899828169081, 
    16.9137054019504, 16.7561863793267, 16.5123842027452, 16.3484032948812, 
    16.2034346262614, 16.205540339152, 16.0671242607964, 15.7848572201199, 
    15.2138847774929, 14.6135743459066, 14.1822698381212, 14.0229782528347, 
    13.8245691723294, 13.6361236572266, 13.361542807685, 13.5420999526978, 
    13.6583212216695, 13.0707894166311, 12.8432679971059, 12.6996172269185, 
    12.8230729897817, 12.5431199073792, 12.2545596758525, 11.8099154559049, 
    16.7619681888156, 16.6501060061985, 16.6135035620795, 16.5191546546088, 
    16.3023495144314, 16.1949738396539, 15.6564608679877, 15.0288678275214, 
    14.5090747409397, 14.2524926927355, 14.2437662548489, 14.2262574301826, 
    14.2550700505575, 14.0618057250977, 13.6228618621826, 13.2174592547947, 
    13.3244410620795, 13.5286852518717, 13.0062580903371, 12.7373469670614, 
    12.8005523681641, 12.5572541554769, 12.4020782311757, 12.0418565273285, 
    16.7299904293484, 16.6391531626383, 16.5906564924452, 16.4295488993327, 
    16.1397125456068, 15.9153903325399, 14.9179495705499, 14.4562714894613, 
    14.2276825375027, 14.0060107972887, 14.2044010162354, 14.1288526323107, 
    14.2445563210381, 14.0602705213759, 13.5728641086155, 13.2653001149495, 
    13.2593864864773, 13.3914142184787, 12.9605952368842, 13.0803106096056, 
    12.95032787323, 12.4206313027276, 16.6830965677897, 16.605015012953, 
    16.5303145514594, 16.261223687066, 15.8899359173245, 15.5614006254408, 
    14.3891898261176, 14.2678381601969, 14.1427737341987, 14.0319456524319, 
    14.2769354714288, 14.1349148220486, 14.1219362682766, 14.0160848829481, 
    13.4087260564168, 13.2726073794895, 13.2335738076104, 13.4217456181844, 
    13.3300819396973, 12.8728590806325, 12.6099591255188, 11.7611373901367, 
    16.5453073713515, 16.6594751146105, 16.504063712226, 16.1471852196587, 
    15.7476727167765, 14.9186386532254, 14.2192540698581, 14.2322626113892, 
    14.1901455985175, 14.1077641381158, 14.2853445476956, 14.2372908062405, 
    13.9810821745131, 13.652629216512, 13.3071416219076, 13.1505865520901, 
    13.3366417355008, 13.3675328890483, 13.2597035566966, 12.7523018230091, 
    16.4850802951389, 16.7009355756972, 16.597372478909, 16.4319118923611, 
    15.7308297687107, 15.0302744971381, 14.3462080425686, 14.3078046374851, 
    14.2378835678101, 14.2541847229004, 14.3674765692817, 14.1940219667223, 
    13.9387115902371, 13.4876976013184, 13.3458997938368, 13.3540137608846, 
    13.3433936436971, 13.0555456876755, 12.7493443489075, 16.3583819071452, 
    16.6582137213813, 16.6750068664551, 16.6297707027859, 16.2797036700779, 
    15.6099002626207, 14.688078350491, 14.5009901258681, 14.3117105695936, 
    14.2169443766276, 14.2467801835802, 14.1134147644043, 14.1093176735772, 
    13.8649740219116, 13.7368135452271, 13.5462412304348, 13.1887452602386, 
    16.1676298777262, 16.1829718483819, 16.4308105044895, 16.5501015981038, 
    16.573269950019, 16.4100894927979, 15.6922904120551, 15.0853894551595, 
    14.4374317593045, 14.2810617023044, 13.9479375415378, 13.7754980723063, 
    13.6865578757392, 13.6298183865017, 13.5630769729614, 13.287286567688, 
    16.1440082126194, 15.9405457178752, 16.1725900438097, 16.4159437815348, 
    16.5625470479329, 16.5255928039551, 16.170125219557, 15.4327919218275, 
    14.7020237180922, 14.5902191797892, 14.023085170322, 13.4801154666477, 
    13.3690653906928, 13.3497232860989, 13.1888695822822, 16.2841705746121, 
    15.991359922621, 15.7365686628554, 16.2172402275933, 16.4982920752631, 
    16.4266986846924, 16.2690940433078, 15.7190099292331, 15.2130666308933, 
    14.4114251666599, 13.792090733846, 13.491589334276, 13.1007482210795, 
    13.0359231630961, 16.3576833936903, 16.2014168633355, 15.7058262295193, 
    15.92268731859, 16.3095866309272, 16.1635761260986, 15.9240901735094, 
    15.4498772091336, 14.9578783247206, 14.1020731396145, 13.4668126106262, 
    13.5386196772257, 16.3922928704156, 16.1941201951769, 15.7281476126777, 
    15.588354534573, 15.6562995910645, 15.4005977842543, 14.9456764856974, 
    14.5571029451158, 14.4692549175686, 13.790209558275, 13.5639472007751, 
    13.6707068549262, 16.3683717515733, 16.1618849436442, 15.706549220615, 
    15.5398908191257, 15.2471912172106, 15.008531888326, 14.8845717112223, 
    14.2954171498617, 14.186283853319, 13.6932436625163, 13.7802093823751, 
    13.5170142915514, 16.2615411546495, 16.0834242502848, 15.6941484875149, 
    15.6018696890937, 15.6059975094265, 15.591246287028, 14.6508352491591, 
    14.1529490152995, 13.8686939875285, 13.7975871827867, 13.9659023284912, 
    16.2397570080227, 15.9259145524767, 15.6842571894328, 15.7019195556641, 
    15.767831908332, 15.6611891852485, 14.3862484825982, 14.4069890975952, 
    14.1475509007772, 14.048377778795, 14.0315143267314, 16.093297428555, 
    15.6071000629001, 15.6697368621826, 15.8300728268094, 15.7446065478855, 
    15.4587413999769, 14.7541980743408, 14.6405990388658, 14.4917744530572, 
    14.4027310477363, 14.2200627326965, 15.7957474390666, 15.479488796658, 
    15.4125658671061, 15.6371079550849, 15.1254260804918, 15.0618999269274, 
    15.0161162482368, 14.9064904318915, 14.8707484006882, 14.5494068463643, 
    15.6825097401937, 15.4692361619737, 15.3576439751519, 15.2585238350762, 
    15.0796634886, 15.1348473230998, 14.9781494140625, 15.0079839494493, 
    15.0627092785305, 15.9849858813816, 15.7069696850247, 15.4619029362996, 
    15.2038567860921, 15.2228181627062, 15.2203339470757, 15.061680369907, 
    15.1132759518094, 14.9453402757645, 16.3220885594686, 16.1109341515435, 
    15.9966684977214, 15.5056640836928, 15.4451687071058, 14.9691705703735, 
    14.8884754180908, 14.8138809204102, 16.5040844811334, 16.2422099643283, 
    15.9943749109904, 15.3377110163371, 14.9511218600803, 16.1232522328695, 
    15.9359462526109, 15.467033068339, 14.8854451179504, 13.5994353294373, 
    13.5979795455933, 13.5995578765869, 13.5986251831055, 9.31532955169678, 
    8.70725421905518, 8.33609848022461, 7.74068880081177, 6.13158750534058, 
    5.19000482559204, 4.59018754959106, 4.12346506118774, 3.58884763717651, 
    3.06718969345093, 2.74898195266724, 2.37187910079956, 2.04651880264282, 
    12.3035481770833, 6.71296739578247, 32.5345001220703, 32.5349998474121, 
    32.5349998474121, 32.5354995727539, 32.9124008178711, 33.6688003540039, 
    33.9573997497559, 34.0235992431641, 34.0849990844727, 34.1889991760254, 
    34.298999786377, 34.3860015869141, 34.4630012512207, 34.4879989624023, 
    34.5289993286133, 34.5589981079102, 34.5810012817383, 32.5649998982747, 
    34.0623334248861, 12.7304906845093, 12.7311878204346, 12.7328443527222, 
    12.72651720047, 11.7412452697754, 8.79164543151856, 7.69488296508789, 
    7.55984725952148, 7.06394948959351, 6.39525003433228, 5.37227010726929, 
    4.68950748443604, 4.17570924758911, 3.81572961807251, 3.30136156082153, 
    2.90579581260681, 2.54541397094727, 2.28822183609009, 2.04689741134644, 
    1.84791898727417, 32.5050010681152, 32.5050010681152, 32.5040016174316, 
    32.5034999847412, 32.5343335469564, 32.823600769043, 33.4916000366211, 
    33.8880004882812, 33.9651992797852, 33.9822006225586, 34.0699996948242, 
    34.1269989013672, 34.2529983520508, 34.3610000610352, 34.4519996643066, 
    34.4970016479492, 34.5349998474121, 34.560001373291, 34.5830001831055, 
    34.6030006408691, 17.6937446594238, 17.730001449585, 17.9029378890991, 
    17.4762090047201, 17.0930430094401, 16.9600601196289, 16.7098439534505, 
    16.5314207077026, 16.6710096995036, 16.526294708252, 16.3527167638143, 
    16.3751169840495, 16.0161083539327, 15.5816133817037, 15.2764863967896, 
    14.8742070198059, 14.4290722211202, 14.3898981412252, 13.8408015569051, 
    13.6516863505046, 13.1773961385091, 13.2379206021627, 13.1906150182088, 
    13.4185662269592, 13.3045722643534, 13.426969687144, 13.8271678288778, 
    12.6630237897237, 12.6465126673381, 12.4903418223063, 11.7005270322164, 
    11.6904576619466, 11.4702774683634, 11.1652231216431, 10.91193262736, 
    10.747181892395, 10.5829645792643, 10.586002667745, 10.5524668693542, 
    10.8295833269755, 10.9150748252869, 10.7833188374837, 10.9186166127523, 
    10.6432709693909, 10.5113304456075, 10.2855242093404, 10.1239002545675, 
    9.7872314453125, 9.7298747698466, 9.59417994817098, 9.1812268892924, 
    17.8198748694526, 17.6392057206896, 17.5643804338243, 17.5420337253147, 
    17.0952847798665, 16.8775628407796, 16.6725476582845, 16.5505373213026, 
    16.5457897186279, 16.4281154208713, 16.343317243788, 16.3123306698269, 
    16.1716673109267, 15.6803780661689, 15.5035287009345, 15.1462027231852, 
    14.5049866570367, 14.5207765897115, 14.2151068051656, 13.8870411713918, 
    13.5750086307526, 13.5723111629486, 13.5509833494822, 13.4924126466115, 
    13.5302048524221, 13.5381878217061, 13.4089523156484, 12.5501164595286, 
    12.3746281464895, 12.2436544895172, 11.954217672348, 11.7154717445374, 
    11.490690946579, 11.5040876865387, 11.0936754544576, 10.8819674650828, 
    10.6620230674744, 10.7876935005188, 10.8478193283081, 10.9172400633494, 
    10.8042500019073, 10.8612916469574, 10.8216832478841, 10.6228350798289, 
    10.3714328606923, 10.3506693840027, 10.0106611251831, 9.81047145525614, 
    9.44192910194397, 9.50626516342163, 9.41678277651469, 17.5836211310493, 
    17.4016123877631, 17.3076881832547, 17.2938783433702, 17.0205296410455, 
    16.5892908308241, 16.444886525472, 16.4671819474962, 16.4605950249566, 
    16.3788876003689, 16.358287387424, 16.2349806891547, 16.3441537221273, 
    15.967924118042, 15.6431670718723, 15.106320699056, 14.8781006071303, 
    14.8887236913045, 14.7658449014028, 14.3005955219269, 13.992699543635, 
    13.8920055230459, 13.9328811168671, 13.8702554702759, 13.563724120458, 
    13.3598176638285, 13.1823342641195, 12.3871296246847, 12.4543976783752, 
    12.3695323467255, 12.1202133496602, 11.8451909224192, 11.7435890038808, 
    11.7068467140198, 11.1854019959768, 11.100014368693, 11.0835076967875, 
    11.0870052178701, 11.290478626887, 11.2015292644501, 10.602162361145, 
    10.6968416372935, 10.5739465554555, 10.5508950551351, 10.2892010211945, 
    10.0159233411153, 9.88308580716451, 9.47754645347595, 9.54642979303996, 
    9.60847687721252, 9.59736084938049, 17.8578737046983, 17.4757580227322, 
    17.3423444959852, 17.136117723253, 16.8266557057699, 16.4237306382921, 
    16.2261781692505, 16.3233759138319, 16.3644104003906, 16.4055105845133, 
    16.2233325110541, 16.1807969411214, 16.2578639984131, 15.9792802598741, 
    15.5553878148397, 15.4405717849731, 15.1334377924601, 15.018320719401, 
    14.1424502266778, 13.5896589491102, 13.6089785893758, 14.0257547166612, 
    13.7773008346558, 13.6662279764811, 13.5769941541884, 13.2475368711683, 
    12.8621546427409, 12.1886682510376, 12.1545068952772, 11.7826271057129, 
    11.4144153594971, 11.2593588299221, 11.4101370705499, 11.8091465632121, 
    11.2342240015666, 11.3353686862522, 11.0408602820502, 11.5133555730184, 
    11.5053944057888, 10.8783693313599, 10.9018621444702, 10.7666864395142, 
    10.5701333151923, 10.2417536841498, 10.0768080817329, 9.78638490041097, 
    9.40688652462429, 9.40613248613146, 9.59667587280273, 9.64232455359565, 
    9.70053556230333, 18.0488764444987, 17.6874226464166, 17.2139708201091, 
    16.7603969573975, 16.5977562798394, 16.5083401997884, 15.9480610953437, 
    16.1968622207642, 16.2883911132812, 16.2963922288683, 16.1492309570312, 
    16.238774617513, 16.1791896820068, 15.8920379214817, 15.6881240208944, 
    15.512035369873, 15.2317394680447, 14.3131673336029, 13.3686785697937, 
    13.0937016010284, 13.1980386575063, 13.5436470508575, 13.6028870741526, 
    13.6169222195943, 13.3935787677765, 12.8424541950226, 12.4858194986979, 
    12.1658274332682, 11.6716759204865, 11.2865296999613, 11.1014885107676, 
    10.9867877960205, 10.9677430788676, 11.1730676492055, 11.2838368415833, 
    11.2536792755127, 10.9494264125824, 11.0426816940308, 11.1063735485077, 
    10.8888674577077, 10.8158638477325, 10.4961854616801, 10.2884578704834, 
    9.84350482622782, 9.5776302019755, 9.37283190091451, 9.34943087895711, 
    9.41421914100647, 9.58926304181417, 9.63160339991252, 9.64310669898987, 
    17.7513412899441, 17.5036349826389, 17.0402200486925, 16.8896609412299, 
    16.7908520168728, 16.6004967159695, 16.1334100299411, 16.2982090844048, 
    16.2104697757297, 16.124932607015, 16.0962270100911, 16.0330641004774, 
    16.0026455985175, 15.6726339128282, 15.5646432240804, 15.1958654191759, 
    14.5252039167616, 13.5518030325572, 13.0654783248901, 12.937236626943, 
    13.1541740894318, 13.4190465609233, 13.46657594045, 13.5723748207092, 
    13.3312193552653, 12.5441193580627, 12.232275724411, 11.79958264033, 
    11.2710422674815, 11.209298213323, 11.0212182998657, 11.0891395409902, 
    10.7412243684133, 10.9143273830414, 11.004249493281, 11.1027876536051, 
    10.9007859230042, 10.8055682182312, 10.8819371859233, 10.7995351950328, 
    10.7382980982463, 10.328110853831, 9.85271469751994, 9.7894766330719, 
    9.698619445165, 9.43217730522156, 9.41277432441711, 9.49573953946432, 
    9.66675964991252, 9.64011073112488, 9.58169007301331, 17.6035073598226, 
    17.5943400065104, 17.3976018693712, 16.8465008205838, 16.9019198947483, 
    16.6852887471517, 16.191753493415, 16.2127687666151, 15.9862818188137, 
    15.8714865578545, 15.8788563410441, 15.9447668923272, 15.5844176610311, 
    15.4065341949463, 15.3983361985948, 15.0272776285807, 13.7392331229316, 
    13.0319796668159, 12.9851797951592, 13.159310552809, 13.3343562020196, 
    13.3898849487305, 13.5241437488132, 13.4872890048557, 13.2164336310493, 
    12.5225928624471, 11.7971421347724, 11.2028819190131, 11.0694305631849, 
    11.1828544404772, 11.1338216993544, 11.1642991171943, 10.9823678334554, 
    10.6853509479099, 10.6373866399129, 10.6441168255276, 10.6786989635891, 
    10.7393777635362, 10.8137979507446, 10.881268925137, 10.6596859825982, 
    10.1933857599894, 9.86532274881999, 9.92752022213406, 9.92485374874539, 
    9.75587452782525, 9.58518674638536, 9.6163420147366, 9.5298408932156, 
    9.55176226298014, 9.59445646074083, 17.8232216305203, 17.7993960910373, 
    17.4004737006293, 16.9378689659966, 16.8744475046794, 16.6244667900933, 
    16.2127684487237, 16.1646341747708, 15.6907200283474, 15.7386397255792, 
    15.8974473741319, 15.7422457800971, 15.5820118586222, 15.4756342569987, 
    15.0400630103217, 14.5560195710924, 13.2131905025906, 12.8973366419474, 
    13.1204452514648, 13.2991565068563, 13.4008554617564, 13.3070964813232, 
    13.3286213080088, 13.1996954282125, 13.053169965744, 12.2082912127177, 
    11.3724638621012, 11.0728227297465, 11.1757430235545, 11.1569720109304, 
    11.1440397898356, 11.1022510528564, 11.1525371869405, 10.7519336541494, 
    10.537723382314, 10.5064031283061, 10.7146492799123, 10.7242278258006, 
    10.606997013092, 11.0008883476257, 10.8405505021413, 10.665420850118, 
    10.175589799881, 9.94765988985697, 10.0212404727936, 9.86375157038371, 
    9.66036359469096, 9.64508748054504, 9.30817635854085, 9.48144205411275, 
    9.91018295288086, 17.9198691050212, 17.6129336886936, 17.6962846120199, 
    17.1957715352376, 17.0172687106662, 16.5033164554172, 16.2304840087891, 
    16.1439954969618, 15.8119518491957, 15.8972210354275, 15.70753426022, 
    14.8973132239448, 15.0877508587307, 15.2614866892497, 15.0096100701226, 
    14.0767629411485, 13.0367517471313, 12.7686416308085, 13.1524867216746, 
    13.4040497144063, 13.381637096405, 13.3032680352529, 13.3224405447642, 
    13.3534615039825, 12.8783390522003, 11.804424683253, 11.1811677614848, 
    11.0586311022441, 11.3020377159119, 11.3470168908437, 11.2274162769318, 
    11.1118377049764, 11.1096940835317, 10.842182079951, 10.6069476604462, 
    10.8009316126506, 10.552343527476, 10.4983580907186, 10.6097234884898, 
    10.8122088909149, 10.9093942642212, 10.68412510554, 10.2358697255452, 
    10.0641175111135, 9.99645884831746, 9.8703285853068, 9.74492979049683, 
    9.42668867111206, 9.14692068099976, 9.47405815124512, 10.0737017790476, 
    17.8784493340386, 17.725341796875, 17.5648905436198, 17.2703062693278, 
    16.694860458374, 16.2659132215712, 16.3099185095893, 16.2484171125624, 
    16.0808562172784, 15.795166015625, 14.9516269895766, 14.6167897118462, 
    14.6110917197333, 15.1670979393853, 15.0547364552816, 13.788050227695, 
    13.0440475675795, 12.5728293524848, 12.9914990531074, 13.3674942652384, 
    13.3184143702189, 13.2921698888143, 13.175066947937, 13.0230136447483, 
    12.6941702100966, 11.6363002989027, 11.0365765889486, 11.0892339282566, 
    11.3495619032118, 11.4744086795383, 11.1871983210246, 11.1445175806681, 
    11.1997865041097, 10.767770131429, 10.6248502731323, 10.5768300162421, 
    10.5051353242662, 10.4831972122192, 10.6759746339586, 10.84071720971, 
    10.9569389555189, 10.5881834030151, 10.3544262780084, 10.3075529734294, 
    9.92250156402588, 9.79712581634521, 9.97758928934733, 9.52689711252848, 
    9.30525557200114, 9.90899011823866, 9.98599296145969, 17.8575579325358, 
    17.5838911268446, 17.5293602413601, 17.1865906185574, 17.177942276001, 
    16.6429621378581, 16.4565052456326, 16.3173242145114, 15.8799634509616, 
    15.4684620963203, 14.7323178185357, 14.6386131710476, 14.3932049009535, 
    14.4424351586236, 14.589706103007, 13.4534349441528, 13.1558331383599, 
    12.6311225891113, 12.5563387870789, 12.9378110567729, 13.1962159474691, 
    13.1397460301717, 13.0272949536641, 12.8885877927144, 12.6423428853353, 
    11.6248348553975, 11.0736499627431, 11.1259814898173, 11.4179697036743, 
    11.6311333179474, 11.3230783939362, 11.5112370649974, 11.2563999493917, 
    11.0130527814229, 10.7334837118785, 10.672067006429, 10.5905209382375, 
    10.5231002966563, 10.9278486569722, 10.6903898715973, 10.4878570238749, 
    10.3676682313283, 10.353929678599, 10.2997822761536, 10.0132249991099, 
    9.90369002024333, 9.89982096354167, 9.60605986913045, 9.69349964459737, 
    10.1795384089152, 9.95627236366272, 17.4917736053467, 17.4664827982585, 
    17.427858988444, 17.3796819051107, 17.4359192318386, 17.1134018368191, 
    16.8423716227214, 16.2502483791775, 15.6992734273275, 15.1520607206557, 
    14.5940441555447, 14.5505153867933, 14.302891837226, 14.0680945714315, 
    13.9383125305176, 13.2382972505358, 13.1347823672824, 12.6253323554993, 
    12.5671638647715, 12.5567539532979, 13.0168108145396, 12.9289659659068, 
    12.8320221106211, 12.8042879899343, 12.491091410319, 11.7960019906362, 
    11.2173762321472, 11.4647114276886, 11.9478599230448, 12.2364477316538, 
    11.2483568986257, 11.3553188641866, 11.3606896400452, 11.1350758075714, 
    10.965448141098, 10.7341481844584, 10.7847356001536, 10.6277194023132, 
    10.8504501183828, 10.6708690325419, 10.4891974131266, 10.3830798467, 
    10.3069052696228, 10.2867267926534, 9.99286468823751, 9.89801359176636, 
    9.98685932159424, 9.39051556587219, 10.1737484137217, 10.2835642496745, 
    10.0157055854797, 17.1913159688314, 17.3917713165283, 17.2457093132867, 
    17.288361231486, 17.3820669386122, 17.1072118547228, 16.7282307942708, 
    16.1454696655273, 15.5512924194336, 14.815819952223, 14.5415954589844, 
    14.5863242679172, 14.2200298309326, 14.230518023173, 14.0888669755724, 
    13.3389869266086, 13.1271486282349, 12.7360253863864, 12.9757295184665, 
    12.7225756115384, 12.7328098085192, 12.8271376291911, 12.6503926383124, 
    12.6276279025608, 12.3777878019545, 12.1371737586127, 11.7804435094198, 
    12.094886885749, 12.3164033889771, 12.221930609809, 11.1599800321791, 
    10.9656209945679, 11.174190097385, 10.9967477586534, 11.1361507839627, 
    10.732189072503, 11.0445665783352, 10.9317961798774, 11.0215794245402, 
    10.9545832739936, 10.6683674918281, 10.4168854819404, 10.4643559985691, 
    10.1686414082845, 9.97388044993083, 10.041015625, 9.90664037068685, 
    9.69203588697645, 10.3209598329332, 10.1847699483236, 9.81614759233263, 
    16.9579802619086, 17.2916526794434, 17.2281307644314, 17.4965534210205, 
    17.4044592115614, 17.1574242909749, 16.4474059210883, 16.1636621687147, 
    15.7707703908285, 14.8302983178033, 14.627046585083, 14.648770014445, 
    14.1851296954685, 14.2288015153673, 14.2114686965942, 13.5477084053887, 
    13.1695155037774, 12.8259863853455, 13.2424849669139, 12.953651825587, 
    12.5603220462799, 12.5214128494263, 12.5291795730591, 12.701931476593, 
    12.7497297128042, 12.720405737559, 12.4349336624146, 11.6567958990733, 
    11.7119430700938, 11.5628360112508, 11.086980899175, 10.9215311209361, 
    10.7400667667389, 10.9284597237905, 10.7274704846469, 10.6769940853119, 
    9.99999986376081, 10.1999998092651, 10.3875000476837, 10.533749961853, 
    10.428658246994, 10.3270554542542, 10.8476403554281, 10.3791363579886, 
    9.9888870716095, 9.83368062973022, 9.34434620539347, 9.67870911684903, 
    10.1049786567688, 9.86479715867476, 9.54644044240316, 16.8101618025038, 
    16.8340515560574, 16.8954230414497, 17.0987381405301, 17.0843221876356, 
    16.6996739705404, 16.4336982303196, 15.9715741475423, 15.8004233042399, 
    15.0859494739109, 14.532747692532, 14.5420604281955, 14.2711844974094, 
    14.2711011038886, 14.2851909001668, 13.6191870371501, 13.3917134602865, 
    12.9598387082418, 13.2413777510325, 13.1666126251221, 12.5602582295736, 
    12.3210634390513, 12.362070719401, 12.4999029636383, 12.8081270853678, 
    12.8076260884603, 12.1857833067576, 11.3487754662832, 11.3504402637482, 
    11.2916509310404, 11.2155196666718, 10.9667645295461, 10.8280895551046, 
    11.1761148626154, 10.672611951828, 10.5407814184825, 10.1969999313354, 
    10.2910714830671, 10.197500038147, 10.375, 10.2679562568665, 
    10.2842186689377, 9.23125004768372, 9.44553579602923, 9.60299987792969, 
    9.40031266212463, 9.75086291631063, 9.67499987284342, 9.70499992370605, 
    16.8869599236382, 16.7085613674588, 16.6881190405952, 16.7675493028429, 
    16.9711772070991, 16.7388899061415, 16.5291025373671, 16.2812351650662, 
    15.8937301635742, 15.1891639497545, 14.7872800827026, 14.5336057874891, 
    14.1863159603543, 14.3047397401598, 14.2858152389526, 13.7970335218641, 
    13.4382271236844, 13.2771546045939, 13.34112962087, 13.2800630993313, 
    12.7100060780843, 12.4916163550483, 12.2745282914903, 12.4712777667575, 
    12.721126238505, 12.8023256725735, 11.7744862238566, 11.2545075946384, 
    11.5732632742988, 11.6051670710246, 11.3573787477281, 10.5458994971381, 
    10.8525001525879, 11.2906250423855, 10.8532552719116, 10.6052098274231, 
    10.3124081747872, 10.0362501144409, 11.0500001907349, 10.2791666984558, 
    10.3552083969116, 9.75, 10.1999998092651, 9.75749988555908, 
    9.70666631062826, 9.76518938276503, 9.78986114925808, 10.1500220828586, 
    9.88437521457672, 9.82392480638292, 9.77708339691162, 16.8460528055827, 
    16.6969028049045, 16.6693053775364, 16.6027007632785, 16.8233432769775, 
    16.4415020412869, 16.0996532440186, 16.230062590705, 16.2292363908556, 
    15.3381661309136, 14.9258574379815, 14.3943520651923, 14.0936975479126, 
    14.3146342171563, 14.4334565268623, 14.0916333728366, 13.6051068835788, 
    13.432475010554, 13.4415332476298, 13.2520198822021, 12.749720176061, 
    12.5567207336426, 12.3796145121257, 12.2824199994405, 12.4724773565928, 
    12.6209418773651, 11.5978225866954, 11.2709999879201, 11.7634595235189, 
    11.7419753869375, 11.3050923877292, 11.4008680184682, 11.0583333969116, 
    11.1414774114435, 10.8548458947076, 9.69999994550433, 9.99892861502511, 
    10.1999998092651, 10.3078126907349, 9.95000004768372, 9.61514854431152, 
    9.58363395267063, 9.91185609499613, 9.77400024731954, 9.18947919209798, 
    9.72964421908061, 9.82457224527995, 9.37186543146769, 16.9208236270481, 
    16.6820299360487, 16.5760112338596, 16.4555568695068, 16.3555111355252, 
    16.1306425730387, 16.0809540218777, 16.3536508348253, 16.5325609842936, 
    15.6816308763292, 15.2450415293376, 14.1262573666043, 13.9475469589233, 
    14.0432411829631, 13.9594891866048, 13.8594152662489, 13.7654229270087, 
    13.6826733748118, 13.4467675685883, 13.3324186007182, 12.8468386332194, 
    12.4868791898092, 12.472663640976, 12.5351433753967, 12.6020941734314, 
    12.4170015652974, 11.8058098951975, 11.5054933230082, 11.5939283370972, 
    10.8580003738403, 11.6250001192093, 11.1625001213767, 10.8682735988072, 
    9.87142876216343, 9.09999990463257, 10.483333269755, 9.8746874332428, 
    9.73693171414462, 9.60545444488525, 9.44629796346029, 8.29400690396627, 
    8.50310778617859, 8.63380159031261, 8.3155323266983, 16.9304105970595, 
    16.7285346984863, 16.718334197998, 16.3896410200331, 16.1789390775892, 
    16.1237291759915, 15.8911561965942, 16.1852672364977, 16.0732000139025, 
    15.7409620285034, 15.2056303024292, 14.1742097006904, 13.7991377512614, 
    13.7555203967624, 13.6778740353054, 13.6212106280857, 13.7321102354262, 
    13.7196203867594, 13.1563532087538, 13.0029147466024, 12.8011322021484, 
    12.4927955203586, 12.3390264511108, 12.2767884996202, 11.9908799065484, 
    11.9892830318875, 11.7705237070719, 11.604575475057, 8.24499979019165, 
    8.83703136444092, 8.65571673711141, 8.13243993123372, 16.9150602552626, 
    16.8731257120768, 16.7148259480794, 16.4834679497613, 16.3424186706543, 
    16.1645090315077, 16.1189714007907, 16.0495785607232, 15.8201479381985, 
    15.2510902616713, 14.5936047236125, 14.1666332880656, 14.0119410620795, 
    13.8103545506795, 13.5956364737617, 13.3327444924249, 13.5320729149712, 
    13.6787450313568, 13.1607396602631, 12.8429358800252, 12.6888354619344, 
    12.8184821605682, 12.5547772248586, 12.2545596758525, 11.8099154559049, 
    16.6500432756212, 16.5723567538791, 16.5567027197944, 16.4666697184245, 
    16.2542209625244, 16.1898556815253, 15.6560639275445, 14.9813301298353, 
    14.5080601374308, 14.2438420189752, 14.205491065979, 14.1945614284939, 
    14.2472356160482, 14.0375741322835, 13.5961010191176, 13.1873145633274, 
    13.3213895161947, 13.5384578704834, 13.0494287014008, 12.7496828238169, 
    12.7807025114695, 12.5487875143687, 12.4100335439046, 12.0418565273285, 
    16.7167063819038, 16.6062689887153, 16.5582692888048, 16.390574561225, 
    16.1514792972141, 15.9296471277873, 14.8804454803467, 14.4534637663099, 
    14.2308008405897, 14.0397000842624, 14.227807574802, 14.1478486590915, 
    14.222783724467, 14.0418914159139, 13.544380929735, 13.2363941404555, 
    13.2634728749593, 13.4129254023234, 12.9704467985365, 13.0891261630588, 
    12.9389547771878, 12.4134928385417, 16.7234944237603, 16.6337297227648, 
    16.5562148623996, 16.251942952474, 15.9043377770318, 15.5893025928073, 
    14.388891643948, 14.289000193278, 14.1575982835558, 14.0553369522095, 
    14.2832481596205, 14.1568938361274, 14.1120427449544, 14.0046656926473, 
    13.3942487504747, 13.2395684983995, 13.2389114167955, 13.4611438115438, 
    13.3420360883077, 12.8663490613302, 12.5922852357229, 11.767521572113, 
    16.5187507205539, 16.6738529205322, 16.5254272884793, 16.1311232248942, 
    15.705591307746, 14.8826036453247, 14.2167616950141, 14.2471878263685, 
    14.2252396477593, 14.1434471342299, 14.3034642537435, 14.2403863271077, 
    13.9984793133206, 13.660028245714, 13.302926381429, 13.1349129147, 
    13.3327792485555, 13.3654622236888, 13.254326581955, 12.7463287006725, 
    16.4282684326172, 16.7031091054281, 16.6201962365044, 16.3743000030518, 
    15.7320693333944, 14.9624101850722, 14.3652086257935, 14.3763501909044, 
    14.2819900512695, 14.2773803075155, 14.357508553399, 14.1819967693753, 
    13.9337762196859, 13.5071983337402, 13.3438786400689, 13.3531330956353, 
    13.3523423936632, 13.0436960458755, 12.7420965433121, 16.3700389862061, 
    16.6647330390082, 16.6897926330566, 16.6506565941705, 16.230073928833, 
    15.5506753921509, 14.8662859598796, 14.6224585639106, 14.4423459370931, 
    14.3043140835232, 14.2257910834418, 14.1017989052667, 14.0819370481703, 
    13.8633456759983, 13.7263580958048, 13.5428926679823, 13.1832609176636, 
    16.1560103098551, 16.1870237986247, 16.4139876895481, 16.5496135287815, 
    16.597290886773, 16.4025463528103, 15.7143149905735, 15.2816406885783, 
    14.548161400689, 14.4151511722141, 14.0122577879164, 13.7738244798448, 
    13.6713432735867, 13.6146290037367, 13.5428795284695, 13.2911334991455, 
    16.1948632134332, 15.9619491365221, 16.1278898451063, 16.4467860327827, 
    16.5890375773112, 16.6035957336426, 16.190395143297, 15.6050075954861, 
    14.7484658559163, 14.6686903635661, 14.1396536297268, 13.4697051578098, 
    13.3605552249485, 13.3454692628649, 13.1741477118598, 16.3400446573893, 
    16.0223497814602, 15.7546922895643, 16.2794257269965, 16.5503819783529, 
    16.4987733629015, 16.3173364003499, 15.8189455668132, 15.2600491841634, 
    14.4556562635634, 13.8633808559842, 13.4991920259264, 13.096159140269, 
    13.0249026616414, 16.370738559299, 16.2104663848877, 15.7471460766262, 
    16.0429756376478, 16.3412776523166, 16.1532973183526, 15.8721218109131, 
    15.4567687776354, 15.0524798499213, 14.1434533860948, 13.4882436990738, 
    13.5612008836534, 16.4268656836616, 16.2122660742866, 15.7546354929606, 
    15.6148114734226, 15.6239806281196, 15.3284576204088, 14.9734172821045, 
    14.699456108941, 14.6190871132745, 13.9916317198012, 13.6137543916702, 
    13.6740821202596, 16.399057176378, 16.2187564637926, 15.7605288823446, 
    15.565821117825, 15.2564761903551, 15.0411933263143, 14.8318073484633, 
    14.3370991812812, 14.254535039266, 13.741199069553, 13.8378376960754, 
    13.5181556277805, 16.2690987057156, 16.0941608217027, 15.7425896326701, 
    15.6051549911499, 15.6006045871311, 15.5933791266547, 14.6668214797974, 
    14.3171984354655, 14.0433803134494, 13.9103853437636, 14.006888601515, 
    16.2057395511203, 15.8962050543891, 15.7133515675863, 15.718627081977, 
    15.767907778422, 15.7143564224243, 14.4076065487332, 14.4246826171875, 
    14.2096020380656, 14.1505030526055, 14.1717019081116, 16.0270653830634, 
    15.5376519097222, 15.7218840916952, 15.859214146932, 15.7409678565131, 
    15.4992487165663, 14.79220061832, 14.6972401936849, 14.540459950765, 
    14.4677571190728, 14.2809767723083, 15.7460888756646, 15.4975696139865, 
    15.4366044998169, 15.6886438793606, 15.1006814108955, 15.0863129297892, 
    15.0219135284424, 14.9261100557115, 14.89275431633, 14.6215642293294, 
    15.6736613379584, 15.5040584140354, 15.3619737625122, 15.3058924145169, 
    15.091618431939, 15.1621013217502, 15.0464191436768, 15.018789185418, 
    15.0707364612155, 15.9488146040175, 15.7705305947198, 15.5051981608073, 
    15.2187773386637, 15.2492617501153, 15.2279349433051, 15.1302349302504, 
    15.1409287982517, 14.9575517177582, 16.3364404042562, 16.1462031470405, 
    16.0858464770847, 15.5420289569431, 15.5157400767008, 14.9886971579658, 
    14.8799578802926, 14.7411727905273, 16.5501147376166, 16.2896082136366, 
    16.0546145968967, 15.3607108857897, 14.9214821921455, 16.1607813305325, 
    15.9212759865655, 15.5850780275133, 14.9529047012329, 13.660737991333, 
    13.6543226242065, 13.6519346237183, 13.6475734710693, 13.5557880401611, 
    12.320969581604, 10.9682931900024, 9.3370189666748, 9.09381484985352, 
    8.71106433868408, 7.90615367889404, 7.44208955764771, 6.51879835128784, 
    6.36768102645874, 5.95759439468384, 5.44174098968506, 5.31588220596313, 
    5.07773685455322, 4.81876945495605, 4.48915863037109, 4.3190770149231, 
    4.09442853927612, 3.94832134246826, 33.0390014648438, 33.0410003662109, 
    33.0419998168945, 33.0429992675781, 33.0460014343262, 33.1069984436035, 
    33.4220008850098, 33.6570014953613, 33.9179992675781, 34.0260009765625, 
    34.0579986572266, 34.1319999694824, 34.1189994812012, 34.226001739502, 
    34.2350006103516, 34.306999206543, 34.3440017700195, 34.3549995422363, 
    34.3779983520508, 34.4150009155273, 34.4290008544922, 34.4309997558594, 
    34.4529991149902, 11.9808597564697, 11.979567527771, 11.9672937393188, 
    11.8038272857666, 11.5040793418884, 11.1912132898966, 8.86040439605713, 
    7.94273729324341, 7.68683080673218, 7.27129459381104, 6.4627062479655, 
    5.905433177948, 4.96015405654907, 4.36980199813843, 3.99167037010193, 
    3.61798858642578, 3.20025634765625, 2.93255996704102, 2.66319346427917, 
    2.38115048408508, 2.12302207946777, 2.01422190666199, 1.83520793914795, 
    32.609001159668, 32.6080017089844, 32.6049995422363, 32.5929985046387, 
    32.5665016174316, 32.5890007019043, 32.863200378418, 33.4963996887207, 
    33.8833999633789, 33.9877998352051, 34.0226669311523, 34.0349998474121, 
    34.1080017089844, 34.1699981689453, 34.2569999694824, 34.3660011291504, 
    34.423999786377, 34.4700012207031, 34.5040016174316, 34.5349998474121, 
    34.5610008239746, 34.576000213623, 34.5909996032715, 8.24374903165377, 
    8.07208486703726, 7.40963862492488, 10.1993227005005, 10.1984163920085, 
    10.1972808837891, 10.1961441040039, 9.74515962600708, 8.72219058445522, 
    8.59093364079793, 8.52049914995829, 8.14381901423136, 7.83411924044291, 
    6.89342304070791, 6.35731637477875, 6.05581331253052, 17.4521064758301, 
    17.5186147689819, 17.7798026402791, 17.2524731953939, 16.8908859888713, 
    16.841423034668, 16.6067616144816, 16.4914929072062, 16.4654572804769, 
    16.3707898457845, 16.310320854187, 16.2978836695353, 15.9055972099304, 
    15.5073030789693, 15.2727502187093, 14.7865436871847, 14.3055931727091, 
    14.2342782020569, 13.8623596827189, 13.5598425865173, 13.2206937472026, 
    13.1862414677938, 13.1362455685933, 13.1925018628438, 13.2313092549642, 
    13.3542019526164, 13.3689521153768, 12.9612310727437, 12.3907348314921, 
    11.9085378646851, 11.7606477737427, 11.8396237691243, 11.6014156341553, 
    11.2889803250631, 11.0234769185384, 10.8983608881632, 10.5983700752258, 
    10.7106485366821, 10.7239500681559, 10.8712759017944, 10.4368408521016, 
    10.269420782725, 10.5252105394999, 10.2006138165792, 10.1269243558248, 
    9.92950487136841, 9.83324750264486, 9.70593372980754, 9.47948582967122, 
    9.28510999679565, 8.92641830444336, 17.6219306521946, 17.4285803900825, 
    17.6011778513591, 17.4277763366699, 16.9896969265408, 16.806791305542, 
    16.5446597205268, 16.4778535630968, 16.4132408565945, 16.3403911590576, 
    16.3200971815321, 16.301718182034, 16.0416741900974, 15.5963178210788, 
    15.4450531005859, 14.9978722466363, 14.3880194558038, 14.4419848124186, 
    14.050444761912, 13.7898867925008, 13.550878127416, 13.4420030117035, 
    13.3393286863963, 13.3702449798584, 13.4143737951914, 13.3680259386698, 
    13.3220423857371, 12.8759008248647, 12.3103707631429, 12.0574643611908, 
    11.7251416842143, 11.6445637543996, 11.4323325157166, 11.4365921815236, 
    11.1384031772614, 10.8755568663279, 10.7099364598592, 10.8574593861898, 
    11.0625181992849, 11.0488599141439, 10.765119155248, 10.4057608445485, 
    10.4253056049347, 10.3070116837819, 10.070229212443, 9.99454148610433, 
    9.66588393847148, 9.56306902567546, 9.2147487004598, 9.27773412068685, 
    9.13771017392476, 17.4306439293755, 17.100271013048, 17.2871918148465, 
    17.294442070855, 16.9547742207845, 16.5289906395806, 16.3720082177056, 
    16.4089387257894, 16.343271891276, 16.2679996490479, 16.2781829833984, 
    16.1842695871989, 15.917549027337, 15.7824754714966, 15.5193818410238, 
    15.1113849216037, 14.7047296100193, 14.6815431118011, 14.4707549413045, 
    14.1779828866323, 13.9392410119375, 13.8542853196462, 13.7608026663462, 
    13.7187414169312, 13.6086111863454, 13.287735303243, 13.1619271437327, 
    12.7353624502818, 12.1838668982188, 11.8532002766927, 11.8354760805766, 
    11.7362672487895, 11.7333873907725, 11.5870920022329, 11.2722353935242, 
    11.0725568135579, 10.9285651048025, 11.0542931556702, 11.1458199818929, 
    11.0035116672516, 10.7099262078603, 10.6812395254771, 10.4409442742666, 
    10.2368634541829, 9.98233977953593, 9.76400502522787, 9.53174328804016, 
    9.26571981112162, 9.24029572804769, 9.33757742245992, 9.35421347618103, 
    17.569976594713, 17.2467642890082, 17.290078692966, 17.1035338507758, 
    16.788572523329, 16.3662221696642, 16.2446363237169, 16.2455399831136, 
    16.1274789174398, 16.2404865688748, 16.1693587832981, 16.0955412122938, 
    16.0071778827243, 15.9049780103895, 15.5378581153022, 15.2406288782756, 
    14.9144949383206, 14.8854532241821, 14.1397955152724, 13.6351191202799, 
    13.6026152504815, 14.0081446965535, 13.8747368918525, 13.7173813713921, 
    13.5757745107015, 13.1989316940308, 12.9187299940321, 12.3610553741455, 
    11.7746045854357, 11.4823514090644, 11.4825720257229, 11.4868247773912, 
    11.4990451600817, 11.7097430759006, 11.2997133466933, 11.2384759055244, 
    10.964741812812, 11.0447864532471, 11.0755052566528, 10.8023805618286, 
    10.8496902253893, 10.8572898440891, 10.2761414845785, 9.75024318695068, 
    9.85389433966743, 9.49061563279894, 9.12722259097629, 9.2241399553087, 
    9.19973776075575, 9.32647874620226, 9.29020108116998, 17.8756773206923, 
    17.6297878689236, 17.0689252217611, 16.7287686665853, 16.5870543585883, 
    16.4807275136312, 16.1611103481717, 16.198420630561, 16.1590167151557, 
    16.0821250279744, 16.0825830035739, 16.0507758458455, 15.9843485090468, 
    15.8028156492445, 15.608029683431, 15.3899722629123, 15.121560520596, 
    14.2839774290721, 13.3028551737467, 13.0803511937459, 13.1461062431335, 
    13.4151796499888, 13.5497903029124, 13.5905869801839, 13.4388221899668, 
    12.8800951639811, 12.587162733078, 12.1518103281657, 11.5915264288584, 
    11.3111531734467, 11.095096429189, 11.0714058081309, 11.0993487040202, 
    11.3157296975454, 11.2154105504354, 11.0974852244059, 10.8645830154419, 
    10.8171068032583, 10.8643432458242, 10.7589556376139, 10.4802484512329, 
    10.6074829101562, 10.0276446342468, 9.64030305544535, 9.38900009791056, 
    9.19114589691162, 9.26121393839518, 9.3174409866333, 9.32460363705953, 
    9.28718034426371, 9.28494834899902, 17.460947672526, 17.2921045091417, 
    16.9064945644803, 16.8219634162055, 16.7925391727024, 16.5447442796495, 
    16.2759034898546, 16.1724580128988, 15.9177476035224, 15.9008036719428, 
    15.866995493571, 15.8210973739624, 15.7004843817817, 15.5838333765666, 
    15.5269913143582, 15.1475962532891, 14.5017631318834, 13.5341317653656, 
    12.9784826437632, 12.9189412593842, 13.1180390516917, 13.3457023302714, 
    13.4151781400045, 13.4620412985484, 13.2540368239085, 12.5827696323395, 
    12.2628451188405, 11.7487033208211, 11.3881251811981, 11.2123995621999, 
    11.060887893041, 11.0526096820831, 10.7692728837331, 11.0099306106567, 
    10.8564976851145, 10.7845520178477, 10.6250243186951, 10.7084084351858, 
    10.7724155584971, 10.4239570299784, 10.3792924880981, 10.0790359179179, 
    9.70093472798665, 9.5265306631724, 9.55407087008158, 9.14119784037272, 
    9.26633985837301, 9.46097207069397, 9.31397517522176, 9.11934463183085, 
    9.28313080469767, 17.3682842254639, 17.2471894158257, 16.9193670484755, 
    16.8115914662679, 16.8810886806912, 16.6719301011827, 16.2131411234538, 
    16.1612383524577, 15.795837826199, 15.6934294170803, 15.6967204411825, 
    15.6943811840481, 15.3774884541829, 15.3446379767524, 15.3773932986789, 
    14.9805707931519, 13.7670423719618, 13.0132239659627, 12.9265489578247, 
    13.1503536436293, 13.295097457038, 13.2833137512207, 13.3486553827922, 
    13.4184143278334, 13.0149866739909, 12.3825714323256, 11.7942488988241, 
    11.2635938856337, 11.0550860299004, 11.1337244245741, 11.1229219436646, 
    11.0452704959446, 10.8799964057075, 10.6041901906331, 10.4979076385498, 
    10.3600741492377, 10.5765366024441, 10.5863953696357, 10.4602131313748, 
    10.6872665617201, 10.4889279471503, 10.1740267011854, 9.657593621148, 
    9.80379030439589, 9.77239269680447, 9.59166929456923, 9.33735423617893, 
    9.36344146728516, 9.21082602606879, 9.00909847683377, 9.38681104448107, 
    17.6048810746935, 17.2099829779731, 16.8422730763753, 16.8244101206462, 
    16.8669668833415, 16.6695868174235, 16.177431318495, 16.1357449425591, 
    15.6615494622125, 15.6309589809842, 15.5704087151421, 15.4403504265679, 
    15.3234673606025, 15.2438584433662, 15.1414667765299, 14.4632595909966, 
    13.1980572806464, 12.8490618069967, 13.0770213603973, 13.2958097457886, 
    13.3580228487651, 13.3060825665792, 13.2893598079681, 13.2881183624268, 
    12.780524969101, 12.1601657072703, 11.3866142431895, 11.1056428750356, 
    11.2059735457102, 11.1468830108643, 11.0570120811462, 11.059386809667, 
    10.9563518365224, 10.6054191589355, 10.3788825670878, 10.3714208602905, 
    10.5570543607076, 10.5125839710236, 10.4468135039012, 10.8159352938334, 
    10.6987140973409, 10.4728709856669, 9.88036672274272, 9.73555493354797, 
    9.77897310256958, 9.55955600738525, 9.44276229540507, 9.36133503913879, 
    9.26112524668376, 9.25328882535299, 9.84788568814596, 17.3467415703668, 
    17.0314617156982, 17.1708937750922, 17.0271538628472, 16.8579906887478, 
    16.3788168165419, 16.1856293148465, 16.1105258729723, 15.544707192315, 
    15.6890062756009, 15.185282919142, 14.6420967313978, 15.0363584094577, 
    15.0997334586249, 15.0147565205892, 14.0352684656779, 12.9967965020074, 
    12.7035621007284, 13.1184571584066, 13.318962097168, 13.3493412335714, 
    13.2460509141286, 13.293865998586, 13.2275763352712, 12.7051961421967, 
    11.8372422854106, 11.1144257386525, 11.0139896869659, 11.2271356582642, 
    11.2823483149211, 10.9825354417165, 10.9881097475688, 11.0766909917196, 
    10.6976267496745, 10.3821472326914, 10.285730044047, 10.5012300014496, 
    10.4193830490112, 10.5050875345866, 10.7123951117198, 10.7778221766154, 
    10.5599930286407, 10.0907887617747, 9.78257417678833, 9.8262669245402, 
    9.6224148273468, 9.54590805371602, 9.23143712679545, 9.25817863146464, 
    9.5073143641154, 10.0336559613546, 17.4319311777751, 17.2045957777235, 
    17.1266655392117, 17.1037693023682, 16.4507217407227, 16.2148696051704, 
    16.2770983378092, 16.2024088965522, 15.8356399536133, 15.6362585491604, 
    14.8103292253282, 14.3505212995741, 14.4962063895331, 15.0458743837145, 
    14.9758562511868, 13.791389465332, 12.9701467090183, 12.5238242679172, 
    12.920093536377, 13.2651773028904, 13.2902026706272, 13.2864519755046, 
    13.1227703094482, 13.1418646706475, 12.5879309972127, 11.6451784769694, 
    10.965217060513, 10.996886783176, 11.1746135287815, 11.2091870837741, 
    11.0596073998345, 11.1919777128432, 11.1708173751831, 10.732323328654, 
    10.383118947347, 10.2475580639309, 10.430459022522, 10.4234550264147, 
    10.5280135472616, 10.6547223197089, 10.4994524849786, 10.4587461683485, 
    10.2879297468397, 9.99062559339735, 9.73448912302653, 9.66484949323866, 
    9.67306031121148, 9.12308523390028, 8.60857031080458, 9.73774878184001, 
    9.93783940209283, 17.7426310645209, 17.2467839982775, 17.2558591630724, 
    17.0870255364312, 16.9140588972304, 16.6114891899957, 16.3309302859836, 
    16.2349757088555, 15.8012108272976, 15.3949406941732, 14.6569734149509, 
    14.4836086697049, 14.2996658749051, 14.3127856784397, 14.631756040785, 
    13.4556488460965, 13.0547329584757, 12.6089690526327, 12.5262390772502, 
    12.9076915582021, 13.1352797349294, 13.0529099305471, 12.9721416632334, 
    12.9142814477285, 12.631405433019, 11.639627456665, 11.005117336909, 
    10.9757498900096, 11.2637555599213, 11.290357430776, 11.1141438484192, 
    11.1396334966024, 11.0966595013936, 10.9864366849264, 10.6796259085337, 
    10.5795420805613, 10.4898873964945, 10.377782980601, 10.740374883016, 
    10.5609070460002, 10.4552805423737, 10.4709061781565, 10.2105224927266, 
    10.1404983997345, 9.89640402793884, 9.55968356132507, 9.61736567815145, 
    9.15096513430277, 9.5605727036794, 10.1349766254425, 9.917990843455, 
    17.3022912343343, 17.2915376027425, 17.3734007941352, 17.1806040869819, 
    17.290882534451, 17.0435678693983, 16.8217046525743, 16.2223552068075, 
    15.646653175354, 15.1500265333388, 14.4833731121487, 14.524974822998, 
    14.2387347751194, 14.0251733991835, 13.9268012576633, 13.2087199952867, 
    13.0942366917928, 12.6067266464233, 12.5793677171071, 12.5140307744344, 
    12.9733895460765, 12.9117290178935, 12.8015755812327, 12.7889177799225, 
    12.4964071114858, 11.8304862181346, 11.1511138280233, 11.2855168978373, 
    11.565601905187, 11.8879539966583, 11.2252229849497, 11.0755345026652, 
    10.9929705460866, 11.0652424494425, 11.0222911039988, 10.652756690979, 
    10.7282264232635, 10.6755494276683, 10.7168610095978, 10.51473681132, 
    10.512821038564, 10.501638174057, 10.0050985018412, 10.1516427199046, 
    9.78515823682149, 9.57314658164978, 9.57317193349203, 9.07371536890666, 
    10.0849494139353, 10.2379088401794, 9.95501446723938, 16.9740746815999, 
    16.8942970699734, 17.1102587381999, 17.2111373477512, 17.0644520653619, 
    16.9884149763319, 16.6795817481147, 16.1292503145006, 15.5100816090902, 
    14.8457256952922, 14.3423201243083, 14.6093082427979, 14.1656976275974, 
    14.2082139121162, 13.9503124025133, 13.2660470538669, 13.0683804617988, 
    12.7118395699395, 12.9518695407444, 12.7414744695028, 12.7286059061686, 
    12.7921856774224, 12.5535247590807, 12.5680008994208, 12.3134245342678, 
    12.077379544576, 11.7108671400282, 11.757499270969, 11.9454306496514, 
    12.0341949462891, 11.376263194614, 10.9505405426025, 11.1207387712267, 
    11.044123755561, 11.0109824074639, 10.6947761111789, 10.9235778384739, 
    10.8852110968696, 11.0443112055461, 10.9042001300388, 10.6588489744398, 
    10.6422628826565, 10.4492073059082, 10.1562774446276, 10.0087998708089, 
    9.61215782165527, 9.40678066677517, 9.37638007269965, 10.2657016118368, 
    10.141212993198, 9.82807985941569, 16.5641589694553, 16.7864089541965, 
    16.769844479031, 17.4961310492622, 17.0218609703912, 17.0287634531657, 
    16.4525731404622, 16.0954038831923, 15.723658879598, 14.8906761805216, 
    14.6168660057916, 14.6325047810872, 14.1287395689223, 14.1722588009304, 
    14.1593129899767, 13.505649778578, 13.077345000373, 12.7536098162333, 
    13.0262541770935, 12.9246857961019, 12.4908056259155, 12.3561503887177, 
    12.3698318799337, 12.5346681276957, 12.5720755259196, 12.3355650901794, 
    12.2937006950378, 11.7628772258759, 11.6831323305766, 11.6334730784098, 
    11.3377277056376, 10.9273862838745, 10.8067313035329, 10.7725114822388, 
    10.7135492960612, 10.6291739940643, 10.224999666214, 10.3875000476837, 
    10.359375, 10.4455355235509, 10.3803132375081, 10.5753334363302, 
    10.2445140566145, 9.7616774559021, 9.48951825228604, 9.23490405082703, 
    9.48468780517578, 10.0812103271484, 9.84556796334007, 9.52770177523295, 
    16.4022036658393, 16.3657383388943, 16.5491631825765, 16.7517846425374, 
    16.8795532650418, 16.6773317125108, 16.4428257412381, 15.9536216523912, 
    15.7590149773492, 15.0648759206136, 14.5261031256782, 14.5532442728678, 
    14.1375183529324, 14.1608899434408, 14.2248752382067, 13.5711562898424, 
    13.2958799997965, 12.9092145760854, 13.1161286036173, 13.1967673301697, 
    12.5328164100647, 12.253123998642, 12.1907619635264, 12.2594504356384, 
    12.7503277460734, 12.7308425108592, 12.3270847002665, 11.2912915547689, 
    11.4126833279928, 11.3542092641195, 11.0436531702677, 10.8888442516327, 
    10.8517874876658, 11.0424999757247, 10.7374998728434, 10.4382292429606, 
    10.1969999313354, 10.3062500953674, 10.197500038147, 10.1999998092651, 
    10.453125, 10.2929686307907, 9.16249990463257, 9.2854167620341, 
    9.59549989700317, 9.39770857493083, 9.78677225112915, 9.67499987284342, 
    9.70499992370605, 16.4472365909153, 16.324092441135, 16.5015936957465, 
    16.6630365583632, 16.5830006069607, 16.64574347602, 16.4932539198134, 
    16.2474066416423, 15.8686803181966, 15.1726971732246, 14.7735238605075, 
    14.5325618320041, 14.1010141372681, 14.2442448933919, 14.2043594784207, 
    13.7759033838908, 13.4057109620836, 13.2190894020928, 13.2015274895562, 
    13.2613598505656, 12.6793841256036, 12.3790841632419, 12.2591648101807, 
    12.3432820638021, 12.768692334493, 13.1034721798367, 11.9586341645983, 
    11.2172819773356, 11.5160697301229, 11.5247788959079, 11.334097120497, 
    10.2851851781209, 10.6541669368744, 10.3499999046326, 10.7302083969116, 
    11.0625, 10.3839288439069, 10.0362501144409, 11.0500001907349, 10.3125, 
    10.3862501144409, 9.75, 10.1999998092651, 9.54166666666667, 
    9.70666631062826, 9.76518938276503, 9.78986114925808, 10.2694665061103, 
    9.81944465637207, 9.82392480638292, 9.77708339691162, 16.3727325863308, 
    16.425689485338, 16.2975966135661, 16.4487592909071, 16.7254473368327, 
    16.3970553080241, 16.1210779613919, 16.212546772427, 16.112735218472, 
    15.3696445888943, 14.9236612319946, 14.3538378609551, 14.0494588216146, 
    14.263196627299, 14.4109831915961, 14.0616061952379, 13.5564122729831, 
    13.4027311007182, 13.4057706197103, 13.2890654404958, 12.7095372676849, 
    12.4876538912455, 12.2729818026225, 12.2731535434723, 12.4404068787893, 
    12.9239672025045, 11.819731314977, 11.1846250693003, 11.8114964167277, 
    11.560378854925, 11.2263888253106, 11.6118750572205, 11.8500003814697, 
    10.8900003433228, 10.4500001271566, 10.0406248569489, 10.1999998092651, 
    10.3078126907349, 10.2000002861023, 9.64204216003418, 9.58363395267063, 
    9.91185609499613, 9.77400024731954, 9.18947919209798, 9.72964421908061, 
    9.82457224527995, 9.37186543146769, 16.5706799825033, 16.604513168335, 
    16.4184457990858, 16.2329580518934, 16.1707442601522, 15.7429925070869, 
    16.0372923745049, 16.3541675143772, 16.4783642027113, 15.6719504462348, 
    15.2432831658257, 14.0683244069417, 13.909828291999, 14.0342269473606, 
    13.9330061806573, 13.8282095591227, 13.7222871780396, 13.6324714024862, 
    13.4452963670095, 13.3711846669515, 12.8486223220825, 12.4256115754445, 
    12.3681372801463, 12.5341523488363, 12.6078248818715, 12.5849274794261, 
    11.9713631470998, 11.4750076135, 11.6180965900421, 10.8225004196167, 
    11.6250001192093, 11.2763890160455, 8.625, 10.875, 9.8746874332428, 
    9.73693171414462, 9.60545444488525, 9.44629796346029, 8.29400690396627, 
    8.50310778617859, 8.63380159031261, 8.3155323266983, 16.6619249979655, 
    16.3247612847222, 16.3966727786594, 16.2913282182482, 16.2184419631958, 
    16.0607453452216, 15.978674782647, 16.1271110110813, 16.0291413201226, 
    15.7388139300876, 15.2097872628106, 14.1112162272135, 13.7374059889052, 
    13.6531474855211, 13.622554037306, 13.6083008448283, 13.725484000312, 
    13.6882996029324, 13.156261338128, 13.0467420154148, 12.7939172320896, 
    12.5313848919339, 12.3456312815348, 12.2808001836141, 12.0348637898763, 
    11.9450873268975, 11.7764410442776, 11.5850460264418, 8.24499979019165, 
    8.83703136444092, 8.65571673711141, 8.13243993123372, 16.5140448676215, 
    16.3230234781901, 16.3522012498644, 16.2969786326091, 16.2689734564887, 
    16.015230178833, 15.8514700995551, 15.931361940172, 15.805475446913, 
    15.2505209181044, 14.5980223549737, 14.1234780417548, 13.9184607399835, 
    13.7328272925483, 13.5142168468899, 13.2741550869412, 13.4903222190009, 
    13.6399835745494, 13.1961416403453, 12.9007976055145, 12.6945463816325, 
    12.8498746554057, 12.5563952128092, 12.2713366349538, 11.8334614146839, 
    16.5331645541721, 16.364187028673, 16.2841521369086, 16.1686462826199, 
    15.92754067315, 15.7410028245714, 15.4230078591241, 14.9539959165785, 
    14.5129081938002, 14.2449222140842, 14.1970852745904, 14.1741861767239, 
    14.1869130664402, 14.0097263124254, 13.5460466808743, 13.2326777776082, 
    13.2805486255222, 13.5336263179779, 13.2016479174296, 12.766566435496, 
    12.8220920562744, 12.5599935849508, 12.4218448003133, 12.07634973526, 
    16.6038597954644, 16.5156673855252, 16.3608623080783, 16.0791866514418, 
    15.8101507822673, 15.499446551005, 14.5192971759372, 14.2581359015571, 
    14.2023625903659, 14.0265281465318, 14.2044197718302, 14.1248016357422, 
    14.1972006691827, 14.1889118618435, 13.6775290171305, 13.2093381881714, 
    13.2615043852064, 13.3953879674276, 13.1230317221748, 13.1849196751912, 
    13.0083642535739, 12.4394025802612, 16.6424590216743, 16.4437077840169, 
    16.5516276889377, 16.087976137797, 15.7279567718506, 15.2799331876967, 
    14.1046301523844, 14.0488941404555, 14.1358157263862, 13.9478526645237, 
    14.1516244676378, 14.0654578738742, 14.2287861506144, 14.1602827707926, 
    13.6579386393229, 13.20754898919, 13.2424987157186, 13.459893544515, 
    13.5103556315104, 12.9808926582336, 12.6556489467621, 11.7840672492981, 
    16.4998965793186, 16.6501901414659, 16.5171930525038, 16.1847087012397, 
    15.5334700478448, 14.8879103130764, 13.9995861053467, 14.1505849626329, 
    14.1780576705933, 13.9164016511705, 14.0218182669746, 13.956203672621, 
    14.0840938356188, 13.7737268871731, 13.4711937374539, 13.1570962270101, 
    13.3236507839627, 13.3783466815948, 13.2886896928151, 12.7979076558893, 
    16.3950642479791, 16.7268986172146, 16.6561029222276, 16.4220485687256, 
    15.7097977532281, 14.9390098783705, 14.1184793048435, 14.2552797529433, 
    14.231750064426, 14.0930458704631, 14.0609507030911, 13.8806876076592, 
    14.0591660605537, 13.5774208704631, 13.4326086044312, 13.5325814353095, 
    13.4106767442491, 13.0715370178223, 12.7530767917633, 16.439006169637, 
    16.7028528849284, 16.7325738271077, 16.6549725002713, 16.1856139500936, 
    15.4497060775757, 14.7032270431519, 14.5607945124308, 14.4572270711263, 
    14.1499063703749, 13.9991596009996, 13.8610765669081, 13.8843505647447, 
    13.9023983213637, 13.735852877299, 13.6126681433784, 13.2512315511703, 
    16.0899913575914, 16.0525305006239, 16.2904851701525, 16.6302602556017, 
    16.6716819339328, 16.3437392976549, 15.6239958869086, 15.2742275661892, 
    14.5786729388767, 14.3867282867432, 13.9765875074599, 13.6398431989882, 
    13.478899108039, 13.5777011447483, 13.5028555128309, 13.3067380905151, 
    16.2068144480387, 15.9232803980509, 16.0462001164754, 16.53820376926, 
    16.6030871073405, 16.5839795006646, 16.1331043243408, 15.5778775744968, 
    14.7687424553765, 14.6740702523126, 14.1620410283407, 13.3845592074924, 
    13.2746832105849, 13.3051026662191, 13.1336999469333, 16.3684741126166, 
    16.0874963336521, 15.7142188813951, 16.3143032921685, 16.5479772355821, 
    16.5178209940592, 16.2935203976101, 15.8225991990831, 15.2659853829278, 
    14.4704221089681, 13.8783077663845, 13.5206939909193, 13.0379188855489, 
    12.8501987457275, 16.394600338406, 16.2023684183757, 15.7180952495999, 
    15.9947347640991, 16.3293688032362, 16.1478969785902, 15.8493882285224, 
    15.4642003377279, 15.0793790817261, 14.161416053772, 13.4991675615311, 
    13.563195016649, 16.4593230353461, 16.1983723110623, 15.750404993693, 
    15.5719236797757, 15.5858874850803, 15.3222267362807, 14.9526377783881, 
    14.7208382288615, 14.6554622650146, 13.9821109771729, 13.6062479019165, 
    13.6595776875814, 16.4533333248562, 16.2513015535143, 15.9043964809842, 
    15.5947280459934, 15.2626521852281, 15.0579289330377, 14.8063691457113, 
    14.3365809122721, 14.2872684266832, 13.7550080617269, 13.8551460901896, 
    13.5207580990261, 16.3158927493625, 16.2043800354004, 15.8539445665148, 
    15.6470822228326, 15.5958701239692, 15.606875843472, 14.6812529034085, 
    14.3407680723402, 14.0926985210843, 13.9365146425035, 14.0482921600342, 
    16.2094508277045, 15.8767967224121, 15.7680886586507, 15.727460331387, 
    15.7971051534017, 15.7167098787096, 14.4850766923692, 14.4568254682753, 
    14.2645647260878, 14.184963438246, 14.2129074732463, 15.9832297431098, 
    15.6064812342326, 15.7826724582248, 15.8883006837633, 15.778157764011, 
    15.5188763936361, 14.8337375852797, 14.752785258823, 14.589465353224, 
    14.5044542948405, 14.3177603085836, 15.764713605245, 15.584216647678, 
    15.4937999513414, 15.737473487854, 15.1769664552477, 15.1558961868286, 
    15.0613864262899, 14.9855097664727, 14.9620975255966, 14.6877051989237, 
    15.4131152894762, 15.5294861263699, 15.2924204932319, 15.3540030585395, 
    15.1913794411553, 15.2409071392483, 15.1095952987671, 15.0799673928155, 
    15.1124964820014, 15.7624419530233, 15.7824169794718, 15.4803779390123, 
    15.1959829330444, 15.2595366372002, 15.259891404046, 15.1860720316569, 
    15.1839969423082, 14.9985092878342, 16.298166486952, 16.1154217190213, 
    16.2535994847616, 15.7027917438083, 15.4867106543647, 15.0263305240207, 
    15.0185871124268, 14.8061496734619, 16.5446578131782, 16.3696399264865, 
    16.5107989841037, 15.477232615153, 14.9267551634047, 16.1303270128038, 
    15.6558390723334, 15.7767386966281, 14.8098753293355, 11.2923981802804, 
    11.2992696762085, 11.2982950210571, 11.2970762252808, 11.2958545684814, 
    11.294629573822, 11.2391742070516, 10.14399822553, 8.83433310190837, 
    7.81750647226969, 9.48060637253981, 8.3945129101093, 7.37896112295297, 
    9.05040022043081, 7.81111368766198, 6.78067544790415, 9.78600271542867, 
    8.49324591954549, 7.2356166044871, 6.28707544008891, 11.3992643356323, 
    11.3982839584351, 11.397057056427, 11.395827293396, 11.3945941925049, 
    11.0060035387675, 11.4494684764317, 14.2498426437378, 14.1591596603394, 
    13.9784469604492, 12.437292098999, 12.0860271453857, 11.6548728942871, 
    11.4536552429199, 33.2130012512207, 33.2099990844727, 33.2060012817383, 
    33.1650009155273, 33.2050018310547, 33.2439994812012, 33.3199996948242, 
    14.5496816635132, 14.5485038757324, 14.547080039978, 14.5456113815308, 
    13.9343614578247, 12.113597869873, 11.5768885612488, 10.8239393234253, 
    10.4896655082703, 33.2140007019043, 33.2169990539551, 33.2190017700195, 
    33.2140007019043, 33.1669998168945, 33.185001373291, 33.2880001068115, 
    33.5415000915527, 33.751501083374, 17.4407428105672, 17.5064427057902, 
    17.764352162679, 17.2335424423218, 16.8680308659871, 16.827561378479, 
    16.5930344263713, 16.4485470453898, 16.3762029012044, 16.3291994730632, 
    16.2919165293376, 16.2883930206299, 15.9193553924561, 15.5074424743652, 
    15.2779763539632, 14.8105263710022, 14.2899905840556, 14.2428450584412, 
    13.9191869099935, 13.5803155899048, 13.2652708689372, 13.2064512570699, 
    13.1351172129313, 13.1786985397339, 13.2495759328206, 13.3462985356649, 
    13.3576793670654, 12.9369489351908, 12.384074529012, 11.8705547650655, 
    11.7326839764913, 11.8096005121867, 11.6234501202901, 11.2959068616231, 
    10.8587563832601, 10.7948732376099, 10.5698078473409, 10.6259299914042, 
    10.7241797447205, 10.8368198076884, 10.4992993672689, 10.4059850374858, 
    10.6148476600647, 10.4257300694784, 10.3511358896891, 10.4992863337199, 
    10.1503248214722, 9.89671421051025, 9.70059219996134, 9.35493564605713, 
    9.22393369674683, 17.5388819376628, 17.3847348954942, 17.5870585971408, 
    17.4175179799398, 16.9635384877523, 16.7779210408529, 16.5465571085612, 
    16.4346084594727, 16.3184941609701, 16.3516354031033, 16.2787736256917, 
    16.2906379699707, 16.0462183422512, 15.6532618204753, 15.4636304643419, 
    14.9801843431261, 14.3810562557644, 14.4178789456685, 14.0910464127858, 
    13.8216909567515, 13.5610047181447, 13.4476498762767, 13.3211879730225, 
    13.361141761144, 13.4090408484141, 13.3806128501892, 13.3229986826579, 
    12.8492257595062, 12.1944622993469, 11.9729450543722, 11.7037199338277, 
    11.6540182431539, 11.3939089775085, 11.3173433144887, 10.9852752685547, 
    10.7588144938151, 10.6383197307587, 10.8193749586741, 11.0014649232229, 
    10.9779201348623, 10.7009816964467, 10.5188834667206, 10.53559923172, 
    10.4537117481232, 10.4813772837321, 10.3381107648214, 9.92720603942871, 
    9.91082525253296, 9.4888121287028, 9.82123525937398, 9.43304228782654, 
    17.2280868954129, 17.0269304911296, 17.2656375037299, 17.2895035213894, 
    16.9593048095703, 16.5276118384467, 16.3826402028402, 16.3707754347059, 
    16.2427618238661, 16.2650176154243, 16.2123875088162, 16.1479350195991, 
    15.9141688876682, 15.7642867830065, 15.5199688805474, 15.134042845832, 
    14.7055932150947, 14.6951745351156, 14.4936854044596, 14.2109311421712, 
    13.9432559013367, 13.8570148150126, 13.7737342516581, 13.6777450243632, 
    13.5949985186259, 13.31573955218, 13.1705929438273, 12.7601448694865, 
    12.0645410219828, 11.772305727005, 11.8752253055573, 11.6757500171661, 
    11.6573831240336, 11.4326567649841, 11.1641902923584, 10.9662425518036, 
    10.8254458109538, 10.9798767566681, 11.1079564889272, 10.98406513532, 
    10.6595888137817, 10.6160031159719, 10.5024708112081, 10.3648361365, 
    10.2591973145803, 10.0444253285726, 9.70507113138835, 9.57716075579325, 
    9.78680316607157, 9.72938895225525, 9.77437766393026, 17.2973376380073, 
    17.1524969736735, 17.2719898223877, 17.0888646443685, 16.7700231340196, 
    16.3436459435357, 16.231930202908, 16.1967368655735, 16.0700204637316, 
    16.2520463731554, 16.1152317259047, 16.0562629699707, 16.0002245373196, 
    15.8805467817518, 15.5060858196682, 15.2457278569539, 14.9094950358073, 
    14.8931783040365, 14.1325806511773, 13.6351594924927, 13.5974298053318, 
    13.9370345009698, 13.9151313569811, 13.7510693868001, 13.5764740837945, 
    13.2057483461168, 12.9598259396023, 12.4068162706163, 11.7518193986681, 
    11.4442266888089, 11.4316877788968, 11.4834878709581, 11.523166762458, 
    11.6120381885105, 11.2007990943061, 11.1372691260444, 10.9677833980984, 
    11.0022110409207, 11.1484022140503, 10.893433464898, 10.7816914452447, 
    10.6569577323066, 10.3810400433011, 10.0717275407579, 9.89221668243408, 
    9.69908693101671, 9.28733942243788, 9.38884109920926, 9.55215930938721, 
    9.75488313039144, 9.34801959991455, 17.7018775939941, 17.4660538567437, 
    17.0549979739719, 16.7113265991211, 16.5339397854275, 16.4405858781603, 
    16.1599079767863, 16.1559916602241, 16.0877589119805, 16.0775277879503, 
    16.0705021752252, 16.0257070329454, 15.9832550684611, 15.8134645885891, 
    15.6235647201538, 15.3505655924479, 15.1098574532403, 14.2944447199504, 
    13.2946399052938, 13.0783290068309, 13.149749994278, 13.388511578242, 
    13.5594705740611, 13.6090795993805, 13.4336241881053, 12.8791151841482, 
    12.6679384708405, 12.1780090332031, 11.5887352625529, 11.3268880049388, 
    11.0781365235647, 11.0822907288869, 11.1047673225403, 11.375014146169, 
    11.216010093689, 11.0769859949748, 10.8608965873718, 10.8306731383006, 
    10.9714101155599, 10.8616866270701, 10.5439930756887, 10.5260449250539, 
    10.1821023623149, 9.71200331052144, 9.47475401560465, 9.3314962387085, 
    9.24781084060669, 9.48219537734985, 9.5135924021403, 9.69603045781454, 
    9.38164075215658, 17.2075252532959, 16.9164377848307, 16.7531000773112, 
    16.5877537197537, 16.7883904774984, 16.5199752383762, 16.2837166256375, 
    16.1371264987522, 15.8683258692423, 15.8821942011515, 15.853571150038, 
    15.8107686572605, 15.7012091742622, 15.6009178161621, 15.5611710018582, 
    15.1619083616469, 14.4493289523655, 13.5348171393077, 12.9620436827342, 
    12.9337914784749, 13.1298352877299, 13.3412856260935, 13.4175929228465, 
    13.4418710072835, 13.1746949354808, 12.5877104600271, 12.3172214031219, 
    11.8356481393178, 11.4718464215597, 11.2276880741119, 11.049028635025, 
    11.045089006424, 10.777866601944, 11.0523693561554, 10.8674148718516, 
    10.7759142716726, 10.638058423996, 10.6974539756775, 10.7858820756276, 
    10.5803984006246, 10.3985203107198, 10.176100174586, 9.82352526982625, 
    9.50128157933553, 9.58844033877055, 9.41781783103943, 9.30671898523966, 
    9.43633111317953, 9.37206546465556, 9.26343854268392, 9.26848371823629, 
    17.1495793660482, 17.160275777181, 16.6843255360921, 16.7523517608643, 
    16.8459964328342, 16.7128092447917, 16.2409269544813, 16.1007401148478, 
    15.760520723131, 15.6748655107286, 15.7049721611871, 15.6856836742825, 
    15.3641019397312, 15.3640046649509, 15.3919418123033, 14.9956979751587, 
    13.8114958869086, 13.0324186748928, 12.9487299389309, 13.1909761428833, 
    13.307394557529, 13.2388354407416, 13.3503861957126, 13.4363278283013, 
    12.8917186525133, 12.3260537253486, 11.8344400193956, 11.3805688222249, 
    11.1254505581326, 11.2302769554986, 11.1426777309842, 11.0945937898424, 
    10.8149979909261, 10.605357170105, 10.4693428675334, 10.3603999879625, 
    10.6697557237413, 10.6357243855794, 10.6634780036079, 10.5452874501546, 
    10.412646399604, 10.0837711758084, 9.7818816502889, 9.75718678368462, 
    9.78448602888319, 9.74895371331109, 9.32527054680718, 9.30478074815538, 
    9.29707770877414, 8.99779510498047, 9.13979456159804, 17.4451722039117, 
    17.2140373653836, 16.7872655656603, 16.7631732092963, 16.7930043538411, 
    16.6958406236437, 16.1672666337755, 16.1281063291762, 15.6475074556139, 
    15.6268667644925, 15.5411672592163, 15.3998907936944, 15.2880375120375, 
    15.2221475177341, 15.1643510394626, 14.420831574334, 13.2205651601156, 
    12.8584336439768, 13.0872968037923, 13.3223929405212, 13.3420946598053, 
    13.2794845104218, 13.3202245235443, 13.393151919047, 12.6596268018087, 
    12.1054422855377, 11.4106761614482, 11.1398917039235, 11.2859503428141, 
    11.1817394892375, 11.0647996266683, 11.0475951830546, 10.9447310765584, 
    10.5362267494202, 10.3696255683899, 10.404568751653, 10.4971151351929, 
    10.5301187038422, 10.5467182000478, 10.7386531829834, 10.6735095977783, 
    10.2884788513184, 9.90359576543172, 9.87823494275411, 9.85761181513468, 
    9.80824685096741, 9.50787790616353, 9.24784366289775, 9.21554613113403, 
    9.22816379865011, 9.68614284197489, 17.2389657762316, 17.332245932685, 
    17.255656560262, 16.7640213436551, 16.6935878329807, 16.249267578125, 
    16.1523412068685, 16.1110719045003, 15.5311112933689, 15.6546027925279, 
    15.165211253696, 14.6333677503798, 15.0711234410604, 15.144739151001, 
    15.1143581602308, 14.0374298095703, 13.0008378558689, 12.7053413391113, 
    13.142558892568, 13.3481151262919, 13.3473348617554, 13.2762741247813, 
    13.3252313931783, 13.280979235967, 12.5711283683777, 11.8401406606038, 
    11.1244633992513, 10.9418803056081, 11.1679409344991, 11.2313680648804, 
    10.8518197536469, 10.9485379060109, 11.0215732256571, 10.6116544405619, 
    10.3708675702413, 10.2186657587687, 10.2908293406169, 10.4383146762848, 
    10.5260616143545, 10.8519035975138, 10.7561483383179, 10.4498000144958, 
    10.1359905401866, 10.1063567002614, 10.1439924240112, 9.93781924247742, 
    9.61387777328491, 9.01830410957336, 9.17745772997538, 9.38219960530599, 
    9.75135882695516, 17.3454564412435, 17.3196603986952, 17.2995476192898, 
    16.920093536377, 16.2710818184747, 16.1630704667833, 16.2776605818007, 
    16.2184268103706, 15.7960197660658, 15.4518435796102, 14.8270867665609, 
    14.3459048800998, 14.5228421952989, 15.0626765357123, 15.0173397064209, 
    13.8168202506171, 12.9780972798665, 12.5278317133586, 12.8998722500271, 
    13.2642650604248, 13.2913848029243, 13.2883005142212, 13.1246996985541, 
    13.2212892108493, 12.6469249725342, 11.6443809933133, 10.9356098175049, 
    10.8593222300212, 10.9832741419474, 11.1199855804443, 10.8565094206068, 
    11.0441283120049, 11.1678572760688, 10.6329860687256, 10.4844217300415, 
    10.2186432944404, 10.3461641735501, 10.5795370737712, 10.6958471934001, 
    10.8045403162638, 10.5442174275716, 10.2853151957194, 10.202297422621, 
    10.216908454895, 9.97555213504367, 9.84572675493028, 9.47333611382378, 
    9.00349892510308, 8.55416059494019, 9.40628221299913, 9.61893325381809, 
    17.3993856641981, 17.3096018897163, 17.1915726131863, 17.1112217373318, 
    16.7407631344265, 16.5061451594035, 16.20858446757, 16.2470009062025, 
    15.8547709782918, 15.295890490214, 14.6251624425252, 14.4858654869927, 
    14.3394242392646, 14.3275000254313, 14.6703714794583, 13.4823314878676, 
    13.0550354851617, 12.6083656946818, 12.5174624125163, 12.9023237228394, 
    13.1393434206645, 13.0521223545074, 13.0329984823863, 12.9624485174815, 
    12.6550550460815, 11.6068156560262, 10.9220371246338, 10.9105775356293, 
    11.112429857254, 11.2496868769328, 11.0048973560333, 11.1257005532583, 
    11.0968091487885, 11.1034553845723, 10.8463124434153, 10.6015605926514, 
    10.3745791912079, 10.3327125708262, 10.724063316981, 10.5063453515371, 
    10.3605902194977, 10.216811577479, 10.2523464361827, 10.1469423770905, 
    9.83370288213094, 9.70165681838989, 9.54609886805216, 8.98902837435404, 
    9.36967412630717, 9.76374459266663, 9.75933615366618, 17.3326816558838, 
    17.1926663716634, 17.2495405409071, 17.1791195339627, 17.1378752390544, 
    16.7347558339437, 16.8453004625108, 16.2091883553399, 15.429412206014, 
    15.2000592549642, 14.4381632275052, 14.5834415223863, 14.2839691374037, 
    14.0598793029785, 13.9551079008314, 13.2249391343859, 13.1161798901028, 
    12.6196520328522, 12.6025187969208, 12.4885989824931, 13.0020501613617, 
    12.9303077061971, 12.8759775161743, 12.8731809457143, 12.5235437552134, 
    11.8249980608622, 11.0693385601044, 11.0548654397329, 11.2647552490234, 
    11.6467224756877, 11.24707086881, 11.1310584545135, 10.982291618983, 
    11.1407237052917, 11.1377499898275, 10.6342956225077, 10.645429054896, 
    10.5664873917898, 10.5935509204865, 10.3854250907898, 10.429660876592, 
    10.1516771316528, 10.0595843791962, 9.98465387026469, 9.75417447090149, 
    9.62610459327698, 9.50410087903341, 8.85821111996969, 9.95434641838074, 
    10.0515115261078, 9.7966882387797, 16.9656567043728, 16.831217235989, 
    16.9842688242594, 17.1450551350911, 17.0702472262912, 16.7899434831407, 
    16.6386144426134, 16.1530777613322, 15.299816555447, 14.9069203270806, 
    14.342488500807, 14.6631540722317, 14.2362846798367, 14.2684552934435, 
    14.0251836776733, 13.2357094022963, 13.054008907742, 12.7317117055257, 
    12.9805680380927, 12.7424490186903, 12.7436338000827, 12.8523179160224, 
    12.6534523434109, 12.6879812876383, 12.3202108807034, 11.9466883341471, 
    11.6239674886068, 11.3508372836643, 11.4637777540419, 11.66117699941, 
    11.3213027318319, 10.9387145572239, 11.0763154559665, 11.1426271862454, 
    10.9717258877224, 10.6548399395413, 10.7726944817437, 10.7227221594916, 
    10.7728110419379, 10.6327815585666, 10.5591249465942, 10.6058443917169, 
    10.0873055987888, 10.0147630903456, 9.80386585659451, 9.53582106696235, 
    9.47573068406847, 9.36817889743381, 9.93648264143202, 9.94683922661675, 
    9.72611151801215, 16.5090866088867, 16.6492144266764, 16.5952010684543, 
    17.0870407952203, 17.0446253882514, 16.9105008443197, 16.5867349836561, 
    16.0734278361003, 15.5878033108181, 14.935258547465, 14.5920299953885, 
    14.7352751625909, 14.19295946757, 14.2609718110826, 14.2289105521308, 
    13.4687583711412, 13.072898334927, 12.7608649730682, 13.0300293763479, 
    12.9030222098033, 12.5059202512105, 12.3714435100555, 12.3716680208842, 
    12.5713256994883, 12.5846848487854, 12.2934060891469, 12.2442331314087, 
    11.5323920683427, 11.5366507371267, 11.2615408463912, 10.8983155091604, 
    10.9227740547874, 10.792551279068, 10.7312454743819, 10.650000163487, 
    10.5281248092651, 10.4249992370605, 10.6836331685384, 10.1145162582397, 
    9.95956659317017, 9.50840441385905, 9.49896543676203, 9.39450287818909, 
    9.59418145815531, 9.91887863477071, 9.61937618255615, 9.44110608100891, 
    16.4035523732503, 16.3142681121826, 16.5729031032986, 16.7710522545709, 
    16.8290365007189, 16.6737128363715, 16.3198290930854, 16.1466997994317, 
    15.6035884221395, 14.8371493021647, 14.4870315127903, 14.5612229241265, 
    14.179835319519, 14.2306594848633, 14.2765067418416, 13.602996190389, 
    13.3350132836236, 12.8932615915934, 13.0981513659159, 13.1980506579081, 
    12.5831123193105, 12.2895526091258, 12.2410128911336, 12.3164131641388, 
    12.7605063120524, 12.7312200069427, 12.7159857749939, 11.3623367656361, 
    11.4062498410543, 11.1837647755941, 10.8795456452803, 10.9799999237061, 
    11.0142856325422, 10.5843750238419, 10.2750002543132, 10.5166666242811, 
    10.3874998092651, 10.03125, 9.65416669845581, 8.96875023841858, 
    9.49319038391113, 9.40146327018738, 9.73913892110189, 9.74921894073486, 
    9.62161461512248, 9.37903650601705, 16.3795827229818, 16.2851816813151, 
    16.5504048665365, 16.6814301808675, 16.5837773217095, 16.3863308164809, 
    16.2746351030138, 16.1323926713732, 15.8835319942898, 15.1011437310113, 
    14.7245102988349, 14.5585074954563, 14.126759952969, 14.3155279159546, 
    14.238107363383, 13.7243324915568, 13.3479553858439, 13.1800669564141, 
    13.1059674157037, 13.2116081449721, 12.6628757052951, 12.4210115008884, 
    12.4139116075304, 12.400127198961, 12.8697915607029, 13.4221063190036, 
    12.3515621423721, 11.2529466152191, 11.6287038591173, 11.5458333151681, 
    10.7699998855591, 10.5, 10.5, 9.63333320617676, 9.37395842870077, 
    9.76518938276503, 9.78986114925808, 10.2694665061103, 9.90138891008165, 
    9.76132678985596, 9.47968745231628, 16.3703763749864, 16.4563965267605, 
    16.3210928175184, 16.4553356170654, 16.6786566840278, 16.3975166744656, 
    16.1324668460422, 16.14061027103, 16.1756214565701, 15.3383597267999, 
    14.9030765957303, 14.3666244082981, 14.0920908186171, 14.329021135966, 
    14.43235206604, 14.0709100299411, 13.505552927653, 13.378001610438, 
    13.3943320115407, 13.2420449256897, 12.7390654881795, 12.5082244873047, 
    12.3541289965312, 12.3027341365814, 12.6718462308248, 13.0088854630788, 
    11.9913904666901, 11.1067533493042, 11.7124998786233, 11.3156249523163, 
    11.7225001335144, 11.8500003814697, 10.1999998092651, 9.62381303310394, 
    9.61759195327759, 9.91185609499613, 9.77400024731954, 9.18947919209798, 
    9.72964421908061, 9.80972862243652, 9.35545913378398, 16.5448188781738, 
    16.5985190073649, 16.4025565253364, 16.2700097825792, 16.2002195782132, 
    15.7051146825155, 16.0710322062174, 16.1290545993381, 16.5095568762885, 
    15.7875632180108, 15.2732830047607, 14.0392749574449, 13.9646011988322, 
    14.0643662346734, 13.9311156802707, 13.703929371304, 13.6686912112766, 
    13.6177020867666, 13.392098903656, 13.3191967010498, 12.8195343812307, 
    12.4510075251261, 12.4402766227722, 12.5910322666168, 12.664484500885, 
    12.7201476891836, 12.1219833691915, 11.2848091920217, 11.44553565979, 
    11.3250001907349, 11.9250001907349, 11.8500003814697, 9.8746874332428, 
    9.73693171414462, 9.60545444488525, 9.44629796346029, 8.29400690396627, 
    8.50310778617859, 8.63380159031261, 8.3155323266983, 16.6686242421468, 
    16.2902003394233, 16.3084083133274, 16.3120678795709, 16.3031611972385, 
    16.0414367251926, 16.0379333496094, 16.1350136862861, 16.0906114578247, 
    15.7648499806722, 15.3466540442573, 14.1293622122871, 13.7447201410929, 
    13.7007037268745, 13.6676157845391, 13.6110110812717, 13.7058689329359, 
    13.7111066182454, 13.178112771776, 13.1209448708428, 13.0040133794149, 
    12.666385544671, 12.4482323328654, 12.3404637442695, 12.1623722712199, 
    11.9744389851888, 11.8500232696533, 11.2524299621582, 8.24499979019165, 
    8.83703136444092, 8.65571673711141, 8.13243993123372, 16.5403406355116, 
    16.2991564008925, 16.3235251108805, 16.2656892140706, 16.2426399654812, 
    15.9517093234592, 15.8531581030952, 15.9068330128988, 15.7737753126356, 
    15.285098499722, 14.560937139723, 14.0976078245375, 13.8938873079088, 
    13.746277279324, 13.5482607947456, 13.3171566857232, 13.4715812471178, 
    13.6405780315399, 13.2797427972158, 13.0696603457133, 12.8959363301595, 
    12.9297362963359, 12.6171340942383, 12.3343273003896, 11.930721282959, 
    16.5466471778022, 16.3573864830865, 16.2689880794949, 16.1528973049588, 
    15.8969090779622, 15.7134613460965, 15.3852313359578, 14.9673113293118, 
    14.5700451533, 14.1746077007718, 14.0748168097602, 14.1612963146634, 
    14.1691550148858, 14.0053785112169, 13.5664491653442, 13.273754119873, 
    13.341518719991, 13.5921570460002, 13.3301290671031, 12.8692685763041, 
    12.974893172582, 12.5955250263214, 12.3460294405619, 11.9625511964162, 
    16.5912823147244, 16.4888617197673, 16.3214685651991, 16.0676229265001, 
    15.811291164822, 15.4803152084351, 14.4917457368639, 14.2731217278375, 
    14.2016354666816, 13.9625874625312, 14.123663160536, 14.1206193500095, 
    14.1267320844862, 13.9399176703559, 13.6106033325195, 13.2470088534885, 
    13.2922394010756, 13.4491234885322, 13.2477052476671, 13.2772703170776, 
    12.8879157172309, 12.101151254442, 16.5681726667616, 16.4052965376112, 
    16.3595566219754, 16.0470709270901, 15.7064392301771, 15.2620561387804, 
    14.0825543933445, 14.0308244493273, 14.1257830725776, 13.9278650283813, 
    14.1307524575127, 14.0774013731215, 14.1947414610121, 13.967144648234, 
    13.5602890650431, 13.082618077596, 13.1582802666558, 13.5898067951202, 
    13.608067035675, 13.0262001355489, 12.7287352879842, 11.4739905463325, 
    16.4649800194634, 16.5980508592394, 16.3801023695204, 16.0660315619575, 
    15.5540285110474, 14.9219880633884, 13.9893618689643, 14.1293178134494, 
    14.1629536946615, 13.9036535686917, 13.9691696166992, 13.9478034973145, 
    13.9750117195977, 13.7919626235962, 13.5572706858317, 13.3497524261475, 
    13.4293732113308, 13.4464832146962, 13.4504771232605, 12.8857918652621, 
    16.3486164940728, 16.6404033237033, 16.4792291853163, 16.2229801813761, 
    15.5113397174411, 14.9442427953084, 14.0887400309245, 14.2185688018799, 
    14.1997281180488, 14.0008041593764, 13.9454485575358, 13.7786398993598, 
    13.8965869479709, 13.5396828121609, 13.4341702991062, 13.6906346215142, 
    13.4519143634372, 13.1300687789917, 12.8366248607635, 16.3872392442491, 
    16.5062005784776, 16.5732460021973, 16.4525623321533, 16.0209333631727, 
    15.3451657825046, 14.5566850238376, 14.3687194188436, 14.2715724309285, 
    14.0126350190904, 13.8952207565308, 13.7502189212375, 13.7664789623684, 
    13.8529929055108, 13.7643551296658, 13.7043863932292, 13.2737722396851, 
    15.9179693857829, 15.9174177381727, 16.184186829461, 16.5807469685872, 
    16.5858296288384, 16.1775312423706, 15.3630091349284, 15.0879450903998, 
    14.529887093438, 14.2942399978638, 14.0433411068386, 13.6355029212104, 
    13.3580771552192, 13.4330078760783, 13.3101497226291, 13.2927070617676, 
    16.1044073104858, 15.8153400421143, 15.8336805767483, 16.4906862046983, 
    16.5301130082872, 16.475759294298, 15.9965153800117, 15.3403729332818, 
    14.7022546132406, 14.6283237669203, 14.183831108941, 13.3352387746175, 
    13.0657759772407, 13.0975022845798, 12.9501637352837, 16.1508238050673, 
    15.9797801971436, 15.533943494161, 16.2363501654731, 16.4382199181451, 
    16.3980880313449, 16.1896562576294, 15.6999911202325, 15.2381004757351, 
    14.4418787426419, 13.8279796176487, 13.4138003455268, 12.935110727946, 
    12.7844624519348, 16.2123974694146, 16.0621469285753, 15.6485826704237, 
    15.908673286438, 16.136890411377, 15.9293148252699, 15.6358903249105, 
    15.5702592002021, 15.0375299453735, 14.1145265367296, 13.4959172010422, 
    13.5376958847046, 16.2105462816026, 16.020029703776, 15.7237539291382, 
    15.3971811930339, 15.4040927886963, 14.8364209069146, 14.515329890781, 
    14.5084833568997, 14.4978573057387, 13.7617637846205, 13.4182469844818, 
    13.5606429841783, 16.2186965942383, 16.1408280266656, 15.8971775902642, 
    15.4921375910441, 15.0573002497355, 14.8071065478855, 14.4910953309801, 
    14.012776904636, 13.9995483822293, 13.4567006429036, 13.6281622250875, 
    13.5268115997314, 16.2446433173286, 16.0896283255683, 15.8415665096707, 
    15.4797661039564, 15.3096743689643, 15.2935651143392, 14.5714815987481, 
    14.0180371602376, 13.8443880081177, 13.6807550854153, 13.9667943318685, 
    16.1735319561428, 15.7790868547228, 15.7452500661214, 15.5913184483846, 
    15.4693118201362, 15.4816409216987, 14.4053270551893, 14.3087112638685, 
    14.1790743933784, 14.1159703996446, 14.2450405756632, 15.9771455128988, 
    15.5414890713162, 15.6925684611003, 15.7076189253065, 15.5450375874837, 
    15.428720580207, 14.8341129091051, 14.6506801181369, 14.5217547946506, 
    14.5445288552178, 14.3421430587769, 15.5865556928847, 15.6450942357381, 
    15.5338409211901, 15.6636292139689, 15.2317417992486, 15.1451901329888, 
    15.0424250496758, 15.1217485004001, 14.9169813394547, 14.5601162910461, 
    15.4519237942166, 15.7415877448188, 15.6251748402913, 15.3610517713759, 
    15.3192720413208, 15.3796740637885, 15.2405783335368, 15.1997252570258, 
    15.0989309946696, 15.8144754833645, 16.1962887446086, 16.1938959757487, 
    15.4698594411214, 15.5309147304959, 15.4333029852973, 15.2230326334635, 
    15.1915273666382, 14.949490070343, 16.700472301907, 16.595744450887, 
    16.7995482550727, 16.1722103754679, 15.5820879406399, 14.944575521681, 
    14.7628289631435, 14.679020690918, 16.8256736331516, 16.7021617889404, 
    16.6389781104194, 15.6932711071438, 14.9854067696465, 16.5309825473362, 
    16.0329845216539, 15.9251018100315, 14.8757115999858, 14.9297780990601, 
    14.8884220123291, 14.8870038986206, 14.8955249786377, 14.8840341567993, 
    13.2351795832316, 11.0896244049072, 10.2727085749308, 9.39949893951416, 
    33.185001373291, 33.185001373291, 33.1860008239746, 33.1839981079102, 
    33.185001373291, 33.1126670837402, 33.2529983520508, 33.6459999084473, 
    34.0149993896484, 14.7791595458984, 14.617115020752, 14.6057024002075, 
    14.6041698455811, 14.4727430343628, 12.4565010070801, 10.8639149665833, 
    10.0750846862793, 9.47451257705688, 9.07508945465088, 8.74132251739502, 
    8.067458152771, 7.35319900512695, 6.89866304397583, 6.34328508377075, 
    33.1900005340576, 33.1889991760254, 33.1940002441406, 33.189998626709, 
    33.1749992370605, 33.1359996795654, 33.4914989471436, 33.8134994506836, 
    34.1079998016357, 34.1990013122559, 34.2270011901855, 34.2589988708496, 
    34.2700004577637, 34.3019981384277, 34.3190002441406, 0.212599942698479, 
    0.192569131261999, 0.186839991967246, 0.1624202385672, 0.17125966474767, 
    0.152691910106491, 0.146031144711369, 0.176656513774725, 0.1348015039948, 
    0.196810728421345, 0.213358404662935, 0.156765985592722, 
    0.180619047954168, 0.226560081928098, 0.207255486524237, 
    0.196013042496556, 0.153787041517729, 0.212368519736534, 
    0.188540460109794, 0.219034055699219, 0.135877917161369, 
    0.203849114453924, 0.192228451632657, 0.159163592833512, 
    0.220391871304086, 0.132698624667742, 0.193613397121513, 
    0.185316122295004, 0.13873319565751, 0.187544003597041, 
    0.206840486321561, 0.140153379016548, 0.178375476378434, 
    0.189879470447559, 0.131266283973526, 0.192476386362354, 
    0.190877864015158, 0.158797417202507, 0.159229716653604, 
    0.186730455619295, 0.161533416395419, 0.133754848955624, 
    0.203181411961557, 0.181360249032948, 0.176701251530931, 
    0.13724620340712, 0.172981160029312, 0.181072427578701, 
    0.147862717384563, 0.195725181429943, 0.170200980298433, 
    0.0912231296053067, 0.172483917087538, 0.123530239580624, 
    0.171583434476126, 0.213740190417576, 0.164966228226658, 
    0.159621184785021, 0.158900262589309, 0.126065558610503, 
    0.150649242556255, 0.130654465431438, 0.182281570045718, 
    0.220499482447659, 0.0843297692879802, 0.163648368880922, 
    0.124864876720244, 0.163739237794475, 0.171729689857581, 
    0.132089284924213, 0.15085291645908, 0.178807922120056, 
    0.182203255578128, 0.116154925343958, 0.144601868916778, 
    0.125835649954296, 0.176666248764831, 0.194565451964035, 
    0.125656084372902, 0.0951966210946208, 0.154974357650454, 
    0.168772842309619, 0.139275560794601, 0.154757899364474, 
    0.129484572267521, 0.152559342177834, 0.176254276864559, 
    0.186633040052655, 0.125069578592439, 0.121059100148645, 
    0.137982911397246, 0.174034401284763, 0.141161124197121, 
    0.171404984700515, 0.128036341067311, 0.109148560224565, 
    0.164344103597518, 0.171835957308029, 0.178019850639175, 
    0.126770975643962, 0.15612172993088, 0.12310014233588, 0.18427215654897, 
    0.176204986264325, 0.173547243987089, 0.130903852754604, 
    0.127725787316048, 0.151375091860373, 0.179945264085907, 
    0.189834190001491, 0.130580396459516, 0.173335984456374, 
    0.125435480471608, 0.184314576186854, 0.120800315709439, 
    0.196173015628708, 0.18358172736331, 0.135984461231908, 
    0.155981523178682, 0.134354566451351, 0.192457189271989, 
    0.213286255193696, 0.137141906313331, 0.174419436369902, 
    0.134747389131557, 0.177906011191179, 0.127593617173957, 
    0.188946197511486, 0.2003258058779, 0.141387771187489, 0.174471591302939, 
    0.131149743454265, 0.198898887094371, 0.111413908850674, 
    0.229361462292454, 0.14757731753431, 0.183833497382841, 
    0.145608789845189, 0.164105325834176, 0.14647705355381, 
    0.168893903303636, 0.21279306882401, 0.144506790450027, 
    0.169930653567971, 0.139393742478665, 0.200723049149477, 
    0.108039058459723, 0.235911675494728, 0.159236916386634, 
    0.202126190399384, 0.150087874947255, 0.130759577328282, 
    0.158447413422126, 0.152873223372957, 0.0867883385720827, 
    0.217450887006753, 0.148472017344834, 0.167502181064347, 
    0.150592866691246, 0.188429626976068, 0.112689401577857, 0.2316305351423, 
    0.16716879307099, 0.214625496802526, 0.146595718672683, 
    0.0887384103705287, 0.148015362405907, 0.150352481363271, 
    0.0923169915991004, 0.227306005377937, 0.151147851548721, 
    0.181857037975724, 0.152515036510108, 0.152791794382232, 
    0.097626915106148, 0.21784515754257, 0.175607888751122, 
    0.0768635644021609, 0.213144551557534, 0.145429414805772, 
    0.0591345235840816, 0.137063634491517, 0.154285576316962, 
    0.0982554816898909, 0.236893961070653, 0.150344228945373, 
    0.198697856801141, 0.143992565215689, 0.11336875028027, 
    0.0678875739619216, 0.20024688042595, 0.191890905029911, 
    0.0826006524877724, 0.214859411139656, 0.142434625230361, 
    0.0408866853814332, 0.143608556730717, 0.152950605022543, 
    0.0798086852914453, 0.236912834747342, 0.151399295782453, 
    0.0844769135886295, 0.199059280511541, 0.13649857726566, 
    0.0904039626149169, 0.054833184914719, 0.181314832557419, 
    0.203360231123154, 0.0876878547367659, 0.224868661998387, 
    0.136521902285216, 0.0313668759942612, 0.157551731513166, 
    0.143161799241976, 0.0448863754235078, 0.227482082648751, 
    0.161822631885461, 0.0843065941059268, 0.19076073107741, 
    0.129524722250593, 0.077314663230628, 0.0600347162776729, 
    0.169021413559023, 0.199461185237027, 0.0732850952035547, 
    0.234648125274686, 0.13494849011839, 0.0857869061906988, 
    0.045490407671542, 0.158706001903253, 0.127696221619965, 
    0.0335974282708369, 0.208846818227487, 0.173393123072065, 
    0.0857374772630198, 0.194658132897222, 0.1238608864997, 
    0.0723668448102527, 0.0667710625878339, 0.162148670409668, 
    0.187840206390679, 0.0451798019371798, 0.236331112189767, 
    0.140228546192102, 0.0885896922599249, 0.0723596192357564, 
    0.149731236287278, 0.112521201061473, 0.0491173789061043, 
    0.187714857740232, 0.179261985413747, 0.0779430055298373, 
    0.21149088844508, 0.124747954069233, 0.0877922016380722, 
    0.0957436113508148, 0.0716862463378918, 0.145759478285662, 
    0.166482136479877, 0.0388148660149774, 0.222461625356393, 
    0.146043422144331, 0.0927576457934852, 0.094395577686176, 
    0.152338314205216, 0.106802271324462, 0.0660189901140265, 
    0.167860888525907, 0.182138687231461, 0.0625148668043827, 
    0.223265285803411, 0.126146296391452, 0.0937729357053701, 
    0.130197392459757, 0.0805622451543081, 0.10486465234704, 
    0.133694999464701, 0.0590632102049324, 0.195817732496092, 
    0.152449699036794, 0.0851876232528266, 0.11309593872781, 
    0.171517987257798, 0.108693977565871, 0.0885101276634629, 
    0.0722875130311398, 0.141939073110885, 0.165418796214676, 
    0.0580573293761953, 0.213639994441002, 0.122421042522264, 
    0.101915876695454, 0.144648333335375, 0.0933086358163868, 
    0.0568254044936266, 0.112786384096192, 0.0816832052019172, 
    0.163785571143094, 0.161106735327164, 0.0649399319516154, 
    0.131719700648381, 0.187228621414072, 0.103242802065824, 
    0.0991830919553701, 0.07461505596538, 0.092007252787039, 
    0.127512181128934, 0.0699976979083551, 0.187407783709607, 
    0.122632612956361, 0.0875321944868269, 0.141514740519587, 0.103262539826, 
    0.0247494439936839, 0.0873945934217513, 0.121148197250351, 
    0.0874974739686398, 0.125611711050338, 0.152932681712723, 
    0.05607569562586, 0.138169020515048, 0.182391995823147, 
    0.0882332081114841, 0.106815016099751, 0.081241909273943, 
    0.0284309582010843, 0.106241530373731, 0.0862088489111991, 
    0.15801593552704, 0.128883398291666, 0.0545201248269491, 
    0.141259482681558, 0.109791761218426, 0.0043857125965379, 
    0.101596832508043, 0.138820465726932, 0.0793458909263174, 
    0.0691428729042265, 0.121878483619169, 0.0592021209211985, 
    0.123216973194215, 0.163126032650346, 0.0820159000542423, 
    0.0873385604536237, 0.0875045596214472, -0.0163261241250303, 
    0.0865503211102296, 0.11820711185942, 0.0917400671408126, 
    0.122703309875294, 0.126858893801642, 0.0347760667238501, 
    0.146201844540412, 0.11571216639536, -0.0113855810564673, 
    0.105144170970055, 0.128169492304487, 0.0762069666469898, 
    0.00509080927530317, 0.105487135842481, 0.0531266274054616, 
    0.0813687791182764, 0.143862095678848, 0.0925961796155693, 
    0.0478868240456991, 0.0909667081392817, -0.0353075618210043, 
    0.110544291129836, 0.131853806605533, 0.0807901147161291, 
    0.0680032705573078, 0.110105537993245, 0.0258587298121571, 
    0.143089549416845, 0.12066470034339, -0.00337777752377674, 
    0.0859380609457383, 0.0797405364228571, 0.0809657107444941, 
    -0.0353269786172177, 0.0902749823574875, 0.122717152142623, 
    0.0472141807872889, 0.0256529024835687, 0.123127309200045, 
    0.0999163246174781, 0.0110716905031469, 0.0974074177763509, 
    -0.0427439984620037, 0.116192917433645, 0.101177705856158, 
    0.0709501347177028, 0.00708054447174309, 0.103176928253667, 
    0.00288715673934535, 0.121676799412608, 0.115205335007285, 
    0.0346594722523939, 0.0499760540532925, 0.0365795248771256, 
    0.0836827725924067, -0.0475048274460043, 0.116136475570454, 
    0.134353806605533, 0.0550519565523709, -0.0327576762995762, 
    0.0847338799894805, 0.0978918201274395, -0.0262031903538584, 
    0.103050625445822, -0.0328043284932975, 0.104838915039341, 
    0.0214630267708272, 0.072262670526513, -0.0280061768495358, 
    0.0982942389492844, 0.120076443514089, -0.0119601807331553, 
    0.0891109471919628, 0.102423887151548, 0.0603047542551269, 
    -0.000356833527703779, 0.0261639717736745, 0.079810982229476, 
    -0.048591471606535, 0.126089091531774, 0.0846135273893609, 
    0.062403282122079, -0.0792766629615696, 0.034422630033488, 
    0.0997354882198928, -0.0704632155751079, 0.0932669119663942, 
    0.00293418471060767, 0.08249379924541, -0.0443960438569357, 
    0.070147624548214, -0.0344510945689051, 0.11726837254311, 
    0.120688343814853, 0.00713949688739561, 0.0491508383795209, 
    0.0875812806660259, 0.0547112517308683, -0.0684239082552415, 
    0.0391179158937507, 0.0676342130923061, -0.0390079417745474, 
    0.111504138091401, -0.0235919048697978, 0.0631233548202655, 
    -0.0997268451033869, 0.00147501256170948, 0.11451068805994, 
    0.106330539959121, -0.0875633606647959, 0.0628643093255001, 
    0.0273970288749848, 0.0286421405015813, -0.0629875009979665, 
    0.0469654823300767, -0.0271670642487514, 0.122992778055211, 
    0.0579111087031687, 0.0364946066367782, 0.0037758445502225, 
    0.0682237510848011, 0.0450187663398328, -0.132511338207424, 
    0.0672459627969688, 0.0404223685093629, -0.0145458262757206, 
    0.086350184406845, -0.113008714755373, 0.0523752407370296, 
    -0.0845728595157573, -0.00510338749735029, 0.112414265012941, 
    0.0839710535073439, -0.0543412160032293, 0.0228331042071658, 
    0.0159090412786291, -0.0641597412089065, -0.0496573356733888, 
    0.00727040264603179, -0.00987128466090484, 0.102806170562104, 
    -0.0521070330618309, 0.0540855733640889, -0.0323412064852972, 
    0.0465286841958633, 0.108692204430391, 0.0355219813041529, 
    -0.148670524816478, 0.10244819846972, -0.00865348242254689, 
    -0.00110089592970274, 0.0456877651649693, -0.141683179708904, 
    0.0184618434508156, -0.0472321368674927, 0.0063137824839318, 
    0.0985993194000374, 0.0103157138925369, -0.00119124541400305, 
    -0.00793274303730017, -0.00481644656039906, -0.146086526629891, 
    -0.00824544477603002, -0.0404157048700442, 0.00859601949064756, 
    0.0788007459302826, -0.141090934104238, 0.0547995564488219, 
    -0.0372972367668081, 0.0296594215337583, 0.10584583804235, 
    0.00268581028206361, -0.100510863769283, 0.13462278521669, 
    -0.0668547009686154, -0.0162216960260585, -0.0285188130124534, 
    -0.126738176737842, -0.0257239041629776, -0.0141823467545363, 
    0.0354883767690438, 0.081240094763644, -0.0782374488925752, 
    0.0389938680418233, -0.0258177585789707, 0.087059056237032, 
    -0.014469244220697, -0.165537512206547, 0.0474237098420337, 
    -0.0902950043163488, 0.0110109249605596, 0.061607870145438, 
    -0.177107318003082, 0.0350047757410135, -0.0132716386302624, 
    0.0264266635645424, 0.0903788233376498, -0.0518185283561811, 
    -0.0276863272151381, 0.141583251148766, -0.103934787715034, 
    -0.0437480261502428, -0.105492506633772, -0.0802335124029831, 
    -0.0645029395879873, 0.00714045361232655, 0.058970481945987, 
    0.0737892355615101, -0.139731878499435, 0.0593068501499937, 
    -0.0348112820127294, 0.0956956915579755, -0.0256693678795052, 
    -0.119323313106812, 0.0975146962882129, -0.131132327728079, 
    -0.00765137101703385, 0.0178704997316872, -0.171291121335519, 
    0.0113813172368638, 0.0164349507991004, 0.0502028777633764, 
    0.0821508833399804, -0.0937522188010662, 0.0287368028069366, 
    0.104673992101793, -0.115115091342642, 0.0645446962981016, 
    -0.0594275877265563, -0.132630259788553, -0.0165098533903884, 
    -0.0781640245735273, 0.00900482431161937, 0.0566905395775436, 
    0.0853433843127985, -0.172976198189294, 0.0601184537195292, 
    -0.0372045929137839, 0.0942150354958528, -0.0459441227775153, 
    -0.0424606491298663, 0.118668441214405, -0.152231759773772, 
    -0.0479802829283275, -0.0492515093193193, -0.134188986887782, 
    -0.00688120817838031, 0.0346376339784631, 0.0772892495462132, 
    0.0892446073811557, -0.112677319477987, 0.0661350270315066, 
    0.0460981865012321, -0.115495180938511, 0.0849958564573901, 
    -0.0590165358482553, -0.0991982497597393, 0.0478616811514942, 
    -0.0679126140191884, -0.0213195391593495, 0.0324155222002493, 
    0.0800877407671267, -0.182710386959751, 0.0558973084478013, 
    -0.0243751865762781, 0.0924153181544336, -0.0623639870786972, 
    0.0256444373090725, 0.0912681059136325, -0.156974685471693, 
    0.0442432526016787, -0.0863495085603242, -0.0872835801010528, 
    -0.0746379596407106, -0.00348372993153055, 0.0314619602513589, 
    0.0763240161044408, 0.115756052067633, -0.123014332169004, 
    0.087461473912577, 0.0171020012619889, -0.115217135638393, 
    0.0943319729489141, -0.0536974186759529, -0.0299716446577413, 
    0.0873708337925302, -0.0617708531230524, -0.0642068845896527, 
    -0.0256830125137786, 0.0398348647067075, -0.16062103384361, 
    0.0547435476809949, -0.00218490243992556, 0.102168801717093, 
    -0.0746326931352005, 0.0696240140900393, 0.0361023937316997, 
    -0.156588936444514, 0.0766140099947058, -0.0941911084231147, 
    -0.0698757399941144, -0.0041565169607127, 0.0114747161845069, 
    -0.00166988432033166, 0.0470633139099867, 0.133121813092228, 
    -0.135755911670089, 0.0972992082776693, 0.025367814177696, 
    -0.107716251029403, 0.0938964991747171, -0.0492876626158066, 
    0.0351160162440884, 0.0782845548882419, -0.0739068850083846, 
    0.0451003387833193, -0.0822611611723553, -0.0931158496226017, 
    0.00290822841658495, -0.110825776895376, 0.0705999797852665, 
    0.0108462488488515, 0.126484659245367, -0.0881312490903048, 
    0.0904203706390785, 0.00432910888308123, -0.156352876138038, 
    0.0916500175663526, -0.0839965545439225, -0.0112840531050068, 
    0.0534895375357919, 0.0119623327935335, -0.0437916963033693, 
    -0.0128314106110337, 0.118064631001535, -0.135365014364471, 
    0.105820566910339, 0.0303113309508253, -0.090912319432113, 
    0.0985504419044934, -0.0537791164750444, 0.0665977201146679, 
    0.0363779674621684, -0.0985074491212009, 0.0775267907564246, 
    -0.0590928170494807, -0.121592024627609, 0.00320159649008188, 
    -0.0492773873818161, 0.0829020233134131, 0.00630694131050501, 
    0.140084245953556, -0.105636481150035, 0.100390246117452, 
    0.00586701652535115, -0.151902667968029, 0.0887951773026146, 
    -0.07382324399899, 0.048341266488229, 0.068244658777988, 
    -0.0128724688103557, 0.047363113323875, -0.0629085949563844, 
    -0.0802930287314033, 0.0902571048188344, -0.116384511085524, 
    0.126648752006957, 0.0114029193163233, -0.0691658055945079, 
    0.110545271329771, -0.0650527883969454, 0.0707320983361994, 
    0.00494113891237812, -0.124265238415449, 0.0997931755253369, 
    -0.0340760232195748, -0.114884985838445, 0.0330085760014328, 
    0.00851530407757918, 0.0702669287407992, -0.0269274165269166, 
    0.125950983540598, -0.115375588727231, 0.111872419670727, 
    0.00227571239498797, -0.143403990408176, 0.0819018788215322, 
    -0.0693323065008059, 0.0691859159154491, 0.0433463071197936, 
    -0.0577059281873746, 0.0746690208633865, -0.0408275921421037, 
    -0.116278206421958, 0.0784395688705087, -0.0923776757681495, 
    0.13294144167469, -0.0218066954048127, -0.0483968855937918, 
    0.113467987717939, -0.0818739689430042, 0.077685164474357, 
    -0.00627012947074257, -0.137328783324833, 0.104720775447146, 
    -0.031408194516804, -0.10722624759526, 0.0611843106337311, 
    0.0380413908959471, 0.0310270673224568, 0.0429429914763443, 
    -0.0716072846559777, 0.0986280764985217, -0.103180846266031, 
    0.127499656305852, -0.0184419722232853, -0.125083343112372, 
    0.0828186431925622, -0.0632060760789571, 0.0601128966760431, 
    0.0152616110538719, -0.101177645704279, 0.103475780388158, 
    -0.0194913708219633, -0.110269104644512, 0.0730296348678434, 
    -0.0680763458217148, 0.108331268793595, -0.0462893870630766, 
    -0.0468694331284791, 0.10001094695184, -0.0980512173893402, 
    0.0910621874868995, -0.0200189043042309, -0.134384340957514, 
    0.0954110951301259, -0.100655994911529, 0.0644342654674867, 
    0.0301023922508332, -0.0277155412244841, 0.0464626084752208, 
    -0.0939884889578605, 0.0802324765853525, -0.0820614057159447, 
    0.11825483843507, -0.0391164252833186, -0.0965133672034531, 
    0.0943796587955442, -0.0645462763211706, 0.0593169393767008, 
    -0.00372496394509453, -0.121607065857804, 0.117238747188321, 
    -0.00659494731126046, -0.0922768180526139, 0.0493610247411094, 
    -0.0394109388562407, 0.0649010527927174, 0.0470744612029068, 
    -0.0577982933209897, -0.0601992036012902, 0.0760004437509048, 
    -0.0931112661879064, 0.097461671436477, -0.0373399824771916, 
    -0.120666430572616, 0.0899266449015466, -0.0855298255248363, 
    0.0505319742571117, 0.0123009718235624, -0.078818331739435, 
    0.0635239054360527, -0.0826700915261183, 0.0624542259322965, 
    -0.0654251758671661, 0.0928283767129976, -0.0485401082541421, 
    -0.0728342728924371, 0.104125342713045, -0.0765212843132895, 
    0.062116264635337, -0.0215230318639828, -0.121052149857672, 
    0.107122070647712, -0.0808185485290903, 0.0241674585061501, 
    -0.0283505123595164, 0.013115699371735, 0.0471599351353772, 
    -0.0579774533606919, -0.0634902894949699, 0.0561753245644529, 
    -0.075071964797976, 0.0806043962903054, -0.0417650458887874, 
    -0.104631442957508, 0.101629414654919, -0.0753886007534449, 
    0.032221250078498, -0.000405695948841567, -0.103545847596085, 
    0.080606179072071, -0.0655681105121444, 0.0252785357274377, 
    -0.0418366731985671, 0.0677628815662848, 0.0561708333513106, 
    -0.0512248567972115, -0.0603253751146246, 0.0897112953039367, 
    -0.0759711341372464, 0.0515891738778832, -0.0352952181302211, 
    -0.110107371796993, 0.0914246077238198, -0.0793116610088547, 
    0.00509556585513413, -0.0222581016959416, -0.0306198798793254, 
    0.0578433634438653, -0.0601279632789866, -0.0489535082741651, 
    0.0379165200751214, -0.0617356006718536, 0.0595897114761648, 
    -0.0351479268576577, -0.0918230142931075, 0.115713324890779, 
    -0.0742024972307032, -0.00451520679631327, -0.0129953073378032, 
    -0.112458247269781, 0.0772561712140156, -0.054254926984503, 
    -0.0104388647360375, -0.0381190125374193, 0.0475851941609274, 
    0.0648227360730963, -0.0553467626832331, -0.0481572567174697, 
    0.0549484492434983, -0.0662620484143279, 0.0262786821789773, 
    -0.0340355222636342, -0.0986273186992354, 0.0919527307374278, 
    -0.0888884969391996, -0.0368089544357442, -0.00855709039348918, 
    -0.06051214740023, 0.0683086632029305, -0.0441578932269881, 
    0.00611219044757472, -0.0405123628958326, 0.0396490554823868, 
    0.0607050318292112, -0.0285962252054147, -0.0800466585496452, 
    0.100564414200421, -0.065254214730441, -0.0538084718701733, 
    -0.0269573087881189, -0.115000102509884, 0.0594321893330042, 
    -0.0494825705901361, -0.0428603667620533, -0.0371225399576368, 
    0.0252654015981332, 0.0738909241637195, -0.0312148580698463, 
    0.0231099644158261, -0.0614565443709571, 0.00793779497225861, 
    -0.0871360126582197, 0.0983612821830744, -0.0885137032311289, 
    -0.11241765224717, -0.00482759404121512, -0.0816066720367744, 
    0.0618237371319845, -0.0494642775704404, -0.0291099553420813, 
    -0.041579095545232, 0.0171400240115436, 0.0793543138789188, 
    -0.04312187865003, -0.062598610911551, 0.0561245967044358, 
    -0.0636566680781261, -0.0901600707468136, -0.0238467158000905, 
    -0.114260405857439, 0.0398099496535075, -0.0618802533535043, 
    -0.10155657406465, -0.00231511464995466, 0.0752103395041276, 
    -0.0346209128235062, -0.00555256005541232, -0.00588988494730074, 
    0.0617130274346799, -0.0746344066706165, 0.085219581594417, 
    -0.0730055287317548, -0.181868665732583, -0.0201383198567652, 
    -0.100194159618408, 0.0435390924091762, -0.0496797141448236, 
    -0.0712715910659562, -0.0459450192056837, -0.00512280424802208, 
    0.0904346784832138, -0.0315532525673187, 0.011906351134576, 
    -0.0710545299555481, -0.103538540338852, -0.101514979943376, 
    0.0212286645638935, -0.0734358490497304, -0.175986530420999, 
    -0.0273520785551247, 0.0618023482476705, -0.0540322166007847, 
    -0.0373300719759971, -0.0241287442990032, 0.0731079759882938, 
    -0.0537708316889471, 0.0472603387103085, -0.0771601349940996, 
    -0.206448217307488, -0.0414527756968616, -0.117953400129699, 
    0.0217546823195233, -0.0600481305507701, -0.137240157636851, 
    -0.0186133546757973, 0.0894358804898526, -0.00707893914496135, 
    -0.0216437160612717, -0.110231052729149, 0.0661062801665477, 
    -0.0750534130182729, 0.0153462353453495, -0.0804836743062159, 
    -0.22445579341813, -0.0485537285080542, 0.0391506285877051, 
    -0.062358754884781, -0.0766131918867235, -0.0399009414550534, 
    0.0768072065593857, -0.0190246638337283, 0.00104761682208946, 
    -0.20963326814997, -0.115973980603232, -0.000230380846262968, 
    -0.073180111745043, -0.196900435633527, -0.0303901257098735, 
    0.0732596012807356, -0.00216163807914405, -0.0516093993685752, 
    -0.111234273878351, 0.0669357297982892, -0.0379238163080876, 
    0.0153549194080557, -0.234828802024284, -0.0795200613045014, 
    0.0129960244731884, -0.0694401887736173, -0.110563325840431, 
    -0.0410834474492346, 0.07410568029454, 0.00501187493042585, 
    -0.0394435209303991, -0.213467509547701, 0.04738910583934, 
    -0.0818239983326247, -0.0105694445862912, -0.218286905968869, 
    -0.0453567465974659, 0.0372830154731377, -0.0398499540621203, 
    -0.0805440085371141, -0.09604428187144, 0.0592069551085165, 
    0.00540053758228723, -0.00213913836414011, -0.234195493491767, 
    -0.105657707207722, -0.0127546729834938, -0.116740936965002, 
    -0.0445933117450299, 0.0607280155873761, 0.00948237365536357, 
    -0.068769039786403, -0.194103833113895, 0.0294459724632242, 
    -0.0325641742249566, -0.0143572998302256, -0.222505603441136, 
    -0.0655928233039834, -0.0135563355479066, -0.0680276194103311, 
    -0.0925822162212905, -0.0709864009027309, 0.0499526799382996, 
    0.0180735509558164, -0.0341801347563096, -0.233404643336763, 
    0.015891760868637, -0.101563514161697, -0.0332699645426877, 
    -0.107200558488745, -0.0516683921052784, 0.0250982620551691, 
    -0.0331732885190191, -0.0864938165814718, -0.142364668398839, 
    0.0134907582939958, 0.00871474730410384, -0.0250799647801557, 
    -0.225816930904478, -0.0772651382873746, -0.0596697344206046, 
    -0.077671570509924, -0.0687157018440337, 0.0357568459302097, 
    0.00578745788387907, -0.0631311749106654, -0.205259228621708, 
    -0.00343687055435381, -0.0693419519124615, -0.0487999067465645, 
    -0.107466501927213, -0.0540950205696083, -0.031648223975641, 
    -0.085651275010767, -0.0917233354560615, 0.00563703228343506, 
    0.00811851624527355, -0.0353471269438095, -0.224257195135527, 
    -0.0394003164929176, -0.0803807952760972, -0.0886116922395639, 
    -0.0610698822192139, -0.0791190760213127, 0.00327330222658251, 
    -0.090856934303305, -0.145677198916417, -0.0124504038153792, 
    -0.0287264825318385, -0.059241509549328, -0.123394422053683, 
    -0.0478713699768278, -0.0854003252409171, -0.0640463823745674, 
    -0.0789483954252614, -0.00679320724223304, -0.0200370417891714, 
    -0.0448409222251185, -0.193067683935661, -0.0641158089093891, 
    -0.0699670943549873, -0.0994220887792265, -0.0615659281967441, 
    -0.074200483490128, -0.0503374082250916, -0.108678129929549, 
    -0.0954399187080147, -0.00955797504078358, -0.052842665670481, 
    -0.133389862065907, -0.0544997838941716, -0.0473020294069567, 
    -0.118428586770814, -0.0447597575604469, -0.0961847253795878, 
    -0.032756670379454, -0.0766110236587738, -0.133800417612521, 
    -0.0671913844067424, -0.0925361874233121, -0.0747802252763389, 
    -0.056310369482163, -0.103030997313027, -0.109910885614386, 
    -0.0843931891264333, -0.0130343571445766, -0.0431450150378105, 
    -0.118170918083353, -0.0816499686934558, -0.0478851851752998, 
    -0.126514526523367, -0.04214708337839, -0.106703068273208, 
    -0.0658644481281602, -0.117897642869002, -0.0925040375199039, 
    -0.051304687237391, -0.0793981236549709, -0.0860970764213753, 
    -0.0684040502515935, -0.0483013513879497, -0.138173857655829, 
    -0.109498015530385, -0.0993097253795879, -0.0315825065610944, 
    -0.0677099996116547, -0.099573324005355, -0.0867928861482574, 
    -0.111849389327609, -0.0510423297953734, -0.0938009761158289, 
    -0.0907540319695819, -0.141494595331183, -0.0885414153836671, 
    -0.0350418427255168, -0.0751053811779882, -0.0911616407396033, 
    -0.0967851615645494, -0.148109263576494, -0.113207210373704, 
    -0.113770176427505, -0.0534245677570663, -0.119066198900008, 
    -0.10559444879555, -0.0715587891949905, -0.0915297764870021, 
    -0.0617722930091569, -0.0896706550246361, -0.0860557443100122, 
    -0.097961899733228, -0.155420561917103, -0.097659542759149, 
    -0.0263606585854969, -0.091110337675674, -0.105281942169417, 
    -0.103283975015445, -0.129861075747254, -0.11370244647679, 
    -0.113137829143173, -0.0634090612664569, -0.160351565233906, 
    -0.124258169432751, -0.0513951878471788, -0.0797831155529881, 
    -0.081634787696809, -0.114618930587339, -0.0876119973151953, 
    -0.166885036301439, -0.105836763430247, -0.0177065712723066, 
    -0.126255197038208, -0.129047207584613, -0.088965405405928, 
    -0.0992152789691814, -0.111335326921726, -0.0820888679152613, 
    -0.112317035813918, -0.0571591348406498, -0.185506175090125, 
    -0.124950148999044, -0.0326782981407527, -0.0847698530565334, 
    -0.117726115931053, -0.109513229377368, -0.0710479220348001, 
    -0.166086174504133, -0.106190135916662, -0.00549898714503639, 
    -0.162112626718784, -0.141806082030407, -0.065300064556163, 
    -0.073670190198921, -0.12047089072895, -0.100082645186949, 
    -0.0423475625007422, -0.198182655089694, -0.108794690079121, 
    -0.0103623178581545, -0.108251351823365, -0.14620636018091, 
    -0.0809954298047246, -0.0582829854442793, -0.152188293230319, 
    -0.0616822752975348, 0.00479040506824083, -0.180969171389469, 
    -0.12866520637209, -0.0388994590294244, -0.0653275283053829, 
    -0.137966897651409, -0.0900070037914307, -0.0324848422008156, 
    -0.195767822707813, 0.0106511565037822, -0.131748246835972, 
    -0.143675779190502, -0.0500729976636619, -0.0508208176853535, 
    -0.14177933189106, -0.0691792627153728, 0.0124303046471256, 
    -0.177074357197241, -0.0997279176181835, -0.0104578378776857, 
    -0.0792804623509891, -0.135188077801881, -0.0578589857129277, 
    -0.0340678975536544, -0.178308402802579, -0.0618313536666755, 
    0.0183421295276062, -0.139244165285953, -0.115445887897359, 
    -0.0309799164640545, -0.0507656886318991, -0.140562875434613, 
    -0.0684147202100926, 0.0136031741880422, -0.164364998327278, 
    -0.088164871710991, 0.0113414641209698, -0.0945613688087048, 
    -0.0999383636907906, -0.0310899959546775, -0.0447113511326191, 
    -0.156059689266054, -0.0604878564653727, 0.0155286469850242, 
    -0.129856949970678, -0.0808026589221384, -0.0216451360456972, 
    -0.0601832528044585, -0.130063260907349, -0.052650788056375, 
    -0.00133406817651547, -0.154873107063183, -0.0692880126454172, 
    0.0136993377795594, -0.0952771596858022, -0.066521104730452, 
    -0.0243763703214763, -0.0588211085537743, -0.143493163750598, 
    -0.0574373947706396, 0.00750756354198772, -0.116672279821419, 
    -0.0684350103136412, -0.0154585658831343, -0.071459339888226, 
    -0.0913746735052436, -0.0407878567659959, -0.0298455093556456, 
    -0.150254112740138, -0.0503358744081328, 0.00244499830338362, 
    -0.0847340874414644, -0.0255602361433535, -0.0744950814177398, 
    -0.13499736889067, -0.0445358588571562, -0.00906417446079648, 
    -0.112319396125683, -0.0911851429041826, -0.0148164655108956, 
    -0.0769575170512615, -0.0552895678652178, -0.0390720922941164, 
    -0.0656406592472309, -0.148151140145609, -0.0345383548174773, 
    -0.0103348436845749, -0.0760286115906381, -0.0220494472307906, 
    -0.086679829390179, -0.105920942126029, -0.0340396573031053, 
    -0.0370121869010767, -0.119055992622951, -0.0580699492469764, 
    -0.0186944368465569, -0.0772588231791748, -0.0351026057741413, 
    -0.103241497543151, -0.131093813716077, -0.0136852932346342, 
    -0.0256698568338434, -0.0818730014623406, -0.125240380221514, 
    -0.0146080304523018, -0.0913186315532146, -0.0736159553687818, 
    -0.0309754736417727, -0.0740213260504744, -0.12460652344639, 
    -0.0266134025567114, -0.0284615378207398, -0.0768928398235867, 
    -0.0263146988440646, -0.126733447620655, -0.0854163328201741, 
    0.00140215111451796, -0.0511859234733423, -0.101023918812267, 
    -0.0872945804748655, -0.00890378743249437, -0.090441959165503, 
    -0.029349889709688, -0.113083215270805, -0.104171664057874, 
    0.00118271322535027, -0.0462346137609926, -0.0886396344803627, 
    -0.0168288437579826, -0.124208270447901, -0.0417727979012361, 
    0.000162298925750664, -0.086022668823912, -0.111129968170324, 
    -0.0488647607270571, -0.0197739462680056, -0.0899918998821803, 
    -0.0281510941077366, -0.137440362316942, -0.0506873289139241, 
    0.0124512289771245, -0.0787666008340579, -0.116527666260296, 
    -0.0117794815918224, -0.105987287511847, -0.0200340176209913, 
    -0.0112219167767725, -0.12296236566143, -0.0875664313468761, 
    -0.0231964016216429, -0.0473056281652895, -0.0961197980545814, 
    -0.0283895127032951, -0.134815087487938, 0.00307110468665448, 
    -6.38382296024986e-05, -0.120124736738472, -0.140661408251265, 
    -0.022421874151389, -0.099709955161841, -0.0221447829920016, 
    -0.146126122814989, -0.0258213128493742, -0.0204647490592673, 
    -0.0853072807656986, -0.113473314453655, -0.0294917313476817, 
    -0.115254840635868, 0.010337839068462, -0.0155624338149381, 
    -0.155738202372373, -0.130892252932326, -0.0464535723222468, 
    -0.107731750791379, -0.031348766611388, -0.14495974080825, 
    0.0391899494469559, -0.0342786849511613, -0.124083324384956, 
    -0.137568299120406, -0.0364962760068579, -0.108259138461534, 
    -0.0209888553279368, -0.168811079627367, -0.0797371918078711, 
    -0.0770381260090228, -0.11271204615583, -0.0385519236532721, 
    -0.126914386534306, 0.0508284220333479, -0.0407805328303598, 
    -0.155846844950498, -0.146052470217482, -0.0484308062089656, 
    -0.116870043172654, -0.0235180431746326, -0.158780279162097, 
    -0.0132875828278238, -0.106076048836427, -0.119052149326779, 
    -0.0402897639227401, -0.118296827670518, -0.0361563395141977, 
    -0.165860945350023, -0.122886148106699, -0.0630261326008196, 
    -0.122550360673447, -0.0310896999723763, -0.131253204751859, 
    0.0184919349798425, -0.127087945537322, -0.125539427641385, 
    -0.036624870515175, -0.125029985799608, -0.0355699213182895, 
    -0.15310721397655, -0.0754947666657144, -0.0796002187583019, 
    -0.124808513011374, -0.0346357830396959, -0.106966981939024, 
    -0.135210468481689, -0.118982365206712, -0.0321226510578052, 
    -0.132410132401963, -0.0462963693333188, -0.122498169351468, 
    -0.0450098045221106, -0.0975823303029465, -0.126621566472464, 
    -0.0305199924153339, -0.101269931489404, -0.127324080293082, 
    -0.0919071751430006, -0.0389361603751569, -0.137736674632467, 
    -0.0569469865842275, -0.094687166265196, -0.0743182818509778, 
    -0.113376514624267, -0.120128285776072, -0.027154781624956, 
    -0.110837895586576, -0.104015029160364, -0.0599775108510164, 
    -0.0608907817070922, -0.140742660222464, -0.0603201279676582, 
    -0.0871430393995601, -0.119163985078238, -0.0953484145035084, 
    -0.0360702744969016, -0.122156347964998, -0.0864705959475676, 
    -0.0604223024500774, -0.0929704488153946, -0.135983693490916, 
    -0.0601844097446401, -0.0997288867975137, -0.111282332627161, 
    -0.0582630921513004, -0.0641817973697749, -0.122136860706985, 
    -0.0914323745641206, -0.12141493806665, -0.112537440382415, 
    -0.0675180976496035, -0.117168097232576, -0.106919204346005, 
    -0.0450502336848722, -0.10556512963921, -0.115464767968473, 
    -0.122155584451712, -0.139564685563659, -0.0711795045048161, 
    -0.0908263502255499, -0.117835865833938, -0.119122041312167, 
    -0.146236334223229, -0.106556749235665, -0.157312540677194, 
    -0.155190689640931, -0.0487530840266691, -0.127009511248762, 
    -0.106708664452848, -0.150703558084525, -0.177301839693579, 
    -0.0894004394874331, -0.169370220994206, -0.170146985466184, 
    -0.158204311414673, -0.0975092028489468, -0.180599283841257, 
    -0.196444079122413, -0.0785797192791569, -0.157804017935279, 
    -0.182180874009614, -0.174968543621036, -0.0882862427100893, 
    -0.184992016648503, -0.202810439644986, -0.133105488497221, 
    -0.183275144499571, -0.185725161691657, -0.0876727368572819, 
    -0.167546754751685, -0.191447358450373, -0.107570014479312, 
    -0.172513107006255, -0.18741050096419, -0.0983527185533028, 
    -0.137693501192534, -0.170734301669822, -0.100561052127719, 
    -0.154384726215119, -0.173844664808549, -0.108596930983218, 
    -0.162051741830596, -0.11261825304721, -0.12164132467203, 
    -0.162515140945505, -0.103719468875766, -0.154917165971101, 
    -0.0864605932026787, -0.168344277971129, -0.118757474238616, 
    -0.11834502907645, -0.0832122670212821, -0.170947922932055, 
    -0.0666492869762032, -0.128208841447852, -0.058881078592658, 
    -0.0600248899686703, -0.0955820169376288, -0.0415603455434485 ;

 obs_lon = -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -125.983334859212, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.987879897609, -125.983334859212, 
    -125.947621663411, -125.833333333333, -125.961906069801, 
    -125.953334554036, -125.945834477743, -125.983334859212, 
    -126.083333333333, -126.047619047619, -125.983334859212, 
    -126.003334554036, -125.983334859212, -125.987879897609, 
    -125.987879897609, -125.996971361565, -125.983334859212, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.678786769058, -125.683331807454, -125.683331807454, 
    -125.71333211263, -125.647618611654, -125.673331197103, 
    -125.799997965495, -125.749997456868, -125.745831807454, 
    -125.683331807454, -125.733331589472, -125.66333211263, 
    -125.683331807454, -125.683331807454, -125.808331807454, 
    -125.653331502279, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.366668701172, -125.333333333333, -125.333333333333, 
    -125.350001017253, -125.3047601609, -125.358334859212, -125.40000406901, 
    -125.233327229818, -125.316665649414, -125.433339436849, 
    -125.283330281576, -125.31333211263, -125.299997965495, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.320832570394, -125.333333333333, -125.333333333333, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.988889906141, -124.983334859212, -124.933333333333, 
    -124.996971361565, -124.988889906142, -124.961906069801, 
    -125.047621227446, -125.133336385091, -125.083333333333, 
    -124.933335622152, -125.000001695421, -124.966668023003, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.683331807454, 
    -124.683331807454, -124.683331807454, -124.683331807454, 
    -124.683331807454, -124.683331807454, -124.683331807454, 
    -124.683331807454, -124.683331807454, -124.683331807454, 
    -124.683331807454, -124.683331807454, -124.753331502279, 
    -124.733332316081, -124.696968309807, -124.733331589472, 
    -124.747618175688, -124.633336385091, -124.799997965495, 
    -124.708331425985, -124.696968309807, -124.683331807454, 
    -124.683331807454, -124.683331807454, -124.683331807454, 
    -124.696968309807, -124.745831807454, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.37333577474, -124.383336385091, -124.383336385091, 
    -124.433339436849, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -123.983334859212, -123.983334859212, -123.983334859212, 
    -123.983334859212, -123.983334859212, -123.983334859212, 
    -123.983334859212, -123.996971361565, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.683331807454, -123.683331807454, 
    -123.683331807454, -123.683331807454, -123.683331807454, 
    -123.683331807454, -123.683331807454, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -122.983334859212, 
    -122.983334859212, -122.983334859212, -122.983334859212, 
    -123.013335164388, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.683331807454, -122.683331807454, -122.696968309807, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.345834096273, 
    -122.345834096273, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.045834859212, 
    -121.633331298828, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.633331298828, -121.633331298828, 
    -121.673329671224, -121.333333333333, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.333333333333, 
    -121.333333333333, -121.033335367839, -121.033335367839, 
    -121.033335367839, -121.033335367839, -121.033335367839, 
    -121.033335367839, -121.033335367839, -121.033335367839, 
    -121.033335367839, -121.033335367839, -121.033335367839, 
    -121.033335367839, -121.083333333333, -121.083333333333, 
    -120.633331298828, -120.633331298828, -120.633331298828, 
    -120.633331298828, -120.633331298828, -120.633331298828, 
    -120.633331298828, -120.633331298828, -120.633331298828, 
    -120.633331298828, -120.645831425985, -120.633331298828, 
    -120.333333333333, -120.333333333333, -120.333333333333, 
    -120.333333333333, -120.333333333333, -120.333333333333, 
    -120.333333333333, -120.333333333333, -120.333333333333, 
    -120.333333333333, -120.320832570394, -120.333333333333, 
    -120.033335367839, -120.033335367839, -120.033335367839, 
    -120.033335367839, -120.033335367839, -120.033335367839, 
    -120.033335367839, -120.033335367839, -120.033335367839, 
    -120.033335367839, -120.033335367839, -120.033335367839, 
    -119.633331298828, -119.633331298828, -119.633331298828, 
    -119.633331298828, -119.633331298828, -119.633331298828, 
    -119.633331298828, -119.633331298828, -119.633331298828, 
    -119.633331298828, -119.633331298828, -119.333333333333, 
    -119.333333333333, -119.333333333333, -119.333333333333, 
    -119.333333333333, -119.333333333333, -119.333333333333, 
    -119.333333333333, -119.333333333333, -119.333333333333, 
    -119.333333333333, -119.033335367839, -119.033335367839, 
    -119.033335367839, -119.033335367839, -119.033335367839, 
    -119.033335367839, -119.033335367839, -119.033335367839, 
    -119.033335367839, -119.033335367839, -119.033335367839, 
    -118.633331298828, -118.633331298828, -118.633331298828, 
    -118.633331298828, -118.633331298828, -118.633331298828, 
    -118.633331298828, -118.633331298828, -118.620831807454, 
    -118.633331298828, -118.333333333333, -118.333333333333, 
    -118.333333333333, -118.333333333333, -118.333333333333, 
    -118.333333333333, -118.333333333333, -118.333333333333, 
    -118.333333333333, -118.033335367839, -118.033335367839, 
    -118.033335367839, -118.033335367839, -118.033335367839, 
    -118.033335367839, -118.033335367839, -118.033335367839, 
    -118.045834859212, -117.633331298828, -117.633331298828, 
    -117.633331298828, -117.633331298828, -117.633331298828, 
    -117.633331298828, -117.661903018043, -117.693330891927, 
    -117.333333333333, -117.333333333333, -117.333333333333, 
    -117.333333333333, -117.333333333333, -117.033335367839, 
    -117.033335367839, -117.033335367839, -117.083333333333, 
    -128.625340779622, -128.625340779622, -128.625340779622, 
    -128.625340779622, -128.625340779622, -128.625340779622, 
    -128.625340779622, -128.625340779622, -128.625340779622, 
    -128.625340779622, -128.625340779622, -128.625340779622, 
    -128.625340779622, -128.625340779622, -128.625340779622, 
    -128.625340779622, -128.625340779622, -128.625340779622, 
    -128.625340779622, -128.625340779622, -128.625340779622, 
    -128.625340779622, -128.625340779622, -128.625340779622, 
    -128.625340779622, -128.625340779622, -128.625340779622, 
    -128.625340779622, -128.625340779622, -128.625340779622, 
    -128.625340779622, -128.625340779622, -128.625340779622, 
    -128.625340779622, -128.625340779622, -128.625340779622, 
    -128.625340779622, -128.625340779622, -127.52333577474, -127.52333577474, 
    -127.52333577474, -127.52333577474, -127.52333577474, -127.52333577474, 
    -127.52333577474, -127.52333577474, -127.52333577474, -127.52333577474, 
    -127.52333577474, -127.52333577474, -127.52333577474, -127.52333577474, 
    -127.52333577474, -127.52333577474, -127.52333577474, -127.52333577474, 
    -127.52333577474, -127.52333577474, -127.52333577474, -127.52333577474, 
    -127.52333577474, -127.52333577474, -127.52333577474, -127.52333577474, 
    -127.52333577474, -127.52333577474, -127.52333577474, -127.52333577474, 
    -127.52333577474, -127.52333577474, -127.52333577474, -127.52333577474, 
    -127.52333577474, -127.52333577474, -127.52333577474, -127.52333577474, 
    -127.52333577474, -127.52333577474, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.983334859212, -125.987879897609, 
    -125.983334859212, -125.947621663411, -125.833333333333, 
    -125.958333333333, -125.953334554036, -125.945834477743, 
    -125.983334859212, -126.083333333333, -126.047619047619, 
    -125.983334859212, -126.003334554036, -125.983334859212, 
    -125.987879897609, -126.003334554036, -125.996971361565, 
    -125.983334859212, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.683331807454, -125.678786769058, -125.683331807454, 
    -125.683331807454, -125.71333211263, -125.647618611654, 
    -125.673331197103, -125.799997965495, -125.749997456868, 
    -125.745831807454, -125.683331807454, -125.733331589472, 
    -125.66333211263, -125.683331807454, -125.683331807454, 
    -125.799997965495, -125.653331502279, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.37333577474, -125.333333333333, 
    -125.333333333333, -125.350001017253, -125.3047601609, -125.358334859212, 
    -125.40000406901, -125.233327229818, -125.316665649414, 
    -125.433339436849, -125.283330281576, -125.31333211263, 
    -125.299997965495, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.320832570394, -125.333333333333, 
    -125.333333333333, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.988889906141, -124.983334859212, 
    -124.933333333333, -124.996971361565, -124.988889906142, 
    -124.961906069801, -125.047621227446, -125.133336385091, 
    -125.083333333333, -124.933335622152, -125.000001695421, 
    -124.966668023003, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.683331807454, -124.683331807454, -124.683331807454, 
    -124.683331807454, -124.683331807454, -124.683331807454, 
    -124.683331807454, -124.683331807454, -124.683331807454, 
    -124.683331807454, -124.683331807454, -124.683331807454, 
    -124.753331502279, -124.733332951864, -124.696968309807, 
    -124.733331589472, -124.747618175688, -124.633336385091, 
    -124.799997965495, -124.708331425985, -124.696968309807, 
    -124.683331807454, -124.683331807454, -124.683331807454, 
    -124.683331807454, -124.696968309807, -124.745831807454, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.37333577474, -124.383336385091, 
    -124.383336385091, -124.433339436849, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -123.983334859212, -123.983334859212, 
    -123.983334859212, -123.983334859212, -123.983334859212, 
    -123.983334859212, -123.983334859212, -123.996971361565, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.683331807454, 
    -123.683331807454, -123.683331807454, -123.683331807454, 
    -123.683331807454, -123.683331807454, -123.683331807454, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -122.983334859212, -122.983334859212, -122.983334859212, 
    -122.983334859212, -123.013335164388, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.683331807454, -122.683331807454, 
    -122.696968309807, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.345834096273, -122.345834096273, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.045834859212, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.673329671224, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.033335367839, 
    -121.033335367839, -121.033335367839, -121.033335367839, 
    -121.033335367839, -121.033335367839, -121.033335367839, 
    -121.033335367839, -121.033335367839, -121.033335367839, 
    -121.033335367839, -121.033335367839, -121.083333333333, 
    -121.083333333333, -120.633331298828, -120.633331298828, 
    -120.633331298828, -120.633331298828, -120.633331298828, 
    -120.633331298828, -120.633331298828, -120.633331298828, 
    -120.633331298828, -120.633331298828, -120.645831425985, 
    -120.633331298828, -120.333333333333, -120.333333333333, 
    -120.333333333333, -120.333333333333, -120.333333333333, 
    -120.333333333333, -120.333333333333, -120.333333333333, 
    -120.333333333333, -120.333333333333, -120.320832570394, 
    -120.333333333333, -120.033335367839, -120.033335367839, 
    -120.033335367839, -120.033335367839, -120.033335367839, 
    -120.033335367839, -120.033335367839, -120.033335367839, 
    -120.033335367839, -120.033335367839, -120.033335367839, 
    -120.033335367839, -119.633331298828, -119.633331298828, 
    -119.633331298828, -119.633331298828, -119.633331298828, 
    -119.633331298828, -119.633331298828, -119.633331298828, 
    -119.633331298828, -119.633331298828, -119.633331298828, 
    -119.333333333333, -119.333333333333, -119.333333333333, 
    -119.333333333333, -119.333333333333, -119.333333333333, 
    -119.333333333333, -119.333333333333, -119.333333333333, 
    -119.333333333333, -119.333333333333, -119.033335367839, 
    -119.033335367839, -119.033335367839, -119.033335367839, 
    -119.033335367839, -119.033335367839, -119.033335367839, 
    -119.033335367839, -119.033335367839, -119.033335367839, 
    -119.033335367839, -118.633331298828, -118.633331298828, 
    -118.633331298828, -118.633331298828, -118.633331298828, 
    -118.633331298828, -118.633331298828, -118.633331298828, 
    -118.620831807454, -118.633331298828, -118.333333333333, 
    -118.333333333333, -118.333333333333, -118.333333333333, 
    -118.333333333333, -118.333333333333, -118.333333333333, 
    -118.333333333333, -118.333333333333, -118.033335367839, 
    -118.033335367839, -118.033335367839, -118.033335367839, 
    -118.033335367839, -118.033335367839, -118.033335367839, 
    -118.033335367839, -118.045834859212, -117.633331298828, 
    -117.633331298828, -117.633331298828, -117.633331298828, 
    -117.633331298828, -117.633331298828, -117.661903018043, 
    -117.693330891927, -117.333333333333, -117.333333333333, 
    -117.333333333333, -117.333333333333, -117.333333333333, 
    -117.033335367839, -117.033335367839, -117.033335367839, 
    -117.083333333333, -122.291333516439, -122.291333516439, 
    -122.291333516439, -122.291333516439, -122.291333516439, 
    -122.291333516439, -122.291333516439, -122.291333516439, 
    -122.291333516439, -122.291333516439, -122.291333516439, 
    -122.291333516439, -122.291333516439, -122.291333516439, 
    -122.291333516439, -122.291333516439, -122.291333516439, 
    -122.291333516439, -122.291333516439, -122.291333516439, 
    -122.291333516439, -122.291333516439, -122.291333516439, 
    -122.291333516439, -122.291333516439, -122.291333516439, 
    -122.291333516439, -122.291333516439, -122.291333516439, 
    -122.291333516439, -122.291333516439, -122.291333516439, 
    -122.291333516439, -122.291333516439, -122.291333516439, 
    -122.291333516439, -122.291333516439, -122.291333516439, 
    -122.291333516439, -122.291333516439, -122.291333516439, 
    -122.291333516439, -122.291333516439, -122.291333516439, 
    -122.291333516439, -122.291333516439, -132.340337117513, 
    -132.340337117513, -132.340337117513, -132.340337117513, 
    -132.340337117513, -132.340337117513, -132.340337117513, 
    -132.340337117513, -132.340337117513, -132.340337117513, 
    -132.340337117513, -132.340337117513, -132.340337117513, 
    -132.340337117513, -132.340337117513, -132.340337117513, 
    -132.340337117513, -132.340337117513, -132.340337117513, 
    -132.340337117513, -132.340337117513, -132.340337117513, 
    -132.340337117513, -132.340337117513, -132.340337117513, 
    -132.340337117513, -132.340337117513, -132.340337117513, 
    -132.340337117513, -132.340337117513, -132.340337117513, 
    -132.340337117513, -132.340337117513, -132.340337117513, 
    -132.340337117513, -132.340337117513, -132.340337117513, 
    -132.340337117513, -132.340337117513, -132.340337117513, 
    -132.340337117513, -132.340337117513, -132.340337117513, 
    -132.340337117513, -132.340337117513, -132.340337117513, 
    -125.530331929525, -125.530331929525, -125.530331929525, 
    -125.530331929525, -125.530331929525, -125.530331929525, 
    -125.530331929525, -125.530331929525, -125.530331929525, 
    -125.530331929525, -125.530331929525, -125.530331929525, 
    -125.530331929525, -125.530331929525, -125.530331929525, 
    -125.530331929525, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.983334859212, -126.022223578559, 
    -125.983334859212, -125.933335622152, -125.958333333333, 
    -125.883336385091, -125.961906069801, -125.983334859212, 
    -126.083333333333, -126.047619047619, -126.003334554036, 
    -125.996971361565, -125.983334859212, -125.987879897609, 
    -126.003334554036, -125.996971361565, -125.983334859212, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.678786769058, -125.644443088108, -125.683331807454, 
    -125.71333211263, -125.61666615804, -125.673331197103, -125.833333333333, 
    -125.833333333333, -125.745831807454, -125.783330281576, 
    -125.716664632161, -125.66333211263, -125.683331807454, 
    -125.683331807454, -125.799997965495, -125.653331502279, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.40833791097, 
    -125.433339436849, -125.350001017253, -125.299997965495, -125.3047601609, 
    -125.358334859212, -125.40000406901, -125.233327229818, 
    -125.333333333333, -125.433339436849, -125.283330281576, 
    -125.333333333333, -125.299997965495, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.978789820816, -124.988889906141, 
    -124.973334248861, -124.833333333333, -125.013335164388, 
    -125.033335367839, -125.058335622152, -125.133336385091, 
    -125.083333333333, -124.983334859212, -124.983334859212, 
    -124.966668023003, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.683331807454, -124.683331807454, -124.683331807454, 
    -124.683331807454, -124.683331807454, -124.683331807454, 
    -124.683331807454, -124.683331807454, -124.683331807454, 
    -124.683331807454, -124.683331807454, -124.683331807454, 
    -124.753331502279, -124.733332951864, -124.666664971246, 
    -124.683331807454, -124.783330281576, -124.708331425985, 
    -124.696968309807, -124.683331807454, -124.683331807454, 
    -124.683331807454, -124.683331807454, -124.696968309807, 
    -124.745831807454, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.37333577474, 
    -124.383336385091, -124.383336385091, -124.433339436849, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -123.983334859212, 
    -123.983334859212, -123.983334859212, -123.983334859212, 
    -123.983334859212, -123.983334859212, -123.983334859212, 
    -123.996971361565, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.683331807454, -123.683331807454, -123.683331807454, 
    -123.683331807454, -123.683331807454, -123.683331807454, 
    -123.683331807454, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -122.983334859212, -122.983334859212, 
    -122.983334859212, -122.983334859212, -123.013335164388, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.683331807454, 
    -122.683331807454, -122.696968309807, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.345834096273, -122.345834096273, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.045834859212, -121.633331298828, 
    -121.633331298828, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.633331298828, -121.673329671224, 
    -121.333333333333, -121.333333333333, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.333333333333, 
    -121.033335367839, -121.033335367839, -121.033335367839, 
    -121.033335367839, -121.033335367839, -121.033335367839, 
    -121.033335367839, -121.033335367839, -121.033335367839, 
    -121.033335367839, -121.033335367839, -121.033335367839, 
    -121.083333333333, -121.083333333333, -120.633331298828, 
    -120.633331298828, -120.633331298828, -120.633331298828, 
    -120.633331298828, -120.633331298828, -120.633331298828, 
    -120.633331298828, -120.633331298828, -120.633331298828, 
    -120.645831425985, -120.633331298828, -120.333333333333, 
    -120.333333333333, -120.333333333333, -120.333333333333, 
    -120.333333333333, -120.333333333333, -120.333333333333, 
    -120.333333333333, -120.333333333333, -120.333333333333, 
    -120.320832570394, -120.333333333333, -120.033335367839, 
    -120.033335367839, -120.033335367839, -120.033335367839, 
    -120.033335367839, -120.033335367839, -120.033335367839, 
    -120.033335367839, -120.033335367839, -120.033335367839, 
    -120.033335367839, -120.033335367839, -119.633331298828, 
    -119.633331298828, -119.633331298828, -119.633331298828, 
    -119.633331298828, -119.633331298828, -119.633331298828, 
    -119.633331298828, -119.633331298828, -119.633331298828, 
    -119.633331298828, -119.333333333333, -119.333333333333, 
    -119.333333333333, -119.333333333333, -119.333333333333, 
    -119.333333333333, -119.333333333333, -119.333333333333, 
    -119.333333333333, -119.333333333333, -119.333333333333, 
    -119.033335367839, -119.033335367839, -119.033335367839, 
    -119.033335367839, -119.033335367839, -119.033335367839, 
    -119.033335367839, -119.033335367839, -119.033335367839, 
    -119.033335367839, -119.033335367839, -118.633331298828, 
    -118.633331298828, -118.633331298828, -118.633331298828, 
    -118.633331298828, -118.633331298828, -118.633331298828, 
    -118.633331298828, -118.620831807454, -118.633331298828, 
    -118.333333333333, -118.333333333333, -118.333333333333, 
    -118.333333333333, -118.333333333333, -118.333333333333, 
    -118.333333333333, -118.333333333333, -118.333333333333, 
    -118.033335367839, -118.033335367839, -118.033335367839, 
    -118.033335367839, -118.033335367839, -118.033335367839, 
    -118.033335367839, -118.033335367839, -118.045834859212, 
    -117.633331298828, -117.633331298828, -117.633331298828, 
    -117.633331298828, -117.633331298828, -117.633331298828, 
    -117.661903018043, -117.693330891927, -117.333333333333, 
    -117.333333333333, -117.333333333333, -117.333333333333, 
    -117.333333333333, -117.033335367839, -117.033335367839, 
    -117.033335367839, -117.083333333333, -125.134335835775, 
    -125.134335835775, -125.134335835775, -125.134335835775, 
    -125.134335835775, -125.134335835775, -125.134335835775, 
    -125.134335835775, -125.134335835775, -125.134335835775, 
    -125.134335835775, -125.134335835775, -125.134335835775, 
    -125.072331746419, -125.072331746419, -125.072331746419, 
    -125.072331746419, -125.072331746419, -125.072331746419, 
    -125.072331746419, -125.072331746419, -125.072331746419, 
    -125.072331746419, -125.072331746419, -125.072331746419, 
    -125.072331746419, -125.072331746419, -117.636334737142, 
    -117.636334737142, -117.636334737142, -117.636334737142, 
    -117.636334737142, -117.636334737142, -117.636334737142, 
    -117.636334737142, -117.636334737142, -117.636334737142, 
    -117.636334737142, -117.636334737142, -117.636334737142, 
    -117.636334737142, -117.748334248861, -117.748334248861, 
    -117.748334248861, -117.748334248861, -117.748334248861, 
    -117.748334248861, -117.748334248861, -117.748334248861, 
    -117.748334248861, -117.748334248861, -117.748334248861, 
    -117.748334248861, -117.748334248861, -117.748334248861, 
    -117.748334248861, -117.748334248861, -117.748334248861, 
    -117.748334248861, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.987879897609, -125.983334859212, 
    -125.987879897609, -125.983334859212, -125.996971361565, 
    -125.983334859212, -125.987879897609, -126.019048055013, 
    -125.983334859212, -125.833333333333, -126.083333333333, 
    -126.013335164388, -126.033334096273, -126.022223578559, 
    -125.987879897609, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.696968309807, -125.683331807454, -125.683331807454, 
    -125.678786769058, -125.733333333333, -125.733331589472, 
    -125.695832570394, -125.766662597656, -125.677776760525, 
    -125.783330281576, -125.733331044515, -125.683331807454, 
    -125.658330281576, -125.673332722982, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.683331807454, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.345834096273, -125.333333333333, 
    -125.361906505766, -125.37333577474, -125.433339436849, 
    -125.433339436849, -125.333333333333, -125.299997965495, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.345834096273, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.96969835686, -124.996971361565, -124.970834096273, 
    -124.973334248861, -124.833333333333, -125.133336385091, 
    -124.983334859212, -124.963335164388, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.683331807454, -124.683331807454, 
    -124.683331807454, -124.683331807454, -124.683331807454, 
    -124.683331807454, -124.683331807454, -124.683331807454, 
    -124.683331807454, -124.683331807454, -124.683331807454, 
    -124.704760596866, -124.753331502279, -124.766665140788, 
    -124.833333333333, -124.708331425985, -124.696968309807, 
    -124.683331807454, -124.683331807454, -124.683331807454, 
    -124.683331807454, -124.696968309807, -124.745831807454, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.37333577474, -124.383336385091, 
    -124.383336385091, -124.433339436849, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -123.983334859212, -123.983334859212, 
    -123.983334859212, -123.983334859212, -123.983334859212, 
    -123.983334859212, -123.983334859212, -123.996971361565, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.683331807454, 
    -123.683331807454, -123.683331807454, -123.683331807454, 
    -123.683331807454, -123.683331807454, -123.683331807454, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -122.983334859212, -122.983334859212, -122.983334859212, 
    -122.983334859212, -123.033335367839, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.683331807454, -122.683331807454, 
    -122.696968309807, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.345834096273, -122.345834096273, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.045834859212, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.673329671224, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.033335367839, 
    -121.033335367839, -121.033335367839, -121.033335367839, 
    -121.033335367839, -121.033335367839, -121.033335367839, 
    -121.033335367839, -121.033335367839, -121.033335367839, 
    -121.033335367839, -121.033335367839, -121.083333333333, 
    -121.083333333333, -120.633331298828, -120.633331298828, 
    -120.633331298828, -120.633331298828, -120.633331298828, 
    -120.633331298828, -120.633331298828, -120.633331298828, 
    -120.633331298828, -120.633331298828, -120.645831425985, 
    -120.633331298828, -120.333333333333, -120.333333333333, 
    -120.333333333333, -120.333333333333, -120.333333333333, 
    -120.333333333333, -120.333333333333, -120.333333333333, 
    -120.333333333333, -120.333333333333, -120.320832570394, 
    -120.333333333333, -120.033335367839, -120.033335367839, 
    -120.033335367839, -120.033335367839, -120.033335367839, 
    -120.033335367839, -120.033335367839, -120.033335367839, 
    -120.033335367839, -120.033335367839, -120.033335367839, 
    -120.033335367839, -119.633331298828, -119.633331298828, 
    -119.633331298828, -119.633331298828, -119.633331298828, 
    -119.633331298828, -119.633331298828, -119.633331298828, 
    -119.633331298828, -119.633331298828, -119.633331298828, 
    -119.333333333333, -119.333333333333, -119.333333333333, 
    -119.333333333333, -119.333333333333, -119.333333333333, 
    -119.333333333333, -119.333333333333, -119.333333333333, 
    -119.333333333333, -119.333333333333, -119.033335367839, 
    -119.033335367839, -119.033335367839, -119.033335367839, 
    -119.033335367839, -119.033335367839, -119.033335367839, 
    -119.033335367839, -119.033335367839, -119.033335367839, 
    -119.033335367839, -118.633331298828, -118.633331298828, 
    -118.633331298828, -118.633331298828, -118.633331298828, 
    -118.633331298828, -118.633331298828, -118.633331298828, 
    -118.620831807454, -118.633331298828, -118.333333333333, 
    -118.333333333333, -118.333333333333, -118.333333333333, 
    -118.333333333333, -118.333333333333, -118.333333333333, 
    -118.333333333333, -118.333333333333, -118.033335367839, 
    -118.033335367839, -118.033335367839, -118.033335367839, 
    -118.033335367839, -118.033335367839, -118.033335367839, 
    -118.033335367839, -118.045834859212, -117.633331298828, 
    -117.633331298828, -117.633331298828, -117.633331298828, 
    -117.633331298828, -117.633331298828, -117.661903018043, 
    -117.693330891927, -117.333333333333, -117.333333333333, 
    -117.333333333333, -117.333333333333, -117.333333333333, 
    -117.033335367839, -117.033335367839, -117.033335367839, 
    -117.083333333333, -118.208333333333, -118.208333333333, 
    -118.208333333333, -118.208333333333, -118.208333333333, 
    -118.208333333333, -118.208333333333, -118.208333333333, 
    -118.208333333333, -118.208333333333, -118.208333333333, 
    -118.208333333333, -118.208333333333, -118.208333333333, 
    -118.208333333333, -118.208333333333, -118.208333333333, 
    -118.208333333333, -118.885335286458, -118.885335286458, 
    -118.885335286458, -118.885335286458, -118.885335286458, 
    -118.885335286458, -118.885335286458, -118.885335286458, 
    -118.885335286458, -118.885335286458, -118.885335286458, 
    -118.885335286458, -118.885335286458, -118.885335286458, 
    -118.885335286458, -118.885335286458, -118.885335286458, 
    -118.885335286458, -118.885335286458, -118.885335286458, 
    -118.885335286458, -118.885335286458, -118.885335286458, 
    -118.885335286458, -118.885335286458, -118.885335286458, 
    -118.885335286458, -118.885335286458, -118.885335286458, 
    -118.885335286458, -133.333333333356, -133.000000000023, 
    -133.333333333356, -132.666666666689, -133.000000000023, 
    -132.333333333356, -132.666666666689, -132.000000000023, 
    -132.333333333356, -133.333333333356, -131.66666666669, 
    -132.000000000023, -133.000000000023, -131.333333333356, 
    -133.333333333356, -131.66666666669, -132.666666666689, 
    -131.000000000023, -133.000000000023, -131.333333333356, 
    -132.333333333356, -133.333333333356, -130.66666666669, 
    -132.666666666689, -131.000000000023, -132.000000000023, 
    -133.000000000023, -130.333333333356, -132.333333333356, 
    -133.333333333356, -130.66666666669, -131.66666666669, -132.666666666689, 
    -130.000000000023, -132.000000000023, -133.000000000023, 
    -130.333333333356, -131.333333333356, -132.333333333356, 
    -129.66666666669, -133.333333333356, -131.66666666669, -132.666666666689, 
    -130.000000000023, -131.000000000023, -132.000000000023, 
    -129.333333333356, -133.000000000023, -131.333333333356, 
    -132.333333333356, -129.66666666669, -133.333333333356, -130.66666666669, 
    -131.66666666669, -129.000000000023, -132.666666666689, 
    -131.000000000023, -132.000000000023, -129.333333333356, 
    -133.000000000023, -130.333333333356, -131.333333333356, 
    -128.66666666669, -132.333333333356, -133.333333333356, -130.66666666669, 
    -131.66666666669, -129.000000000023, -132.666666666689, 
    -130.000000000023, -131.000000000023, -128.333333333357, 
    -132.000000000023, -133.000000000023, -130.333333333356, 
    -131.333333333356, -128.66666666669, -132.333333333356, -129.66666666669, 
    -133.333333333356, -130.66666666669, -128.000000000023, -131.66666666669, 
    -132.666666666689, -130.000000000023, -131.000000000023, 
    -128.333333333357, -132.000000000023, -129.333333333356, 
    -133.000000000023, -130.333333333356, -127.66666666669, 
    -131.333333333356, -132.333333333356, -129.66666666669, 
    -133.333333333356, -130.66666666669, -128.000000000023, -131.66666666669, 
    -129.000000000023, -132.666666666689, -130.000000000023, 
    -127.333333333357, -131.000000000023, -132.000000000023, 
    -129.333333333356, -133.000000000023, -130.333333333356, 
    -127.66666666669, -131.333333333356, -128.66666666669, -132.333333333356, 
    -129.66666666669, -127.000000000023, -133.333333333356, -130.66666666669, 
    -131.66666666669, -129.000000000023, -132.666666666689, 
    -130.000000000023, -127.333333333357, -131.000000000023, 
    -128.333333333357, -132.000000000023, -129.333333333356, 
    -126.66666666669, -133.000000000023, -130.333333333356, 
    -131.333333333356, -128.66666666669, -132.333333333356, -129.66666666669, 
    -127.000000000023, -133.333333333356, -130.66666666669, 
    -128.000000000023, -131.66666666669, -129.000000000023, 
    -126.333333333357, -132.666666666689, -130.000000000023, 
    -131.000000000023, -128.333333333357, -132.000000000023, 
    -129.333333333356, -126.66666666669, -133.000000000023, 
    -130.333333333356, -127.66666666669, -131.333333333356, -128.66666666669, 
    -126.000000000023, -132.333333333356, -129.66666666669, 
    -133.333333333356, -130.66666666669, -128.000000000023, -131.66666666669, 
    -129.000000000023, -126.333333333357, -132.666666666689, 
    -130.000000000023, -127.333333333357, -131.000000000023, 
    -128.333333333357, -125.66666666669, -132.000000000023, 
    -129.333333333356, -133.000000000023, -130.333333333356, 
    -127.66666666669, -131.333333333356, -128.66666666669, -126.000000000023, 
    -132.333333333356, -129.66666666669, -127.000000000023, 
    -133.333333333356, -130.66666666669, -128.000000000023, 
    -125.333333333357, -131.66666666669, -129.000000000023, 
    -132.666666666689, -130.000000000023, -127.333333333357, 
    -131.000000000023, -128.333333333357, -125.66666666669, 
    -132.000000000023, -129.333333333356, -126.66666666669, 
    -133.000000000023, -130.333333333356, -127.66666666669, 
    -125.000000000024, -131.333333333356, -128.66666666669, 
    -132.333333333356, -129.66666666669, -127.000000000023, 
    -133.333333333356, -130.66666666669, -128.000000000023, 
    -125.333333333357, -131.66666666669, -129.000000000023, 
    -126.333333333357, -132.666666666689, -130.000000000023, 
    -127.333333333357, -124.66666666669, -131.000000000023, 
    -128.333333333357, -132.000000000023, -129.333333333356, 
    -126.66666666669, -133.000000000023, -130.333333333356, -127.66666666669, 
    -125.000000000024, -131.333333333356, -128.66666666669, 
    -126.000000000023, -132.333333333356, -129.66666666669, 
    -127.000000000023, -133.333333333356, -124.333333333357, 
    -130.66666666669, -128.000000000023, -131.66666666669, -129.000000000023, 
    -126.333333333357, -132.666666666689, -130.000000000023, 
    -127.333333333357, -124.66666666669, -131.000000000023, 
    -128.333333333357, -125.66666666669, -132.000000000023, 
    -129.333333333356, -126.66666666669, -133.000000000023, 
    -124.000000000024, -130.333333333356, -127.66666666669, 
    -131.333333333356, -128.66666666669, -126.000000000023, 
    -132.333333333356, -129.66666666669, -127.000000000023, 
    -133.333333333356, -124.333333333357, -130.66666666669, 
    -128.000000000023, -125.333333333357, -131.66666666669, 
    -129.000000000023, -126.333333333357, -132.666666666689, 
    -123.66666666669, -130.000000000023, -127.333333333357, 
    -131.000000000023, -128.333333333357, -125.66666666669, 
    -132.000000000023, -129.333333333356, -126.66666666669, 
    -133.000000000023, -124.000000000024, -130.333333333356, 
    -127.66666666669, -125.000000000024, -131.333333333356, -128.66666666669, 
    -126.000000000023, -132.333333333356, -123.333333333357, 
    -129.66666666669, -127.000000000023, -133.333333333356, -130.66666666669, 
    -128.000000000023, -125.333333333357, -131.66666666669, 
    -129.000000000023, -126.333333333357, -132.666666666689, 
    -123.66666666669, -130.000000000023, -127.333333333357, -124.66666666669, 
    -131.000000000023, -128.333333333357, -125.66666666669, 
    -132.000000000023, -123.000000000024, -129.333333333356, 
    -126.66666666669, -133.000000000023, -130.333333333356, -127.66666666669, 
    -125.000000000024, -131.333333333356, -128.66666666669, 
    -126.000000000023, -132.333333333356, -123.333333333357, 
    -129.66666666669, -127.000000000023, -133.333333333356, 
    -124.333333333357, -130.66666666669, -128.000000000023, 
    -125.333333333357, -131.66666666669, -122.66666666669, -129.000000000023, 
    -126.333333333357, -132.666666666689, -130.000000000023, 
    -127.333333333357, -124.66666666669, -131.000000000023, 
    -128.333333333357, -125.66666666669, -132.000000000023, 
    -123.000000000024, -129.333333333356, -126.66666666669, 
    -133.000000000023, -124.000000000024, -130.333333333356, 
    -127.66666666669, -125.000000000024, -131.333333333356, 
    -122.333333333357, -128.66666666669, -126.000000000023, 
    -132.333333333356, -129.66666666669, -127.000000000023, 
    -133.333333333356, -124.333333333357, -130.66666666669, 
    -128.000000000023, -125.333333333357, -131.66666666669, -122.66666666669, 
    -129.000000000023, -126.333333333357, -132.666666666689, 
    -123.66666666669, -130.000000000023, -127.333333333357, -124.66666666669, 
    -131.000000000023, -122.000000000024, -128.333333333357, 
    -125.66666666669, -132.000000000023, -129.333333333356, -126.66666666669, 
    -133.000000000023, -124.000000000024, -130.333333333356, 
    -127.66666666669, -125.000000000024, -131.333333333356, 
    -122.333333333357, -128.66666666669, -126.000000000023, 
    -132.333333333356, -123.333333333357, -129.66666666669, 
    -127.000000000023, -133.333333333356, -124.333333333357, 
    -130.66666666669, -121.666666666691, -128.000000000023, 
    -125.333333333357, -131.66666666669, -129.000000000023, 
    -126.333333333357, -132.666666666689, -123.66666666669, 
    -130.000000000023, -127.333333333357, -124.66666666669, 
    -131.000000000023, -122.000000000024, -128.333333333357, 
    -125.66666666669, -132.000000000023, -123.000000000024, 
    -129.333333333356, -126.66666666669, -133.000000000023, 
    -124.000000000024, -130.333333333356, -121.333333333357, 
    -127.66666666669, -125.000000000024, -131.333333333356, -128.66666666669, 
    -126.000000000023, -132.333333333356, -123.333333333357, 
    -129.66666666669, -127.000000000023, -133.333333333356, 
    -124.333333333357, -130.66666666669, -121.666666666691, 
    -128.000000000023, -125.333333333357, -131.66666666669, -122.66666666669, 
    -129.000000000023, -126.333333333357, -132.666666666689, 
    -123.66666666669, -130.000000000023, -121.000000000024, 
    -127.333333333357, -124.66666666669, -131.000000000023, 
    -128.333333333357, -125.66666666669, -132.000000000023, 
    -123.000000000024, -129.333333333356, -126.66666666669, 
    -133.000000000023, -124.000000000024, -130.333333333356, 
    -121.333333333357, -127.66666666669, -125.000000000024, 
    -131.333333333356, -122.333333333357, -128.66666666669, 
    -126.000000000023, -132.333333333356, -123.333333333357, 
    -129.66666666669, -120.666666666691, -127.000000000023, 
    -133.333333333356, -124.333333333357, -130.66666666669, 
    -128.000000000023, -125.333333333357, -131.66666666669, -122.66666666669, 
    -129.000000000023, -126.333333333357, -132.666666666689, 
    -123.66666666669, -130.000000000023, -121.000000000024, 
    -127.333333333357, -124.66666666669, -131.000000000023, 
    -122.000000000024, -128.333333333357, -125.66666666669, 
    -132.000000000023, -123.000000000024, -129.333333333356, 
    -120.333333333357, -126.66666666669, -133.000000000023, 
    -124.000000000024, -130.333333333356, -127.66666666669, 
    -125.000000000024, -131.333333333356, -122.333333333357, 
    -128.66666666669, -126.000000000023, -132.333333333356, 
    -123.333333333357, -129.66666666669, -120.666666666691, 
    -127.000000000023, -133.333333333356, -124.333333333357, 
    -130.66666666669, -121.666666666691, -128.000000000023, 
    -125.333333333357, -131.666666666689, -122.66666666669, 
    -129.000000000023, -120.000000000024, -126.333333333357, 
    -132.666666666689, -123.66666666669, -130.000000000023, 
    -127.333333333357, -124.66666666669, -131.000000000023, 
    -122.000000000024, -128.333333333357, -125.66666666669, 
    -132.000000000023, -123.000000000024, -129.333333333356, 
    -120.333333333357, -126.66666666669, -133.000000000023, 
    -124.000000000024, -130.333333333356, -121.333333333357, 
    -127.66666666669, -125.000000000024, -131.333333333356, 
    -122.333333333357, -128.66666666669, -119.666666666691, 
    -126.000000000023, -132.333333333356, -123.333333333357, 
    -129.66666666669, -127.000000000023, -133.333333333356, 
    -124.333333333357, -130.66666666669, -121.666666666691, 
    -128.000000000023, -125.333333333357, -131.66666666669, -122.66666666669, 
    -129.000000000023, -120.000000000024, -126.333333333357, 
    -132.666666666689, -123.66666666669, -130.000000000023, 
    -121.000000000024, -127.333333333357, -124.66666666669, 
    -131.000000000023, -122.000000000024, -128.333333333357, 
    -119.333333333357, -125.66666666669, -132.000000000023, 
    -123.000000000024, -129.333333333356, -126.66666666669, 
    -133.000000000023, -124.000000000024, -130.333333333356, 
    -121.333333333357, -127.66666666669, -125.000000000024, 
    -131.333333333356, -122.333333333357, -128.66666666669, 
    -119.666666666691, -126.000000000023, -132.333333333356, 
    -123.333333333357, -129.66666666669, -120.666666666691, 
    -127.000000000023, -133.333333333356, -124.333333333357, 
    -130.66666666669, -121.666666666691, -128.000000000023, 
    -119.000000000024, -125.333333333357, -131.666666666689, 
    -122.66666666669, -129.000000000023, -126.333333333357, 
    -132.666666666689, -123.66666666669, -130.000000000023, 
    -121.000000000024, -127.333333333357, -124.66666666669, 
    -131.000000000023, -122.000000000024, -128.333333333357, 
    -119.333333333357, -125.66666666669, -132.000000000023, 
    -123.000000000024, -129.333333333356, -120.333333333357, 
    -126.66666666669, -133.000000000023, -124.000000000024, 
    -130.333333333356, -121.333333333357, -127.66666666669, 
    -118.666666666691, -125.000000000024, -131.333333333356, 
    -122.333333333357, -128.66666666669, -126.000000000023, 
    -132.333333333356, -123.333333333357, -129.66666666669, 
    -120.666666666691, -127.000000000023, -133.333333333356, 
    -124.333333333357, -130.66666666669, -121.666666666691, 
    -128.000000000023, -119.000000000024, -125.333333333357, 
    -131.66666666669, -122.66666666669, -129.000000000023, -120.000000000024, 
    -126.333333333357, -132.666666666689, -123.66666666669, 
    -130.000000000023, -121.000000000024, -127.333333333357, 
    -118.333333333358, -124.66666666669, -131.000000000023, 
    -122.000000000024, -128.333333333357, -125.66666666669, 
    -132.000000000023, -123.000000000024, -129.333333333356, 
    -120.333333333357, -126.66666666669, -133.000000000023, 
    -124.000000000024, -130.333333333356, -121.333333333357, 
    -127.66666666669, -118.666666666691, -125.000000000024, 
    -131.333333333356, -122.333333333357, -128.66666666669, 
    -119.666666666691, -126.000000000023, -132.333333333356, 
    -123.333333333357, -129.66666666669, -120.666666666691, 
    -127.000000000023, -133.333333333356, -118.000000000024, 
    -124.333333333357, -130.66666666669, -121.666666666691, 
    -128.000000000023, -125.333333333357, -131.66666666669, -122.66666666669, 
    -129.000000000023, -120.000000000024, -126.333333333357, 
    -132.666666666689, -123.66666666669, -130.000000000023, 
    -121.000000000024, -127.333333333357, -118.333333333358, 
    -124.66666666669, -131.000000000023, -122.000000000024, 
    -128.333333333357, -119.333333333357, -125.66666666669, 
    -132.000000000023, -123.000000000024, -129.333333333356, 
    -120.333333333357, -126.66666666669, -133.000000000023, 
    -117.666666666691, -124.000000000024, -130.333333333356, 
    -121.333333333357, -127.66666666669, -125.000000000024, 
    -131.333333333356, -122.333333333357, -128.66666666669, 
    -119.666666666691, -126.000000000023, -132.333333333356, 
    -123.333333333357, -129.66666666669, -120.666666666691, 
    -127.000000000023, -133.333333333356, -118.000000000024, 
    -124.333333333357, -130.66666666669, -121.666666666691, 
    -128.000000000023, -119.000000000024, -125.333333333357, 
    -131.66666666669, -122.66666666669, -129.000000000023, -120.000000000024, 
    -126.333333333357, -132.666666666689, -117.333333333358, 
    -123.66666666669, -130.000000000023, -121.000000000024, 
    -127.333333333357, -124.66666666669, -131.000000000023, 
    -122.000000000024, -128.333333333357, -119.333333333357, 
    -125.66666666669, -132.000000000023, -123.000000000024, 
    -129.333333333356, -120.333333333357, -126.66666666669, 
    -133.000000000023, -117.666666666691, -124.000000000024, 
    -130.333333333356, -121.333333333357, -127.66666666669, 
    -118.666666666691, -125.000000000024, -131.333333333356, 
    -122.333333333357, -128.66666666669, -119.666666666691, 
    -126.000000000023, -132.333333333356, -117.000000000024, 
    -123.333333333357, -129.66666666669, -120.666666666691, 
    -127.000000000023, -133.333333333356, -124.333333333357, 
    -130.66666666669, -121.666666666691, -128.000000000023, 
    -119.000000000024, -125.333333333357, -131.66666666669, -122.66666666669, 
    -129.000000000023, -120.000000000024, -126.333333333357, 
    -132.666666666689, -117.333333333358, -123.66666666669, 
    -130.000000000023, -121.000000000024, -127.333333333357, 
    -118.333333333358, -124.66666666669, -131.000000000023, 
    -122.000000000024, -128.333333333357, -119.333333333357, 
    -125.66666666669, -132.000000000023, -123.000000000024, 
    -129.333333333356, -120.333333333357, -126.66666666669, 
    -133.000000000023, -124.000000000024, -130.333333333356, 
    -121.333333333357, -127.66666666669, -118.666666666691, 
    -125.000000000024, -131.333333333356, -122.333333333357, 
    -128.66666666669, -119.666666666691, -126.000000000023, 
    -132.333333333356, -117.000000000024, -123.333333333357, 
    -129.66666666669, -120.666666666691, -127.000000000023, 
    -133.333333333356, -118.000000000024, -124.333333333357, 
    -130.66666666669, -121.666666666691, -128.000000000023, 
    -119.000000000024, -125.333333333357, -131.66666666669, -122.66666666669, 
    -129.000000000023, -120.000000000024, -126.333333333357, 
    -132.666666666689, -123.66666666669, -130.000000000023, 
    -121.000000000024, -127.333333333357, -118.333333333358, 
    -124.66666666669, -131.000000000023, -122.000000000024, 
    -128.333333333357, -119.333333333357, -125.66666666669, 
    -132.000000000023, -123.000000000024, -129.333333333356, 
    -120.333333333357, -126.66666666669, -133.000000000023, 
    -117.666666666691, -124.000000000024, -130.333333333356, 
    -121.333333333357, -127.66666666669, -118.666666666691, 
    -125.000000000024, -131.333333333356, -122.333333333357, 
    -128.66666666669, -119.666666666691, -126.000000000023, 
    -132.333333333356, -123.333333333357, -129.66666666669, 
    -120.666666666691, -127.000000000023, -133.333333333356, 
    -118.000000000024, -124.333333333357, -130.66666666669, 
    -121.666666666691, -128.000000000023, -119.000000000024, 
    -125.333333333357, -131.66666666669, -122.66666666669, -129.000000000023, 
    -120.000000000024, -126.333333333357, -132.666666666689, 
    -117.333333333358, -123.66666666669, -130.000000000023, 
    -121.000000000024, -127.333333333357, -118.333333333358, 
    -124.66666666669, -131.000000000023, -122.000000000024, 
    -128.333333333357, -119.333333333357, -125.66666666669, 
    -132.000000000023, -123.000000000024, -129.333333333356, 
    -120.333333333357, -126.66666666669, -133.000000000023, 
    -117.666666666691, -124.000000000024, -130.333333333356, 
    -121.333333333357, -127.66666666669, -118.666666666691, 
    -125.000000000024, -131.333333333356, -122.333333333357, 
    -128.66666666669, -119.666666666691, -126.000000000023, 
    -132.333333333356, -123.333333333357, -129.66666666669, 
    -120.666666666691, -127.000000000023, -133.333333333356, 
    -118.000000000024, -124.333333333357, -130.66666666669, 
    -121.666666666691, -128.000000000023, -119.000000000024, 
    -125.333333333357, -131.66666666669, -122.66666666669, -129.000000000023, 
    -120.000000000024, -126.333333333357, -132.666666666689, 
    -123.66666666669, -130.000000000023, -121.000000000024, 
    -127.333333333357, -124.66666666669, -131.000000000023, 
    -122.000000000024, -128.333333333357, -119.333333333357, 
    -125.66666666669, -132.000000000023, -123.000000000024, 
    -129.333333333356, -120.333333333357, -126.66666666669, 
    -133.000000000023, -117.666666666691, -124.000000000024, 
    -130.333333333356, -121.333333333357, -127.66666666669, 
    -118.666666666691, -125.000000000024, -131.333333333356, 
    -122.333333333357, -128.66666666669, -126.000000000023, 
    -132.333333333356, -123.333333333357, -129.66666666669, 
    -127.000000000023, -133.333333333356, -124.333333333357, 
    -130.66666666669, -121.666666666691, -128.000000000023, 
    -119.000000000024, -125.333333333357, -131.66666666669, -122.66666666669, 
    -129.000000000023, -120.000000000024, -126.333333333357, 
    -132.666666666689, -123.66666666669, -130.000000000023, 
    -121.000000000024, -127.333333333357, -124.66666666669, 
    -131.000000000023, -122.000000000024, -128.333333333357, 
    -125.66666666669, -132.000000000023, -123.000000000024, 
    -129.333333333356, -126.66666666669, -133.000000000023, 
    -124.000000000024, -130.333333333356, -121.333333333357, 
    -127.66666666669, -118.666666666691, -125.000000000024, 
    -131.333333333356, -122.333333333357, -128.66666666669, 
    -126.000000000023, -132.333333333356, -123.333333333357, 
    -129.66666666669, -127.000000000023, -133.333333333356, 
    -124.333333333357, -130.66666666669, -121.666666666691, 
    -128.000000000023, -125.333333333357, -131.66666666669, -122.66666666669, 
    -129.000000000023, -126.333333333357, -132.666666666689, 
    -123.66666666669, -130.000000000023, -127.333333333357, -124.66666666669, 
    -131.000000000023, -122.000000000024, -128.333333333357, 
    -125.66666666669, -132.000000000023, -123.000000000024, 
    -129.333333333356, -126.66666666669, -133.000000000023, 
    -124.000000000024, -130.333333333356, -127.66666666669, 
    -125.000000000024, -131.333333333356, -122.333333333357, 
    -128.66666666669, -126.000000000023, -132.333333333356, 
    -123.333333333357, -129.66666666669, -127.000000000023, 
    -133.333333333356, -124.333333333357, -130.66666666669, 
    -128.000000000023, -125.333333333357, -131.66666666669, -122.66666666669, 
    -129.000000000023, -126.333333333357, -132.666666666689, 
    -123.66666666669, -130.000000000023, -127.333333333357, -124.66666666669, 
    -131.000000000023, -128.333333333357, -125.66666666669, 
    -132.000000000023, -123.000000000024, -129.333333333356, 
    -126.66666666669, -133.000000000023, -124.000000000024, 
    -130.333333333356, -127.66666666669, -125.000000000024, 
    -131.333333333356, -122.333333333357, -128.66666666669, 
    -126.000000000023, -132.333333333356, -123.333333333357, 
    -129.66666666669, -127.000000000023, -133.333333333356, 
    -124.333333333357, -130.66666666669, -128.000000000023, 
    -125.333333333357, -131.66666666669, -122.66666666669, -129.000000000023, 
    -126.333333333357, -132.666666666689, -123.66666666669, 
    -130.000000000023, -127.333333333357, -124.66666666669, 
    -131.000000000023, -128.333333333357, -125.66666666669, 
    -132.000000000023, -123.000000000024, -129.333333333356, 
    -126.66666666669, -133.000000000023, -124.000000000024, 
    -130.333333333356, -127.66666666669, -125.000000000024, 
    -131.333333333356, -128.66666666669, -126.000000000023, 
    -132.333333333356, -123.333333333357, -129.66666666669, 
    -127.000000000023, -133.333333333356, -124.333333333357, 
    -130.66666666669, -128.000000000023, -125.333333333357, -131.66666666669, 
    -129.000000000023, -126.333333333357, -132.666666666689, 
    -123.66666666669, -130.000000000023, -127.333333333357, -124.66666666669, 
    -131.000000000023, -128.333333333357, -125.66666666669, 
    -132.000000000023, -123.000000000024, -129.333333333356, 
    -126.66666666669, -133.000000000023, -124.000000000024, 
    -130.333333333356, -127.66666666669, -125.000000000024, 
    -131.333333333356, -128.66666666669, -126.000000000023, 
    -132.333333333356, -129.66666666669, -127.000000000023, 
    -133.333333333356, -124.333333333357, -130.66666666669, 
    -128.000000000023, -125.333333333357, -131.66666666669, 
    -129.000000000023, -126.333333333357, -132.666666666689, 
    -130.000000000023, -127.333333333357, -124.66666666669, 
    -131.000000000023, -128.333333333357, -125.66666666669, 
    -132.000000000023, -129.333333333356, -126.66666666669, 
    -133.000000000023, -124.000000000024, -130.333333333356, 
    -127.66666666669, -125.000000000024, -131.333333333356, -128.66666666669, 
    -126.000000000023, -132.333333333356, -129.66666666669, 
    -127.000000000023, -133.333333333356, -124.333333333357, 
    -130.66666666669, -128.000000000023, -125.333333333357, -131.66666666669, 
    -129.000000000023, -126.333333333357, -132.666666666689, 
    -130.000000000023, -127.333333333357, -124.66666666669, 
    -131.000000000023, -128.333333333357, -125.66666666669, 
    -132.000000000023, -129.333333333356, -126.66666666669, 
    -133.000000000023, -130.333333333356, -127.66666666669, 
    -125.000000000024, -131.333333333356, -128.66666666669, 
    -126.000000000023, -132.333333333356, -129.66666666669, 
    -127.000000000023, -133.333333333356, -124.333333333357, 
    -130.66666666669, -128.000000000023, -125.333333333357, -131.66666666669, 
    -129.000000000023, -126.333333333357, -132.666666666689, 
    -130.000000000023, -127.333333333357, -124.66666666669, 
    -131.000000000023, -128.333333333357, -125.66666666669, 
    -132.000000000023, -129.333333333356, -126.66666666669, 
    -133.000000000023, -130.333333333356, -127.66666666669, 
    -125.000000000024, -131.333333333356, -128.66666666669, 
    -126.000000000023, -132.333333333356, -129.66666666669, 
    -127.000000000023, -133.333333333356, -124.333333333357, 
    -130.66666666669, -128.000000000023, -125.333333333357, -131.66666666669, 
    -129.000000000023, -126.333333333357, -132.666666666689, 
    -130.000000000023, -127.333333333357, -124.66666666669, 
    -131.000000000023, -128.333333333357, -125.66666666669, 
    -132.000000000023, -129.333333333356, -126.66666666669, 
    -133.000000000023, -130.333333333356, -127.66666666669, 
    -125.000000000024, -131.333333333356, -128.66666666669, 
    -126.000000000023, -132.333333333356, -129.66666666669, 
    -127.000000000023, -133.333333333356, -130.66666666669, 
    -128.000000000023, -125.333333333357, -131.66666666669, 
    -129.000000000023, -126.333333333357, -132.666666666689, 
    -130.000000000023, -127.333333333357, -131.000000000023, 
    -128.333333333357, -125.66666666669, -132.000000000023, 
    -129.333333333356, -126.66666666669, -133.000000000023, 
    -130.333333333356, -127.66666666669, -125.000000000024, 
    -131.333333333356, -128.66666666669, -126.000000000023, 
    -132.333333333356, -129.66666666669, -127.000000000023, 
    -133.333333333356, -130.66666666669, -128.000000000023, 
    -125.333333333357, -131.66666666669, -129.000000000023, 
    -126.333333333357, -132.666666666689, -130.000000000023, 
    -127.333333333357, -124.66666666669, -131.000000000023, 
    -128.333333333357, -125.66666666669, -132.000000000023, 
    -129.333333333356, -126.66666666669, -133.000000000023, 
    -130.333333333356, -127.66666666669, -125.000000000024, 
    -131.333333333356, -128.66666666669, -126.000000000023, 
    -132.333333333356, -129.66666666669, -127.000000000023, 
    -133.333333333356, -130.66666666669, -128.000000000023, 
    -125.333333333357, -131.66666666669, -129.000000000023, 
    -126.333333333357, -132.666666666689, -130.000000000023, 
    -127.333333333357, -124.66666666669, -131.000000000023, 
    -128.333333333357, -125.66666666669, -132.000000000023, 
    -129.333333333356, -126.66666666669, -133.000000000023, 
    -130.333333333356, -127.66666666669, -131.333333333356, -128.66666666669, 
    -126.000000000023, -132.333333333356, -129.66666666669, 
    -127.000000000023, -133.333333333356, -130.66666666669, 
    -128.000000000023, -125.333333333357, -131.66666666669, 
    -129.000000000023, -126.333333333357, -132.666666666689, 
    -130.000000000023, -127.333333333357, -131.000000000023, 
    -128.333333333357, -125.66666666669, -132.000000000023, 
    -129.333333333356, -126.66666666669, -133.000000000023, 
    -130.333333333356, -127.66666666669, -131.333333333356, -128.66666666669, 
    -126.000000000023, -132.333333333356, -129.66666666669, 
    -127.000000000023, -133.333333333356, -130.66666666669, 
    -128.000000000023, -125.333333333357, -131.66666666669, 
    -129.000000000023, -126.333333333357, -132.666666666689, 
    -130.000000000023, -127.333333333357, -131.000000000023, 
    -128.333333333357, -125.66666666669, -132.000000000023, 
    -129.333333333356, -126.66666666669, -133.000000000023, 
    -130.333333333356, -127.66666666669, -131.333333333356, -128.66666666669, 
    -126.000000000023, -132.333333333356, -129.66666666669, 
    -127.000000000023, -130.66666666669, -128.000000000023, 
    -125.333333333357, -131.66666666669, -129.000000000023, 
    -126.333333333357, -132.666666666689, -130.000000000023, 
    -127.333333333357, -131.000000000023, -128.333333333357, 
    -125.66666666669, -132.000000000023, -129.333333333356, -126.66666666669, 
    -130.333333333356, -127.66666666669, -125.000000000024, 
    -131.333333333356, -128.66666666669, -126.000000000023, 
    -132.333333333356, -129.66666666669, -127.000000000023, -130.66666666669, 
    -128.000000000023, -125.333333333357, -131.66666666669, 
    -129.000000000023, -126.333333333357, -130.000000000023, 
    -127.333333333357, -131.000000000023, -128.333333333357, 
    -125.66666666669, -132.000000000023, -129.333333333356, -126.66666666669, 
    -130.333333333356, -127.66666666669, -125.000000000024, 
    -131.333333333356, -128.66666666669, -126.000000000023, -129.66666666669, 
    -127.000000000023, -130.66666666669, -128.000000000023, 
    -125.333333333357, -131.66666666669, -129.000000000023, 
    -126.333333333357, -130.000000000023, -127.333333333357, 
    -131.000000000023, -128.333333333357, -125.66666666669, 
    -129.333333333356, -126.66666666669, -130.333333333356, -127.66666666669, 
    -125.000000000024, -131.333333333356, -128.66666666669, 
    -126.000000000023, -129.66666666669, -127.000000000023, -130.66666666669, 
    -128.000000000023, -125.333333333357, -129.000000000023, 
    -126.333333333357, -130.000000000023, -127.333333333357, 
    -131.000000000023, -128.333333333357, -125.66666666669, 
    -129.333333333356, -126.66666666669, -130.333333333356, -127.66666666669, 
    -125.000000000024, -128.66666666669, -126.000000000023, -129.66666666669, 
    -127.000000000023, -130.66666666669, -128.000000000023, 
    -125.333333333357, -129.000000000023, -126.333333333357, 
    -130.000000000023, -127.333333333357, -128.333333333357, 
    -125.66666666669, -129.333333333356, -126.66666666669, -130.333333333356, 
    -127.66666666669, -125.000000000024, -128.66666666669, -126.000000000023, 
    -129.66666666669, -127.000000000023, -128.000000000023, 
    -125.333333333357, -129.000000000023, -126.333333333357, 
    -130.000000000023, -127.333333333357, -124.66666666669, 
    -128.333333333357, -125.66666666669, -129.333333333356, -126.66666666669, 
    -127.66666666669, -125.000000000024, -128.66666666669, -126.000000000023, 
    -129.66666666669, -127.000000000023, -128.000000000023, 
    -125.333333333357, -129.000000000023, -126.333333333357, 
    -127.333333333357, -124.66666666669, -128.333333333357, -125.66666666669, 
    -129.333333333356, -126.66666666669, -127.66666666669, -125.000000000024, 
    -128.66666666669, -126.000000000023, -127.000000000023, 
    -128.000000000023, -125.333333333357, -129.000000000023, 
    -126.333333333357, -127.333333333357, -124.66666666669, 
    -128.333333333357, -125.66666666669, -126.66666666669, -127.66666666669, 
    -125.000000000024, -128.66666666669, -126.000000000023, 
    -127.000000000023, -128.000000000023, -125.333333333357, 
    -126.333333333357, -127.333333333357, -124.66666666669, 
    -128.333333333357, -125.66666666669, -126.66666666669, -127.66666666669, 
    -125.000000000024, -126.000000000023, -127.000000000023, 
    -128.000000000023, -125.333333333357, -126.333333333357, 
    -127.333333333357, -124.66666666669, -125.66666666669, -126.66666666669, 
    -127.66666666669, -125.000000000024, -126.000000000023, 
    -127.000000000023, -125.333333333357, -126.333333333357, 
    -127.333333333357, -124.66666666669, -125.66666666669, -126.66666666669, 
    -125.000000000024, -126.000000000023, -127.000000000023, 
    -124.333333333357, -125.333333333357, -126.333333333357, 
    -124.66666666669, -125.66666666669, -126.66666666669, -125.000000000024, 
    -126.000000000023, -124.333333333357, -125.333333333357, 
    -126.333333333357, -124.66666666669, -125.66666666669, -125.000000000024, 
    -126.000000000023, -124.333333333357, -125.333333333357, 
    -124.66666666669, -125.66666666669, -125.000000000024, -125.333333333357, 
    -124.66666666669, -125.000000000024, -124.333333333357, -124.66666666669 ;

 obs_lat = 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3666661580404, 38.6666666666667, 38.966667175293, 
    39.3666661580404, 39.6666666666667, 39.966667175293, 40.3666661580404, 
    40.6666666666667, 40.966667175293, 41.3666661580404, 41.6666666666667, 
    41.966667175293, 42.3666661580404, 42.6666666666667, 42.966667175293, 
    43.3666661580404, 43.6666666666667, 43.966667175293, 44.3666661580404, 
    44.6666666666667, 44.966667175293, 45.3666661580404, 45.6666666666667, 
    45.966667175293, 46.3666661580404, 46.6666666666667, 46.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.966667175293, 41.3666661580404, 41.6666666666667, 41.966667175293, 
    42.3666661580404, 42.6666666666667, 42.966667175293, 43.3666661580404, 
    43.6666666666667, 43.966667175293, 44.3666661580404, 44.6666666666667, 
    44.966667175293, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    39.966667175293, 40.3666661580404, 40.6666666666667, 40.966667175293, 
    41.3666661580404, 41.6666666666667, 41.966667175293, 42.3666661580404, 
    42.6666666666667, 42.966667175293, 43.3666661580404, 43.6666666666667, 
    43.966667175293, 44.3666661580404, 44.6666666666667, 44.966667175293, 
    45.3666661580404, 45.6666666666667, 45.966667175293, 46.3666661580404, 
    46.6666666666667, 46.966667175293, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 38.3666661580404, 38.6666666666667, 
    38.966667175293, 39.3666661580404, 39.6666666666667, 39.966667175293, 
    40.3666661580404, 40.6666666666667, 40.966667175293, 41.3666661580404, 
    41.6666666666667, 41.966667175293, 42.3666661580404, 42.6666666666667, 
    42.966667175293, 43.3666661580404, 43.6666666666667, 43.966667175293, 
    44.3666661580404, 44.6666666666667, 44.966667175293, 45.3666661580404, 
    45.6666666666667, 45.966667175293, 46.3666661580404, 46.6666666666667, 
    46.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3666661580404, 38.6666666666667, 38.966667175293, 
    39.3666661580404, 39.6666666666667, 39.966667175293, 40.3666661580404, 
    40.6666666666667, 40.966667175293, 41.3666661580404, 41.6666666666667, 
    41.966667175293, 42.3666661580404, 42.6666666666667, 42.966667175293, 
    43.3666661580404, 43.6666666666667, 43.966667175293, 44.3666661580404, 
    44.6666666666667, 44.966667175293, 45.3666661580404, 45.6666666666667, 
    45.966667175293, 46.3666661580404, 46.6666666666667, 46.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.966667175293, 41.3666661580404, 41.6666666666667, 41.966667175293, 
    42.3666661580404, 42.6666666666667, 42.966667175293, 43.3666661580404, 
    43.6666666666667, 43.966667175293, 44.3666661580404, 44.6666666666667, 
    44.966667175293, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    39.966667175293, 40.3666661580404, 40.6666666666667, 40.966667175293, 
    41.3666661580404, 41.6666666666667, 41.966667175293, 42.3666661580404, 
    42.6666666666667, 42.966667175293, 43.3666661580404, 43.6666666666667, 
    43.966667175293, 44.3666661580404, 44.6666666666667, 44.966667175293, 
    45.3666661580404, 45.6666666666667, 45.966667175293, 46.3666661580404, 
    46.6666666666667, 46.966667175293, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 38.3666661580404, 38.6666666666667, 
    38.966667175293, 39.3666661580404, 39.6666666666667, 39.966667175293, 
    40.3666661580404, 40.6666666666667, 40.966667175293, 41.3666661580404, 
    41.6666666666667, 41.966667175293, 42.3666661580404, 42.6666666666667, 
    42.966667175293, 43.3666661580404, 43.6666666666667, 43.966667175293, 
    44.3666661580404, 44.6666666666667, 44.966667175293, 45.3666661580404, 
    45.6666666666667, 45.966667175293, 46.3666661580404, 46.6666666666667, 
    46.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3666661580404, 38.6666666666667, 38.966667175293, 
    39.3666661580404, 39.6666666666667, 39.966667175293, 40.3666661580404, 
    40.6666666666667, 40.966667175293, 41.3666661580404, 41.6666666666667, 
    41.966667175293, 42.3666661580404, 42.6666666666667, 42.966667175293, 
    43.3666661580404, 43.6666666666667, 43.966667175293, 44.3666661580404, 
    44.6666666666667, 44.966667175293, 45.3666661580404, 45.6666666666667, 
    45.966667175293, 46.3666661580404, 46.6666666666667, 46.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.966667175293, 41.3666661580404, 41.6666666666667, 41.966667175293, 
    42.3666661580404, 42.6666666666667, 42.966667175293, 43.3666661580404, 
    43.6666666666667, 43.966667175293, 44.3666661580404, 44.6666666666667, 
    44.966667175293, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    39.966667175293, 40.3666661580404, 40.6666666666667, 40.966667175293, 
    41.3666661580404, 41.6666666666667, 41.966667175293, 42.3666661580404, 
    42.6666666666667, 42.966667175293, 43.3666661580404, 43.6666666666667, 
    43.966667175293, 44.3666661580404, 44.6666666666667, 44.966667175293, 
    45.3666661580404, 45.6666666666667, 45.966667175293, 46.3666661580404, 
    46.6666666666667, 46.966667175293, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 38.3666661580404, 38.6666666666667, 
    38.966667175293, 39.3666661580404, 39.6666666666667, 39.966667175293, 
    40.3666661580404, 40.6666666666667, 40.966667175293, 41.3666661580404, 
    41.6666666666667, 41.966667175293, 42.3666661580404, 42.6666666666667, 
    42.966667175293, 43.3666661580404, 43.6666666666667, 43.966667175293, 
    44.3666661580404, 44.6666666666667, 44.966667175293, 45.3666661580404, 
    45.6666666666667, 45.966667175293, 46.3666661580404, 46.6666666666667, 
    46.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3666661580404, 38.6666666666667, 38.966667175293, 
    39.3666661580404, 39.6666666666667, 39.966667175293, 40.3666661580404, 
    40.6666666666667, 40.966667175293, 41.3666661580404, 41.6666666666667, 
    41.966667175293, 42.3666661580404, 42.6666666666667, 42.966667175293, 
    43.3666661580404, 43.6666666666667, 43.966667175293, 44.3666661580404, 
    44.6666666666667, 44.966667175293, 45.3666661580404, 45.6666666666667, 
    45.966667175293, 46.3666661580404, 46.6666666666667, 46.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.966667175293, 41.3666661580404, 41.6757574370413, 41.966667175293, 
    42.3523802984328, 42.5666681925456, 42.9952385312035, 43.3666659037272, 
    43.6291672388713, 43.966667175293, 44.3666661580404, 44.6809521629697, 
    44.966667175293, 45.3566660563151, 45.6666666666667, 45.9666672908899, 
    46.3757571596088, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    39.966667175293, 40.3666661580404, 40.6666666666667, 40.966667175293, 
    41.3575752720688, 41.6666666666667, 41.966667175293, 42.3666659037272, 
    42.6380956740606, 42.9666670481364, 43.3999989827474, 43.6999994913737, 
    43.9541670481364, 44.7666651407878, 44.9666675385975, 45.3666659037272, 
    45.6666666666667, 45.966667175293, 46.3666664759318, 46.6666666666667, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.966667175293, 41.3666661580404, 41.6666666666667, 41.9333337148031, 
    42.3809518359956, 42.5916678110759, 43.0333340962728, 43.3166662851969, 
    43.6999994913737, 43.9166666666667, 44.2666651407878, 44.6866663614909, 
    45.0000012715658, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3791662851969, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    39.966667175293, 40.3888884650336, 40.6666666666667, 41.006667582194, 
    41.3575752720688, 41.6444447835286, 41.9952385312035, 42.3952378772554, 
    42.5666681925456, 43.3166662851969, 43.6416670481364, 44.6999994913737, 
    44.9666675991482, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    40.4266665140788, 40.6666666666667, 40.9757580612645, 41.3380948021298, 
    41.6380956740606, 43.3166662851969, 43.6666666666667, 44.7041660944621, 
    44.9757580612645, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.657575896292, 46.9541670481364, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 44.9866671244303, 
    45.3666661580404, 45.6666666666667, 46.3666661580404, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3575752720688, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3766661326091, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.657575896292, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.9541670481364, 36.3791662851969, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6541668574015, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3266657511393, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6166674296061, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6166674296061, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.9541670481364, 33.3166662851969, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.9541670481364, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3523802984329, 32.6466669718424, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 37.5846659342448, 
    37.5846659342448, 37.5846659342448, 37.5846659342448, 37.5846659342448, 
    37.5846659342448, 37.5846659342448, 37.5846659342448, 37.5846659342448, 
    37.5846659342448, 37.5846659342448, 37.5846659342448, 37.5846659342448, 
    37.5846659342448, 37.5846659342448, 37.5846659342448, 37.5846659342448, 
    37.5846659342448, 37.5846659342448, 37.5846659342448, 37.5846659342448, 
    37.5846659342448, 37.5846659342448, 37.5846659342448, 37.5846659342448, 
    37.5846659342448, 37.5846659342448, 37.5846659342448, 37.5846659342448, 
    37.5846659342448, 37.5846659342448, 37.5846659342448, 37.5846659342448, 
    37.5846659342448, 37.5846659342448, 37.5846659342448, 37.5846659342448, 
    37.5846659342448, 38.4526659647624, 38.4526659647624, 38.4526659647624, 
    38.4526659647624, 38.4526659647624, 38.4526659647624, 38.4526659647624, 
    38.4526659647624, 38.4526659647624, 38.4526659647624, 38.4526659647624, 
    38.4526659647624, 38.4526659647624, 38.4526659647624, 38.4526659647624, 
    38.4526659647624, 38.4526659647624, 38.4526659647624, 38.4526659647624, 
    38.4526659647624, 38.4526659647624, 38.4526659647624, 38.4526659647624, 
    38.4526659647624, 38.4526659647624, 38.4526659647624, 38.4526659647624, 
    38.4526659647624, 38.4526659647624, 38.4526659647624, 38.4526659647624, 
    38.4526659647624, 38.4526659647624, 38.4526659647624, 38.4526659647624, 
    38.4526659647624, 38.4526659647624, 38.4526659647624, 38.4526659647624, 
    38.4526659647624, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3666661580404, 38.6666666666667, 38.966667175293, 
    39.3666661580404, 39.6666666666667, 39.966667175293, 40.3666661580404, 
    40.6666666666667, 40.966667175293, 41.3666661580404, 41.6666666666667, 
    41.966667175293, 42.3666661580404, 42.6666666666667, 42.966667175293, 
    43.3666661580404, 43.6666666666667, 43.966667175293, 44.3666661580404, 
    44.6666666666667, 44.966667175293, 45.3666661580404, 45.6666666666667, 
    45.966667175293, 46.3666661580404, 46.6666666666667, 46.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.966667175293, 41.3666661580404, 41.6666666666667, 41.966667175293, 
    42.3666661580404, 42.6666666666667, 42.966667175293, 43.3666661580404, 
    43.6666666666667, 43.966667175293, 44.3666661580404, 44.6666666666667, 
    44.966667175293, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    39.966667175293, 40.3666661580404, 40.6666666666667, 40.966667175293, 
    41.3666661580404, 41.6666666666667, 41.966667175293, 42.3666661580404, 
    42.6666666666667, 42.966667175293, 43.3666661580404, 43.6666666666667, 
    43.966667175293, 44.3666661580404, 44.6666666666667, 44.966667175293, 
    45.3666661580404, 45.6666666666667, 45.966667175293, 46.3666661580404, 
    46.6666666666667, 46.966667175293, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 38.3666661580404, 38.6666666666667, 
    38.966667175293, 39.3666661580404, 39.6666666666667, 39.966667175293, 
    40.3666661580404, 40.6666666666667, 40.966667175293, 41.3666661580404, 
    41.6666666666667, 41.966667175293, 42.3666661580404, 42.6666666666667, 
    42.966667175293, 43.3666661580404, 43.6666666666667, 43.966667175293, 
    44.3666661580404, 44.6666666666667, 44.966667175293, 45.3666661580404, 
    45.6666666666667, 45.966667175293, 46.3666661580404, 46.6666666666667, 
    46.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3666661580404, 38.6666666666667, 38.966667175293, 
    39.3666661580404, 39.6666666666667, 39.966667175293, 40.3666661580404, 
    40.6666666666667, 40.966667175293, 41.3666661580404, 41.6666666666667, 
    41.966667175293, 42.3666661580404, 42.6666666666667, 42.966667175293, 
    43.3666661580404, 43.6666666666667, 43.966667175293, 44.3666661580404, 
    44.6666666666667, 44.966667175293, 45.3666661580404, 45.6666666666667, 
    45.966667175293, 46.3666661580404, 46.6666666666667, 46.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.966667175293, 41.3666661580404, 41.6666666666667, 41.966667175293, 
    42.3666661580404, 42.6666666666667, 42.966667175293, 43.3666661580404, 
    43.6666666666667, 43.966667175293, 44.3666661580404, 44.6666666666667, 
    44.966667175293, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    39.966667175293, 40.3666661580404, 40.6666666666667, 40.966667175293, 
    41.3666661580404, 41.6666666666667, 41.966667175293, 42.3666661580404, 
    42.6666666666667, 42.966667175293, 43.3666661580404, 43.6666666666667, 
    43.966667175293, 44.3666661580404, 44.6666666666667, 44.966667175293, 
    45.3666661580404, 45.6666666666667, 45.966667175293, 46.3666661580404, 
    46.6666666666667, 46.966667175293, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 38.3666661580404, 38.6666666666667, 
    38.966667175293, 39.3666661580404, 39.6666666666667, 39.966667175293, 
    40.3666661580404, 40.6666666666667, 40.966667175293, 41.3666661580404, 
    41.6666666666667, 41.966667175293, 42.3666661580404, 42.6666666666667, 
    42.966667175293, 43.3666661580404, 43.6666666666667, 43.966667175293, 
    44.3666661580404, 44.6666666666667, 44.966667175293, 45.3666661580404, 
    45.6666666666667, 45.966667175293, 46.3666661580404, 46.6666666666667, 
    46.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3666661580404, 38.6666666666667, 38.966667175293, 
    39.3666661580404, 39.6666666666667, 39.966667175293, 40.3666661580404, 
    40.6666666666667, 40.966667175293, 41.3666661580404, 41.6666666666667, 
    41.966667175293, 42.3666661580404, 42.6666666666667, 42.966667175293, 
    43.3666661580404, 43.6666666666667, 43.966667175293, 44.3666661580404, 
    44.6666666666667, 44.966667175293, 45.3666661580404, 45.6666666666667, 
    45.966667175293, 46.3666661580404, 46.6666666666667, 46.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.966667175293, 41.3666661580404, 41.6666666666667, 41.966667175293, 
    42.3666661580404, 42.6666666666667, 42.966667175293, 43.3666661580404, 
    43.6666666666667, 43.966667175293, 44.3666661580404, 44.6666666666667, 
    44.966667175293, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    39.966667175293, 40.3666661580404, 40.6666666666667, 40.966667175293, 
    41.3666661580404, 41.6666666666667, 41.966667175293, 42.3666661580404, 
    42.6666666666667, 42.966667175293, 43.3666661580404, 43.6666666666667, 
    43.966667175293, 44.3666661580404, 44.6666666666667, 44.966667175293, 
    45.3666661580404, 45.6666666666667, 45.966667175293, 46.3666661580404, 
    46.6666666666667, 46.966667175293, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 38.3666661580404, 38.6666666666667, 
    38.966667175293, 39.3666661580404, 39.6666666666667, 39.966667175293, 
    40.3666661580404, 40.6666666666667, 40.966667175293, 41.3666661580404, 
    41.6666666666667, 41.966667175293, 42.3666661580404, 42.6666666666667, 
    42.966667175293, 43.3666661580404, 43.6666666666667, 43.966667175293, 
    44.3666661580404, 44.6666666666667, 44.966667175293, 45.3666661580404, 
    45.6666666666667, 45.966667175293, 46.3666661580404, 46.6666666666667, 
    46.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3666661580404, 38.6666666666667, 38.966667175293, 
    39.3666661580404, 39.6666666666667, 39.966667175293, 40.3666661580404, 
    40.6666666666667, 40.966667175293, 41.3666661580404, 41.6666666666667, 
    41.966667175293, 42.3666661580404, 42.6666666666667, 42.966667175293, 
    43.3666661580404, 43.6666666666667, 43.966667175293, 44.3666661580404, 
    44.6666666666667, 44.966667175293, 45.3666661580404, 45.6666666666667, 
    45.966667175293, 46.3666661580404, 46.6666666666667, 46.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.966667175293, 41.3666661580404, 41.6757574370413, 41.966667175293, 
    42.3523802984328, 42.5666681925456, 42.9666668574015, 43.3666659037272, 
    43.6291672388713, 43.966667175293, 44.3666661580404, 44.6809521629697, 
    44.966667175293, 45.3566660563151, 45.6666666666667, 45.9666672908899, 
    46.3866663614909, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    39.966667175293, 40.3666661580404, 40.6666666666667, 40.966667175293, 
    41.3575752720688, 41.6666666666667, 41.966667175293, 42.3666659037272, 
    42.6380956740606, 42.9666670481364, 43.3999989827474, 43.6999994913737, 
    43.9541670481364, 44.7666651407878, 44.9666675385975, 45.3666659037272, 
    45.6666666666667, 45.966667175293, 46.4000002543131, 46.6666666666667, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.9666674296061, 41.3666661580404, 41.6666666666667, 41.9333337148031, 
    42.3809518359956, 42.5916678110759, 43.0333340962728, 43.3166662851969, 
    43.6999994913737, 43.9166666666667, 44.2666651407878, 44.6866663614909, 
    45.0000012715658, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3791662851969, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    39.966667175293, 40.3888884650336, 40.6666666666667, 41.006667582194, 
    41.3575752720688, 41.6444447835286, 41.9952385312035, 42.3952378772554, 
    42.5666681925456, 43.3166662851969, 43.6416670481364, 44.6999994913737, 
    44.9666675991482, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    40.4266665140788, 40.6791664759318, 40.9757580612645, 41.3380948021298, 
    41.6380956740606, 43.3166662851969, 43.6666666666667, 44.7041660944621, 
    44.9757580612645, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.657575896292, 46.9541670481364, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 44.9866671244303, 
    45.3666661580404, 45.6666666666667, 46.3666661580404, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3575752720688, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3766661326091, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.657575896292, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.9541670481364, 36.3791662851969, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6541668574015, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3266657511393, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6166674296061, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6166674296061, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.9541670481364, 33.3166662851969, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.9541670481364, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3523802984329, 32.6466669718424, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 34.122667948405, 
    34.122667948405, 34.122667948405, 34.122667948405, 34.122667948405, 
    34.122667948405, 34.122667948405, 34.122667948405, 34.122667948405, 
    34.122667948405, 34.122667948405, 34.122667948405, 34.122667948405, 
    34.122667948405, 34.122667948405, 34.122667948405, 34.122667948405, 
    34.122667948405, 34.122667948405, 34.122667948405, 34.122667948405, 
    34.122667948405, 34.122667948405, 34.122667948405, 34.122667948405, 
    34.122667948405, 34.122667948405, 34.122667948405, 34.122667948405, 
    34.122667948405, 34.122667948405, 34.122667948405, 34.122667948405, 
    34.122667948405, 34.122667948405, 34.122667948405, 34.122667948405, 
    34.122667948405, 34.122667948405, 34.122667948405, 34.122667948405, 
    34.122667948405, 34.122667948405, 34.122667948405, 34.122667948405, 
    34.122667948405, 42.2416674296061, 42.2416674296061, 42.2416674296061, 
    42.2416674296061, 42.2416674296061, 42.2416674296061, 42.2416674296061, 
    42.2416674296061, 42.2416674296061, 42.2416674296061, 42.2416674296061, 
    42.2416674296061, 42.2416674296061, 42.2416674296061, 42.2416674296061, 
    42.2416674296061, 42.2416674296061, 42.2416674296061, 42.2416674296061, 
    42.2416674296061, 42.2416674296061, 42.2416674296061, 42.2416674296061, 
    42.2416674296061, 42.2416674296061, 42.2416674296061, 42.2416674296061, 
    42.2416674296061, 42.2416674296061, 42.2416674296061, 42.2416674296061, 
    42.2416674296061, 42.2416674296061, 42.2416674296061, 42.2416674296061, 
    42.2416674296061, 42.2416674296061, 42.2416674296061, 42.2416674296061, 
    42.2416674296061, 42.2416674296061, 42.2416674296061, 42.2416674296061, 
    42.2416674296061, 42.2416674296061, 42.2416674296061, 44.8956667582194, 
    44.8956667582194, 44.8956667582194, 44.8956667582194, 44.8956667582194, 
    44.8956667582194, 44.8956667582194, 44.8956667582194, 44.8956667582194, 
    44.8956667582194, 44.8956667582194, 44.8956667582194, 44.8956667582194, 
    44.8956667582194, 44.8956667582194, 44.8956667582194, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    39.966667175293, 40.3666661580404, 40.6666666666667, 40.966667175293, 
    41.3666661580404, 41.6666666666667, 41.966667175293, 42.3666661580404, 
    42.6666666666667, 42.966667175293, 43.3666661580404, 43.6666666666667, 
    43.966667175293, 44.3666661580404, 44.6666666666667, 44.966667175293, 
    45.3666661580404, 45.6666666666667, 45.966667175293, 46.3666661580404, 
    46.6666666666667, 46.966667175293, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 38.3666661580404, 38.6666666666667, 
    38.966667175293, 39.3666661580404, 39.6666666666667, 39.966667175293, 
    40.3666661580404, 40.6666666666667, 40.966667175293, 41.3666661580404, 
    41.6666666666667, 41.966667175293, 42.3666661580404, 42.6666666666667, 
    42.966667175293, 43.3666661580404, 43.6666666666667, 43.966667175293, 
    44.3666661580404, 44.6666666666667, 44.966667175293, 45.3666661580404, 
    45.6666666666667, 45.966667175293, 46.3666661580404, 46.6666666666667, 
    46.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3666661580404, 38.6666666666667, 38.966667175293, 
    39.3666661580404, 39.6666666666667, 39.966667175293, 40.3666661580404, 
    40.6666666666667, 40.966667175293, 41.3666661580404, 41.6666666666667, 
    41.966667175293, 42.3666661580404, 42.6666666666667, 42.966667175293, 
    43.3666661580404, 43.6666666666667, 43.966667175293, 44.3666661580404, 
    44.6666666666667, 44.966667175293, 45.3666661580404, 45.6666666666667, 
    45.966667175293, 46.3666661580404, 46.6666666666667, 46.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.966667175293, 41.3666661580404, 41.6666666666667, 41.966667175293, 
    42.3666661580404, 42.6666666666667, 42.966667175293, 43.3666661580404, 
    43.6666666666667, 43.966667175293, 44.3666661580404, 44.6666666666667, 
    44.966667175293, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    39.966667175293, 40.3666661580404, 40.6666666666667, 40.966667175293, 
    41.3666661580404, 41.6666666666667, 41.966667175293, 42.3666661580404, 
    42.6666666666667, 42.966667175293, 43.3666661580404, 43.6666666666667, 
    43.966667175293, 44.3666661580404, 44.6666666666667, 44.966667175293, 
    45.3666661580404, 45.6666666666667, 45.966667175293, 46.3666661580404, 
    46.6666666666667, 46.966667175293, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 38.3666661580404, 38.6666666666667, 
    38.966667175293, 39.3666661580404, 39.6666666666667, 39.966667175293, 
    40.3666661580404, 40.6666666666667, 40.966667175293, 41.3666661580404, 
    41.6666666666667, 41.966667175293, 42.3666661580404, 42.6666666666667, 
    42.966667175293, 43.3666661580404, 43.6666666666667, 43.966667175293, 
    44.3666661580404, 44.6666666666667, 44.966667175293, 45.3666661580404, 
    45.6666666666667, 45.966667175293, 46.3666661580404, 46.6666666666667, 
    46.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3666661580404, 38.6666666666667, 38.966667175293, 
    39.3666661580404, 39.6666666666667, 39.966667175293, 40.3666661580404, 
    40.6666666666667, 40.966667175293, 41.3666661580404, 41.6666666666667, 
    41.966667175293, 42.3666661580404, 42.6666666666667, 42.966667175293, 
    43.3666661580404, 43.6666666666667, 43.966667175293, 44.3666661580404, 
    44.6666666666667, 44.966667175293, 45.3666661580404, 45.6666666666667, 
    45.966667175293, 46.3666661580404, 46.6666666666667, 46.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.966667175293, 41.3666661580404, 41.6666666666667, 41.966667175293, 
    42.3666661580404, 42.6666666666667, 42.966667175293, 43.3666661580404, 
    43.6666666666667, 43.966667175293, 44.3666661580404, 44.6666666666667, 
    44.966667175293, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    39.966667175293, 40.3666661580404, 40.6666666666667, 40.966667175293, 
    41.3666661580404, 41.6666666666667, 41.966667175293, 42.3666661580404, 
    42.6666666666667, 42.966667175293, 43.3666661580404, 43.6666666666667, 
    43.966667175293, 44.3666661580404, 44.6666666666667, 44.966667175293, 
    45.3666661580404, 45.6666666666667, 45.966667175293, 46.3666661580404, 
    46.6666666666667, 46.966667175293, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 38.3666661580404, 38.6666666666667, 
    38.966667175293, 39.3666661580404, 39.6666666666667, 39.966667175293, 
    40.3666661580404, 40.6666666666667, 40.966667175293, 41.3666661580404, 
    41.6666666666667, 41.966667175293, 42.3666661580404, 42.6666666666667, 
    42.966667175293, 43.3666661580404, 43.6666666666667, 43.966667175293, 
    44.3666661580404, 44.6666666666667, 44.966667175293, 45.3666661580404, 
    45.6666666666667, 45.966667175293, 46.3666661580404, 46.6666666666667, 
    46.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3666661580404, 38.6666666666667, 38.966667175293, 
    39.3666661580404, 39.6666666666667, 39.966667175293, 40.3666661580404, 
    40.6666666666667, 40.966667175293, 41.3666661580404, 41.6666666666667, 
    41.966667175293, 42.3666661580404, 42.6666666666667, 42.966667175293, 
    43.3666661580404, 43.6666666666667, 43.966667175293, 44.3666661580404, 
    44.6666666666667, 44.966667175293, 45.3666661580404, 45.6666666666667, 
    45.966667175293, 46.3666661580404, 46.6666666666667, 46.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.966667175293, 41.3666661580404, 41.6666666666667, 41.966667175293, 
    42.3666661580404, 42.6666666666667, 42.966667175293, 43.3666661580404, 
    43.6666666666667, 43.966667175293, 44.3666661580404, 44.6666666666667, 
    44.966667175293, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    39.966667175293, 40.3666661580404, 40.6666666666667, 40.966667175293, 
    41.3666661580404, 41.6666666666667, 41.966667175293, 42.3666661580404, 
    42.6666666666667, 42.966667175293, 43.3666661580404, 43.6666666666667, 
    43.966667175293, 44.3666661580404, 44.6666666666667, 44.966667175293, 
    45.3666661580404, 45.6666666666667, 45.966667175293, 46.3666661580404, 
    46.6666666666667, 46.966667175293, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 38.3666661580404, 38.6666666666667, 
    38.966667175293, 39.3666661580404, 39.6666666666667, 39.966667175293, 
    40.3666661580404, 40.6666666666667, 40.966667175293, 41.3666661580404, 
    41.6888885498047, 41.966667175293, 42.2916657129923, 42.9666668574015, 
    43.2666651407878, 43.6095246814546, 43.966667175293, 44.3666661580404, 
    44.6809521629697, 44.9666674296061, 45.3666660424435, 45.6666666666667, 
    45.9666672908899, 46.3866663614909, 46.6666666666667, 46.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.966667175293, 41.3575752720688, 41.6777776082357, 41.966667175293, 
    42.3666659037272, 42.6500002543132, 42.9666670481364, 43.2666651407878, 
    43.6166674296061, 43.9541670481364, 44.7666651407878, 44.9666678110758, 
    45.3666659037272, 45.6666666666667, 45.966667175293, 46.4000002543131, 
    46.6666666666667, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3666661580404, 38.6666666666667, 38.966667175293, 
    39.3666661580404, 39.6666666666667, 39.966667175293, 40.3666661580404, 
    40.6666666666667, 40.9416672388713, 41.3666655222575, 41.6999994913737, 
    41.9000002543132, 42.3809518359956, 42.5916678110759, 43.0333340962728, 
    43.3666674296061, 43.6866663614909, 43.9166666666667, 44.2666651407878, 
    44.7666651407878, 45.0000012715658, 45.3666661580404, 45.6666666666667, 
    45.966667175293, 46.3666661580404, 46.6666666666667, 46.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.9575761737245, 40.3888884650336, 40.6566668192546, 
    40.8666674296061, 41.3466654459635, 41.5666681925456, 42.3916670481364, 
    42.5666681925456, 43.3166662851969, 43.7166659037272, 44.7166659037272, 
    44.9666675991482, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    40.4266665140788, 40.6791664759318, 40.966667175293, 41.6666666666667, 
    43.7166659037272, 44.7041660944621, 44.9757580612645, 45.3666661580404, 
    45.6666666666667, 45.966667175293, 46.3666661580404, 46.657575896292, 
    46.9541670481364, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3666661580404, 38.6666666666667, 38.966667175293, 
    39.3666661580404, 44.9866671244303, 45.3666661580404, 45.6666666666667, 
    46.3666661580404, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3575752720688, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3766661326091, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.657575896292, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.9541670481364, 
    36.3791662851969, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6541668574015, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3266657511393, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6166674296061, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6166674296061, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.9541670481364, 33.3166662851969, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.9541670481364, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3523802984329, 32.6466669718424, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 41.2626673380534, 41.2626673380534, 41.2626673380534, 
    41.2626673380534, 41.2626673380534, 41.2626673380534, 41.2626673380534, 
    41.2626673380534, 41.2626673380534, 41.2626673380534, 41.2626673380534, 
    41.2626673380534, 41.2626673380534, 40.8836657206217, 40.8836657206217, 
    40.8836657206217, 40.8836657206217, 40.8836657206217, 40.8836657206217, 
    40.8836657206217, 40.8836657206217, 40.8836657206217, 40.8836657206217, 
    40.8836657206217, 40.8836657206217, 40.8836657206217, 40.8836657206217, 
    32.6146685282389, 32.6146685282389, 32.6146685282389, 32.6146685282389, 
    32.6146685282389, 32.6146685282389, 32.6146685282389, 32.6146685282389, 
    32.6146685282389, 32.6146685282389, 32.6146685282389, 32.6146685282389, 
    32.6146685282389, 32.6146685282389, 32.5836664835612, 32.5836664835612, 
    32.5836664835612, 32.5836664835612, 32.5836664835612, 32.5836664835612, 
    32.5836664835612, 32.5836664835612, 32.5836664835612, 32.5836664835612, 
    32.5836664835612, 32.5836664835612, 32.5836664835612, 32.5836664835612, 
    32.5836664835612, 32.5836664835612, 32.5836664835612, 32.5836664835612, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.966667175293, 41.3666661580404, 41.6666666666667, 41.966667175293, 
    42.3666661580404, 42.6666666666667, 42.966667175293, 43.3666661580404, 
    43.6666666666667, 43.966667175293, 44.3666661580404, 44.6666666666667, 
    44.966667175293, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    39.966667175293, 40.3666661580404, 40.6666666666667, 40.966667175293, 
    41.3666661580404, 41.6666666666667, 41.966667175293, 42.3666661580404, 
    42.6666666666667, 42.966667175293, 43.3666661580404, 43.6666666666667, 
    43.966667175293, 44.3666661580404, 44.6666666666667, 44.966667175293, 
    45.3666661580404, 45.6666666666667, 45.966667175293, 46.3666661580404, 
    46.6666666666667, 46.966667175293, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 38.3666661580404, 38.6666666666667, 
    38.966667175293, 39.3666661580404, 39.6666666666667, 39.966667175293, 
    40.3666661580404, 40.6666666666667, 40.966667175293, 41.3666661580404, 
    41.6666666666667, 41.966667175293, 42.3666661580404, 42.6666666666667, 
    42.966667175293, 43.3666661580404, 43.6666666666667, 43.966667175293, 
    44.3666661580404, 44.6666666666667, 44.966667175293, 45.3666661580404, 
    45.6666666666667, 45.966667175293, 46.3666661580404, 46.6666666666667, 
    46.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3666661580404, 38.6666666666667, 38.966667175293, 
    39.3666661580404, 39.6666666666667, 39.966667175293, 40.3666661580404, 
    40.6666666666667, 40.966667175293, 41.3666661580404, 41.6666666666667, 
    41.966667175293, 42.3666661580404, 42.6666666666667, 42.966667175293, 
    43.3666661580404, 43.6666666666667, 43.966667175293, 44.3666661580404, 
    44.6666666666667, 44.966667175293, 45.3666661580404, 45.6666666666667, 
    45.966667175293, 46.3666661580404, 46.6666666666667, 46.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.966667175293, 41.3666661580404, 41.6666666666667, 41.966667175293, 
    42.3666661580404, 42.6666666666667, 42.966667175293, 43.3666661580404, 
    43.6666666666667, 43.966667175293, 44.3666661580404, 44.6666666666667, 
    44.966667175293, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    39.966667175293, 40.3666661580404, 40.6666666666667, 40.966667175293, 
    41.3666661580404, 41.6666666666667, 41.966667175293, 42.3666661580404, 
    42.6666666666667, 42.966667175293, 43.3666661580404, 43.6666666666667, 
    43.966667175293, 44.3666661580404, 44.6666666666667, 44.966667175293, 
    45.3666661580404, 45.6666666666667, 45.966667175293, 46.3666661580404, 
    46.6666666666667, 46.966667175293, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 38.3666661580404, 38.6666666666667, 
    38.966667175293, 39.3666661580404, 39.6666666666667, 39.966667175293, 
    40.3666661580404, 40.6666666666667, 40.966667175293, 41.3666661580404, 
    41.6666666666667, 41.966667175293, 42.3666661580404, 42.6666666666667, 
    42.966667175293, 43.3666661580404, 43.6666666666667, 43.966667175293, 
    44.3666661580404, 44.6666666666667, 44.966667175293, 45.3666661580404, 
    45.6666666666667, 45.966667175293, 46.3666661580404, 46.6666666666667, 
    46.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3666661580404, 38.6666666666667, 38.966667175293, 
    39.3666661580404, 39.6666666666667, 39.966667175293, 40.3666661580404, 
    40.6666666666667, 40.966667175293, 41.3666661580404, 41.6666666666667, 
    41.966667175293, 42.3666661580404, 42.6666666666667, 42.966667175293, 
    43.3666661580404, 43.6666666666667, 43.966667175293, 44.3666661580404, 
    44.6666666666667, 44.966667175293, 45.3666661580404, 45.6666666666667, 
    45.966667175293, 46.3666661580404, 46.6666666666667, 46.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.966667175293, 41.3666661580404, 41.6666666666667, 41.966667175293, 
    42.3666661580404, 42.6666666666667, 42.966667175293, 43.3666661580404, 
    43.6666666666667, 43.966667175293, 44.3666661580404, 44.6666666666667, 
    44.966667175293, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    39.966667175293, 40.3666661580404, 40.6666666666667, 40.966667175293, 
    41.3666661580404, 41.6666666666667, 41.966667175293, 42.3666661580404, 
    42.6666666666667, 42.966667175293, 43.3666661580404, 43.6666666666667, 
    43.966667175293, 44.3666661580404, 44.6666666666667, 44.966667175293, 
    45.3666661580404, 45.6666666666667, 45.966667175293, 46.3666661580404, 
    46.6666666666667, 46.966667175293, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 38.3666661580404, 38.6666666666667, 
    38.966667175293, 39.3666661580404, 39.6666666666667, 39.966667175293, 
    40.3666661580404, 40.6666666666667, 40.966667175293, 41.3666661580404, 
    41.6666666666667, 41.966667175293, 42.3666661580404, 42.6666666666667, 
    42.966667175293, 43.3666661580404, 43.6666666666667, 43.966667175293, 
    44.3666661580404, 44.6666666666667, 44.966667175293, 45.3666661580404, 
    45.6666666666667, 45.966667175293, 46.3666661580404, 46.6666666666667, 
    46.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3666661580404, 38.6666666666667, 38.966667175293, 
    39.3666661580404, 39.6666666666667, 39.966667175293, 40.3666661580404, 
    40.6666666666667, 40.966667175293, 41.3666661580404, 41.6666666666667, 
    41.966667175293, 42.3666661580404, 42.6666666666667, 42.966667175293, 
    43.3666661580404, 43.6666666666667, 43.966667175293, 44.3666661580404, 
    44.6666666666667, 44.966667175293, 45.3666661580404, 45.6666666666667, 
    45.966667175293, 46.3666661580404, 46.6666666666667, 46.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.966667175293, 41.3666661580404, 41.6666666666667, 41.966667175293, 
    42.3666661580404, 42.6666666666667, 42.966667175293, 43.3666661580404, 
    43.6666666666667, 43.966667175293, 44.3666661580404, 44.6666666666667, 
    44.966667175293, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666660424435, 39.6666666666667, 
    39.9575761737245, 40.3666661580404, 40.6666666666667, 40.966667175293, 
    41.3575752720688, 41.6809521629697, 41.9541670481364, 42.3666674296061, 
    43.966667175293, 44.3666662851969, 44.6791664759318, 44.955556233724, 
    45.3666660424435, 45.6666666666667, 45.966667175293, 46.3666661580404, 
    46.6666666666667, 46.966667175293, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 38.3666661580404, 38.6666666666667, 
    38.966667175293, 39.3666660424435, 39.6666666666667, 39.966667175293, 
    40.3666660424435, 40.6266672770182, 41.0095245724633, 41.3291660944621, 
    41.6999994913737, 41.9333335028754, 42.3166662851969, 44.3916670481364, 
    44.7166659037272, 44.916667620341, 45.3766661326091, 45.6666666666667, 
    45.966667175293, 46.3666661580403, 46.6666666666667, 46.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.9541670481364, 39.3541661898295, 
    39.6666666666667, 39.9523814973377, 40.3266657511393, 41.2666651407878, 
    41.7666651407878, 44.7166659037272, 45.0000006357829, 45.3666661580404, 
    45.6666666666667, 45.966667175293, 46.3666661580404, 46.6666666666667, 
    46.9541670481364, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3666661580404, 38.6666666666667, 38.966667175293, 
    39.3575752720688, 39.657575896292, 40.4041663805644, 40.6566668192546, 
    40.8666674296061, 42.5666681925456, 44.7166659037272, 44.9666674296061, 
    45.3666661580404, 45.6666666666667, 45.966667175293, 46.3666661580404, 
    46.6666666666667, 46.966667175293, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 38.3666661580404, 38.6666666666667, 
    38.966667175293, 39.3666661580404, 39.6380956740606, 40.4266665140788, 
    40.6666666666667, 40.8666674296061, 44.7041660944621, 44.9757580612645, 
    45.3666661580404, 45.6666666666667, 45.966667175293, 46.3666661580404, 
    46.657575896292, 46.9541670481364, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 38.3666661580404, 38.6666666666667, 
    38.966667175293, 39.3666661580404, 44.9866671244303, 45.3666661580404, 
    45.6666666666667, 46.3666661580404, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 38.3575752720688, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.657575896292, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.9541670481364, 36.3791662851969, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6541668574015, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3266657511393, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6166674296061, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6166674296061, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.9541670481364, 33.3166662851969, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.9541670481364, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3523802984329, 
    32.6466669718424, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 32.3496653238932, 32.3496653238932, 
    32.3496653238932, 32.3496653238932, 32.3496653238932, 32.3496653238932, 
    32.3496653238932, 32.3496653238932, 32.3496653238932, 32.3496653238932, 
    32.3496653238932, 32.3496653238932, 32.3496653238932, 32.3496653238932, 
    32.3496653238932, 32.3496653238932, 32.3496653238932, 32.3496653238932, 
    32.013666788737, 32.013666788737, 32.013666788737, 32.013666788737, 
    32.013666788737, 32.013666788737, 32.013666788737, 32.013666788737, 
    32.013666788737, 32.013666788737, 32.013666788737, 32.013666788737, 
    32.013666788737, 32.013666788737, 32.013666788737, 32.013666788737, 
    32.013666788737, 32.013666788737, 32.013666788737, 32.013666788737, 
    32.013666788737, 32.013666788737, 32.013666788737, 32.013666788737, 
    32.013666788737, 32.013666788737, 32.013666788737, 32.013666788737, 
    32.013666788737, 32.013666788737, 30.6170631237561, 30.6170631237561, 
    30.9025056550392, 30.6170631237561, 30.9025056550392, 30.6170631237561, 
    30.9025056550392, 30.6170631237561, 30.9025056550392, 31.7536566677173, 
    30.6170631237561, 30.9025056550392, 31.7536566677173, 30.6170631237561, 
    32.0356337743697, 30.9025056550392, 31.7536566677173, 30.6170631237561, 
    32.0356337743697, 30.9025056550392, 31.7536566677173, 32.3167339917995, 
    30.6170631237561, 32.0356337743697, 30.9025056550392, 31.7536566677173, 
    32.3167339917995, 30.6170631237561, 32.0356337743697, 32.5969533019733, 
    30.9025056550392, 31.7536566677173, 32.3167339917995, 30.6170631237561, 
    32.0356337743697, 32.5969533019733, 30.9025056550392, 31.7536566677173, 
    32.3167339917995, 30.6170631237561, 32.8762877838633, 32.0356337743697, 
    32.5969533019733, 30.9025056550392, 31.7536566677173, 32.3167339917995, 
    30.6170631237561, 32.8762877838633, 32.0356337743697, 32.5969533019733, 
    30.9025056550392, 33.432287061478, 31.7536566677173, 32.3167339917995, 
    30.6170631237561, 32.8762877838633, 32.0356337743697, 32.5969533019733, 
    30.9025056550392, 33.432287061478, 31.7536566677173, 32.3167339917995, 
    30.6170631237561, 32.8762877838633, 33.7089444967663, 32.0356337743697, 
    32.5969533019733, 30.9025056550392, 33.432287061478, 31.7536566677173, 
    32.3167339917995, 30.6170631237561, 32.8762877838633, 33.7089444967663, 
    32.0356337743697, 32.5969533019733, 30.9025056550392, 33.432287061478, 
    31.7536566677173, 33.9847023820702, 32.3167339917995, 30.6170631237561, 
    32.8762877838633, 33.7089444967663, 32.0356337743697, 32.5969533019733, 
    30.9025056550392, 33.432287061478, 31.7536566677173, 33.9847023820702, 
    32.3167339917995, 30.6170631237561, 32.8762877838633, 33.7089444967663, 
    32.0356337743697, 34.2595572754987, 32.5969533019733, 30.9025056550392, 
    33.432287061478, 31.7536566677173, 33.9847023820702, 32.3167339917995, 
    30.6170631237561, 32.8762877838633, 33.7089444967663, 32.0356337743697, 
    34.2595572754987, 32.5969533019733, 30.9025056550392, 33.432287061478, 
    31.7536566677173, 33.9847023820702, 32.3167339917995, 30.6170631237561, 
    34.5335058296867, 32.8762877838633, 33.7089444967663, 32.0356337743697, 
    34.2595572754987, 32.5969533019733, 30.9025056550392, 33.432287061478, 
    31.7536566677173, 33.9847023820702, 32.3167339917995, 30.6170631237561, 
    34.5335058296867, 32.8762877838633, 33.7089444967663, 32.0356337743697, 
    34.2595572754987, 32.5969533019733, 30.9025056550392, 35.0786710006513, 
    33.432287061478, 31.7536566677173, 33.9847023820702, 32.3167339917995, 
    30.6170631237561, 34.5335058296867, 32.8762877838633, 33.7089444967663, 
    32.0356337743697, 34.2595572754987, 32.5969533019733, 30.9025056550392, 
    35.0786710006513, 33.432287061478, 31.7536566677173, 33.9847023820702, 
    32.3167339917995, 30.6170631237561, 34.5335058296867, 32.8762877838633, 
    35.3498813909852, 33.7089444967663, 32.0356337743697, 34.2595572754987, 
    32.5969533019733, 30.9025056550392, 35.0786710006513, 33.432287061478, 
    31.7536566677173, 33.9847023820702, 32.3167339917995, 30.6170631237561, 
    34.5335058296867, 32.8762877838633, 35.3498813909852, 33.7089444967663, 
    32.0356337743697, 34.2595572754987, 32.5969533019733, 30.9025056550392, 
    35.0786710006513, 33.432287061478, 31.7536566677173, 35.620172988168, 
    33.9847023820702, 32.3167339917995, 30.6170631237561, 34.5335058296867, 
    32.8762877838633, 35.3498813909853, 33.7089444967663, 32.0356337743697, 
    34.2595572754987, 32.5969533019733, 30.9025056550392, 35.0786710006513, 
    33.432287061478, 31.7536566677173, 35.620172988168, 33.9847023820702, 
    32.3167339917995, 30.6170631237561, 34.5335058296867, 32.8762877838633, 
    35.3498813909852, 33.7089444967663, 32.0356337743697, 35.8895429100474, 
    34.2595572754987, 32.5969533019733, 30.9025056550392, 35.0786710006513, 
    33.432287061478, 31.7536566677173, 35.620172988168, 33.9847023820702, 
    32.3167339917995, 30.6170631237561, 34.5335058296867, 32.8762877838633, 
    35.3498813909852, 33.7089444967663, 32.0356337743697, 35.8895429100474, 
    34.2595572754987, 32.5969533019733, 30.9025056550392, 35.0786710006513, 
    33.432287061478, 31.7536566677173, 35.620172988168, 33.9847023820702, 
    32.3167339917995, 36.4255066559906, 30.6170631237561, 34.5335058296867, 
    32.8762877838633, 35.3498813909852, 33.7089444967663, 32.0356337743697, 
    35.8895429100474, 34.2595572754987, 32.5969533019733, 30.9025056550392, 
    35.0786710006513, 33.432287061478, 31.7536566677173, 35.620172988168, 
    33.9847023820702, 32.3167339917995, 36.4255066559906, 30.6170631237561, 
    34.5335058296867, 32.8762877838633, 35.3498813909852, 33.7089444967663, 
    32.0356337743697, 35.8895429100474, 34.2595572754987, 32.5969533019733, 
    36.6920951707497, 30.9025056550392, 35.0786710006513, 33.432287061478, 
    31.7536566677173, 35.620172988168, 33.9847023820702, 32.3167339917995, 
    36.4255066559906, 30.6170631237561, 34.5335058296867, 32.8762877838633, 
    35.3498813909852, 33.7089444967663, 32.0356337743697, 35.8895429100474, 
    34.2595572754987, 32.5969533019733, 36.6920951707497, 30.9025056550392, 
    35.0786710006513, 33.432287061478, 31.7536566677173, 35.620172988168, 
    33.9847023820702, 32.3167339917995, 36.4255066559906, 30.6170631237561, 
    34.5335058296867, 32.8762877838633, 36.9577513904295, 35.3498813909852, 
    33.7089444967663, 32.0356337743697, 35.8895429100474, 34.2595572754987, 
    32.5969533019733, 36.6920951707497, 30.9025056550392, 35.0786710006513, 
    33.432287061478, 31.7536566677173, 35.620172988168, 33.9847023820702, 
    32.3167339917995, 36.4255066559906, 30.6170631237561, 34.5335058296867, 
    32.8762877838633, 36.9577513904295, 35.3498813909852, 33.7089444967663, 
    32.0356337743697, 35.8895429100474, 34.2595572754987, 32.5969533019733, 
    36.6920951707497, 30.9025056550392, 35.0786710006513, 33.432287061478, 
    37.2224728843778, 31.7536566677173, 35.620172988168, 33.9847023820702, 
    32.3167339917995, 36.4255066559906, 30.6170631237561, 34.5335058296867, 
    32.8762877838633, 36.9577513904295, 35.3498813909853, 33.7089444967663, 
    32.0356337743697, 35.8895429100474, 34.2595572754987, 32.5969533019733, 
    36.6920951707497, 30.9025056550392, 35.0786710006513, 33.432287061478, 
    37.2224728843778, 31.7536566677173, 35.620172988168, 33.9847023820702, 
    32.3167339917995, 36.4255066559906, 30.6170631237561, 34.5335058296867, 
    32.8762877838633, 36.9577513904295, 35.3498813909852, 33.7089444967663, 
    37.7491024143739, 32.0356337743697, 35.8895429100474, 34.2595572754987, 
    32.5969533019733, 36.6920951707497, 30.9025056550392, 35.0786710006513, 
    33.432287061478, 37.2224728843778, 31.7536566677173, 35.620172988168, 
    33.9847023820702, 32.3167339917995, 36.4255066559906, 30.6170631237561, 
    34.5335058296867, 32.8762877838633, 36.9577513904295, 35.3498813909852, 
    33.7089444967663, 37.749102414374, 32.0356337743697, 35.8895429100474, 
    34.2595572754987, 32.5969533019733, 36.6920951707497, 30.9025056550392, 
    35.0786710006513, 33.432287061478, 37.2224728843778, 31.7536566677173, 
    35.620172988168, 33.9847023820702, 38.0110060291271, 32.3167339917995, 
    36.4255066559906, 30.6170631237561, 34.5335058296867, 32.8762877838633, 
    36.9577513904295, 35.3498813909852, 33.7089444967663, 37.7491024143739, 
    32.0356337743697, 35.8895429100474, 34.2595572754987, 32.5969533019733, 
    36.6920951707497, 30.9025056550392, 35.0786710006513, 33.432287061478, 
    37.2224728843778, 31.7536566677173, 35.620172988168, 33.9847023820702, 
    38.0110060291271, 32.3167339917995, 36.4255066559906, 30.6170631237561, 
    34.5335058296867, 32.8762877838633, 36.9577513904295, 35.3498813909852, 
    33.7089444967663, 37.7491024143739, 32.0356337743697, 35.8895429100474, 
    34.2595572754987, 38.2719660742721, 32.5969533019733, 36.6920951707497, 
    30.9025056550392, 35.0786710006513, 33.432287061478, 37.2224728843778, 
    31.7536566677173, 35.620172988168, 33.9847023820702, 38.0110060291271, 
    32.3167339917995, 36.4255066559906, 30.6170631237561, 34.5335058296867, 
    32.8762877838633, 36.9577513904295, 35.3498813909852, 33.7089444967663, 
    37.7491024143739, 32.0356337743697, 35.8895429100474, 34.2595572754987, 
    38.2719660742721, 32.5969533019733, 36.6920951707497, 30.9025056550392, 
    35.0786710006513, 33.432287061478, 37.2224728843778, 31.7536566677173, 
    35.620172988168, 33.9847023820702, 38.0110060291271, 32.3167339917995, 
    36.4255066559906, 30.6170631237561, 34.5335058296867, 38.6615140591414, 
    32.8762877838633, 36.9577513904295, 35.3498813909852, 33.7089444967663, 
    37.7491024143739, 32.0356337743697, 35.8895429100474, 34.2595572754987, 
    38.2719660742721, 32.5969533019733, 36.6920951707497, 30.9025056550392, 
    35.0786710006513, 33.432287061478, 37.2224728843778, 31.7536566677173, 
    35.620172988168, 33.9847023820702, 38.0110060291271, 32.3167339917995, 
    36.4255066559906, 30.6170631237561, 34.5335058296867, 38.6615140591413, 
    32.8762877838633, 36.9577513904295, 35.3498813909852, 33.7089444967663, 
    37.7491024143739, 32.0356337743697, 35.8895429100474, 34.2595572754987, 
    38.2719660742721, 32.5969533019733, 36.6920951707497, 30.9025056550392, 
    35.0786710006513, 39.049165272633, 33.432287061478, 37.2224728843778, 
    31.7536566677173, 35.620172988168, 33.9847023820702, 38.0110060291271, 
    32.3167339917995, 36.4255066559906, 30.6170631237561, 34.5335058296867, 
    38.6615140591414, 32.8762877838633, 36.9577513904295, 35.3498813909852, 
    33.7089444967663, 37.7491024143739, 32.0356337743697, 35.8895429100474, 
    34.2595572754987, 38.2719660742721, 32.5969533019733, 36.6920951707497, 
    30.9025056550392, 35.0786710006513, 39.049165272633, 33.432287061478, 
    37.2224728843778, 31.7536566677173, 35.620172988168, 33.9847023820702, 
    38.0110060291271, 32.3167339917995, 36.4255066559906, 30.6170631237561, 
    34.5335058296867, 38.6615140591414, 32.8762877838633, 36.9577513904295, 
    35.3498813909853, 39.3063319434942, 33.7089444967663, 37.7491024143739, 
    32.0356337743697, 35.8895429100474, 34.2595572754987, 38.2719660742721, 
    32.5969533019733, 36.6920951707497, 30.9025056550392, 35.0786710006513, 
    39.049165272633, 33.432287061478, 37.2224728843778, 31.7536566677173, 
    35.620172988168, 33.9847023820702, 38.0110060291271, 32.3167339917995, 
    36.4255066559906, 30.6170631237561, 34.5335058296867, 38.6615140591414, 
    32.8762877838633, 36.9577513904295, 35.3498813909852, 39.3063319434942, 
    33.7089444967663, 37.7491024143739, 32.0356337743697, 35.8895429100474, 
    34.2595572754987, 38.2719660742721, 32.5969533019733, 36.6920951707497, 
    30.9025056550392, 35.0786710006513, 39.049165272633, 33.432287061478, 
    37.2224728843778, 31.7536566677173, 35.620172988168, 39.5625459179821, 
    33.9847023820702, 38.0110060291271, 32.3167339917995, 36.4255066559906, 
    30.6170631237561, 34.5335058296867, 38.6615140591414, 32.8762877838633, 
    36.9577513904295, 35.3498813909852, 39.3063319434942, 33.7089444967663, 
    37.7491024143739, 32.0356337743697, 35.8895429100474, 34.2595572754987, 
    38.2719660742721, 32.5969533019733, 36.6920951707497, 30.9025056550392, 
    35.0786710006513, 39.049165272633, 33.432287061478, 37.2224728843778, 
    31.7536566677173, 35.620172988168, 39.5625459179821, 33.9847023820702, 
    38.0110060291271, 32.3167339917995, 36.4255066559906, 30.6170631237561, 
    34.5335058296867, 38.6615140591414, 32.8762877838633, 36.9577513904295, 
    35.3498813909853, 39.3063319434942, 33.7089444967663, 37.7491024143739, 
    32.0356337743697, 35.8895429100474, 40.0721095592252, 34.2595572754987, 
    38.2719660742721, 32.5969533019733, 36.6920951707497, 30.9025056550392, 
    35.0786710006513, 39.049165272633, 33.432287061478, 37.2224728843778, 
    31.7536566677173, 35.620172988168, 39.5625459179821, 33.9847023820702, 
    38.0110060291271, 32.3167339917995, 36.4255066559906, 30.6170631237561, 
    34.5335058296867, 38.6615140591414, 32.8762877838633, 36.9577513904295, 
    35.3498813909852, 39.3063319434942, 33.7089444967663, 37.749102414374, 
    32.0356337743697, 35.8895429100474, 40.0721095592252, 34.2595572754987, 
    38.2719660742721, 32.5969533019733, 36.6920951707497, 30.9025056550392, 
    35.0786710006513, 39.049165272633, 33.432287061478, 37.2224728843778, 
    31.7536566677173, 35.620172988168, 39.5625459179821, 33.9847023820702, 
    38.0110060291271, 32.3167339917995, 36.4255066559906, 40.3254563203728, 
    30.6170631237561, 34.5335058296867, 38.6615140591414, 32.8762877838633, 
    36.9577513904295, 35.3498813909852, 39.3063319434942, 33.7089444967663, 
    37.7491024143739, 32.0356337743697, 35.8895429100474, 40.0721095592252, 
    34.2595572754987, 38.2719660742721, 32.5969533019733, 36.6920951707497, 
    30.9025056550392, 35.0786710006513, 39.049165272633, 33.432287061478, 
    37.2224728843778, 31.7536566677173, 35.620172988168, 39.5625459179821, 
    33.9847023820702, 38.0110060291271, 32.3167339917995, 36.4255066559906, 
    40.3254563203728, 30.6170631237561, 34.5335058296867, 38.6615140591413, 
    32.8762877838633, 36.9577513904295, 35.3498813909852, 39.3063319434942, 
    33.7089444967663, 37.7491024143739, 32.0356337743697, 35.8895429100474, 
    40.0721095592252, 34.2595572754987, 38.2719660742721, 32.5969533019733, 
    36.6920951707497, 40.5778445724771, 30.9025056550392, 35.0786710006513, 
    39.049165272633, 33.432287061478, 37.2224728843778, 31.7536566677173, 
    35.620172988168, 39.5625459179821, 33.9847023820702, 38.0110060291271, 
    32.3167339917995, 36.4255066559906, 40.3254563203728, 30.6170631237561, 
    34.5335058296867, 38.6615140591414, 32.8762877838633, 36.9577513904294, 
    35.3498813909852, 39.3063319434942, 33.7089444967663, 37.7491024143739, 
    32.0356337743697, 35.8895429100474, 40.0721095592252, 34.2595572754987, 
    38.2719660742721, 32.5969533019733, 36.6920951707497, 40.5778445724771, 
    30.9025056550392, 35.0786710006513, 39.049165272633, 33.432287061478, 
    37.2224728843778, 31.7536566677173, 35.620172988168, 39.5625459179821, 
    33.9847023820702, 38.0110060291271, 32.3167339917995, 36.4255066559906, 
    40.3254563203728, 30.6170631237561, 34.5335058296867, 38.6615140591414, 
    32.8762877838633, 36.9577513904295, 41.0797406188206, 35.3498813909852, 
    39.3063319434942, 33.7089444967663, 37.7491024143739, 32.0356337743697, 
    35.8895429100474, 40.0721095592252, 34.2595572754987, 38.2719660742721, 
    32.5969533019733, 36.6920951707497, 40.5778445724771, 30.9025056550392, 
    35.0786710006513, 39.049165272633, 33.432287061478, 37.2224728843778, 
    31.7536566677173, 35.620172988168, 39.5625459179821, 33.9847023820702, 
    38.0110060291271, 32.3167339917995, 36.4255066559906, 40.3254563203728, 
    34.5335058296867, 38.6615140591414, 32.8762877838633, 36.9577513904295, 
    41.0797406188206, 35.3498813909852, 39.3063319434942, 33.7089444967663, 
    37.7491024143739, 32.0356337743697, 35.8895429100474, 40.0721095592252, 
    34.2595572754987, 38.2719660742721, 32.5969533019733, 36.6920951707497, 
    40.5778445724771, 30.9025056550392, 35.0786710006513, 39.049165272633, 
    33.432287061478, 37.2224728843778, 41.3292461440167, 31.7536566677173, 
    35.620172988168, 39.5625459179821, 33.9847023820702, 38.0110060291271, 
    32.3167339917995, 36.4255066559906, 40.3254563203728, 34.5335058296867, 
    38.6615140591414, 32.8762877838633, 36.9577513904295, 41.0797406188206, 
    35.3498813909852, 39.3063319434942, 33.7089444967663, 37.7491024143739, 
    32.0356337743697, 35.8895429100474, 40.0721095592252, 34.2595572754987, 
    38.2719660742721, 32.5969533019733, 36.6920951707497, 40.5778445724771, 
    35.0786710006513, 39.049165272633, 33.432287061478, 37.2224728843778, 
    41.3292461440167, 31.7536566677173, 35.620172988168, 39.5625459179821, 
    33.9847023820702, 38.0110060291271, 32.3167339917995, 36.4255066559906, 
    40.3254563203728, 34.5335058296867, 38.6615140591413, 32.8762877838633, 
    36.9577513904295, 41.0797406188206, 35.3498813909852, 39.3063319434942, 
    33.7089444967663, 37.7491024143739, 41.5777886205734, 32.0356337743697, 
    35.8895429100474, 40.0721095592252, 34.2595572754987, 38.2719660742721, 
    32.5969533019733, 36.6920951707497, 40.5778445724771, 35.0786710006513, 
    39.049165272633, 33.432287061478, 37.2224728843778, 41.3292461440167, 
    31.7536566677173, 35.620172988168, 39.5625459179821, 33.9847023820702, 
    38.0110060291271, 32.3167339917995, 36.4255066559906, 40.3254563203728, 
    34.5335058296867, 38.6615140591414, 32.8762877838633, 36.9577513904295, 
    41.0797406188206, 35.3498813909852, 39.3063319434942, 33.7089444967663, 
    37.7491024143739, 41.5777886205734, 32.0356337743697, 35.8895429100474, 
    40.0721095592252, 34.2595572754987, 38.2719660742721, 32.5969533019733, 
    36.6920951707497, 40.5778445724771, 35.0786710006513, 39.049165272633, 
    33.432287061478, 37.2224728843778, 41.3292461440167, 35.620172988168, 
    39.5625459179821, 33.9847023820702, 38.0110060291271, 42.0719807371405, 
    32.3167339917995, 36.4255066559906, 40.3254563203728, 34.5335058296867, 
    38.6615140591414, 32.8762877838633, 36.9577513904295, 41.0797406188206, 
    35.3498813909852, 39.3063319434942, 33.7089444967663, 37.7491024143739, 
    41.5777886205734, 35.8895429100474, 40.0721095592252, 34.2595572754987, 
    38.2719660742721, 36.6920951707497, 40.5778445724771, 35.0786710006513, 
    39.049165272633, 33.432287061478, 37.2224728843778, 41.3292461440167, 
    35.620172988168, 39.5625459179821, 33.9847023820702, 38.0110060291271, 
    42.0719807371405, 32.3167339917995, 36.4255066559906, 40.3254563203728, 
    34.5335058296867, 38.6615140591413, 32.8762877838633, 36.9577513904295, 
    41.0797406188206, 35.3498813909852, 39.3063319434942, 37.749102414374, 
    41.5777886205734, 35.8895429100474, 40.0721095592252, 38.2719660742721, 
    42.3176287205335, 36.6920951707497, 40.5778445724771, 35.0786710006513, 
    39.049165272633, 33.432287061478, 37.2224728843778, 41.3292461440167, 
    35.620172988168, 39.5625459179821, 33.9847023820702, 38.0110060291271, 
    42.0719807371405, 36.4255066559906, 40.3254563203728, 34.5335058296867, 
    38.6615140591414, 36.9577513904295, 41.0797406188206, 35.3498813909852, 
    39.3063319434942, 37.7491024143739, 41.5777886205734, 35.8895429100474, 
    40.0721095592252, 38.2719660742721, 42.3176287205335, 36.6920951707497, 
    40.5778445724771, 35.0786710006513, 39.049165272633, 33.432287061478, 
    37.2224728843778, 41.3292461440167, 35.620172988168, 39.5625459179821, 
    38.0110060291271, 42.0719807371405, 36.4255066559906, 40.3254563203728, 
    38.6615140591414, 42.5623103404995, 36.9577513904295, 41.0797406188206, 
    35.3498813909852, 39.3063319434942, 37.7491024143739, 41.5777886205734, 
    35.8895429100474, 40.0721095592252, 38.2719660742721, 42.3176287205335, 
    36.6920951707497, 40.5778445724771, 39.049165272633, 37.2224728843778, 
    41.3292461440167, 35.620172988168, 39.5625459179821, 38.0110060291271, 
    42.0719807371405, 36.4255066559906, 40.3254563203728, 38.6615140591414, 
    42.5623103404995, 36.9577513904295, 41.0797406188206, 39.3063319434942, 
    37.7491024143739, 41.5777886205734, 35.8895429100474, 40.0721095592252, 
    38.2719660742721, 42.3176287205335, 36.6920951707497, 40.5778445724771, 
    39.049165272633, 43.0487719903617, 37.2224728843778, 41.3292461440167, 
    39.5625459179821, 38.0110060291271, 42.0719807371405, 36.4255066559906, 
    40.3254563203728, 38.6615140591414, 42.5623103404995, 36.9577513904295, 
    41.0797406188206, 39.3063319434942, 37.749102414374, 41.5777886205734, 
    40.0721095592252, 38.2719660742721, 42.3176287205335, 36.6920951707497, 
    40.5778445724771, 39.049165272633, 43.0487719903617, 37.2224728843778, 
    41.3292461440167, 39.5625459179821, 38.0110060291271, 42.0719807371405, 
    36.4255066559906, 40.3254563203728, 38.6615140591414, 42.5623103404995, 
    36.9577513904295, 41.0797406188206, 39.3063319434942, 43.2905509512355, 
    37.7491024143739, 41.5777886205734, 40.0721095592252, 38.2719660742721, 
    42.3176287205335, 36.6920951707497, 40.5778445724771, 39.049165272633, 
    43.0487719903617, 37.2224728843778, 41.3292461440167, 39.5625459179821, 
    38.0110060291271, 42.0719807371405, 40.3254563203728, 38.6615140591414, 
    42.5623103404995, 36.9577513904295, 41.0797406188206, 39.3063319434942, 
    43.2905509512355, 37.7491024143739, 41.5777886205734, 40.0721095592252, 
    38.2719660742721, 42.3176287205335, 40.5778445724771, 39.049165272633, 
    43.0487719903617, 37.2224728843778, 41.3292461440167, 39.5625459179821, 
    43.7712030066013, 38.0110060291271, 42.0719807371405, 40.3254563203728, 
    38.6615140591414, 42.5623103404995, 41.0797406188206, 39.3063319434942, 
    43.2905509512355, 37.749102414374, 41.5777886205734, 40.0721095592252, 
    38.2719660742721, 42.3176287205335, 40.5778445724771, 39.049165272633, 
    43.0487719903617, 37.2224728843778, 41.3292461440167, 39.5625459179821, 
    43.7712030066013, 38.0110060291271, 42.0719807371405, 40.3254563203728, 
    38.6615140591414, 42.5623103404995, 41.0797406188206, 39.3063319434942, 
    43.2905509512355, 41.5777886205734, 40.0721095592252, 44.0100754561533, 
    38.2719660742721, 42.3176287205335, 40.5778445724771, 39.049165272633, 
    43.0487719903617, 41.3292461440167, 39.5625459179821, 43.7712030066013, 
    42.0719807371405, 40.3254563203728, 38.6615140591414, 42.5623103404995, 
    41.0797406188206, 39.3063319434942, 43.2905509512355, 41.5777886205734, 
    40.0721095592252, 44.0100754561533, 38.2719660742721, 42.3176287205335, 
    40.5778445724771, 39.049165272633, 43.0487719903617, 41.3292461440167, 
    39.5625459179821, 43.7712030066013, 42.0719807371405, 40.3254563203728, 
    44.2479785386593, 38.6615140591414, 42.5623103404995, 41.0797406188206, 
    39.3063319434942, 43.2905509512355, 41.5777886205734, 40.0721095592252, 
    44.0100754561533, 42.3176287205335, 40.5778445724771, 39.049165272633, 
    43.0487719903617, 41.3292461440167, 39.5625459179821, 43.7712030066013, 
    42.0719807371405, 40.3254563203728, 44.2479785386593, 42.5623103404995, 
    41.0797406188206, 39.3063319434942, 43.2905509512355, 41.5777886205734, 
    40.0721095592252, 44.0100754561533, 42.3176287205335, 40.5778445724771, 
    44.7208760649052, 39.049165272633, 43.0487719903617, 41.3292461440167, 
    39.5625459179821, 43.7712030066013, 42.0719807371405, 40.3254563203728, 
    44.2479785386593, 42.5623103404995, 41.0797406188206, 39.3063319434942, 
    43.2905509512354, 41.5777886205734, 40.0721095592252, 44.0100754561533, 
    42.3176287205335, 40.5778445724771, 44.7208760649052, 43.0487719903617, 
    41.3292461440167, 39.5625459179821, 43.7712030066013, 42.0719807371405, 
    40.3254563203728, 44.2479785386593, 42.5623103404995, 41.0797406188206, 
    44.9558704066931, 39.3063319434942, 43.2905509512355, 41.5777886205734, 
    40.0721095592252, 44.0100754561533, 42.3176287205335, 40.5778445724771, 
    44.7208760649052, 43.0487719903617, 41.3292461440167, 39.5625459179821, 
    43.7712030066013, 42.0719807371405, 40.3254563203728, 44.2479785386593, 
    42.5623103404995, 41.0797406188206, 44.9558704066931, 43.2905509512355, 
    41.5777886205734, 40.0721095592252, 44.0100754561533, 42.3176287205335, 
    40.5778445724771, 44.7208760649052, 43.0487719903617, 41.3292461440167, 
    45.4229504848083, 43.7712030066013, 42.0719807371405, 40.3254563203728, 
    44.2479785386593, 42.5623103404995, 41.0797406188206, 44.9558704066931, 
    43.2905509512355, 41.5777886205734, 44.0100754561533, 42.3176287205335, 
    40.5778445724771, 44.7208760649052, 43.0487719903617, 41.3292461440167, 
    45.4229504848083, 43.7712030066013, 42.0719807371405, 40.3254563203728, 
    44.2479785386593, 42.5623103404995, 41.0797406188206, 44.9558704066931, 
    43.2905509512355, 41.5777886205734, 45.6550365094507, 44.0100754561533, 
    42.3176287205335, 40.5778445724771, 44.7208760649052, 43.0487719903617, 
    41.3292461440167, 45.4229504848083, 43.7712030066013, 42.0719807371405, 
    40.3254563203728, 44.2479785386593, 42.5623103404995, 41.0797406188206, 
    44.9558704066931, 43.2905509512355, 41.5777886205734, 45.6550365094507, 
    44.0100754561533, 42.3176287205335, 40.5778445724771, 44.7208760649052, 
    43.0487719903617, 41.3292461440167, 45.4229504848083, 43.7712030066013, 
    42.0719807371405, 46.0012276067282, 44.2479785386593, 42.5623103404995, 
    41.0797406188206, 44.9558704066931, 43.2905509512354, 41.5777886205734, 
    45.6550365094507, 44.0100754561533, 42.3176287205335, 40.5778445724771, 
    44.7208760649052, 43.0487719903617, 41.3292461440167, 45.4229504848083, 
    43.7712030066013, 42.0719807371405, 46.0012276067282, 44.2479785386593, 
    42.5623103404995, 44.9558704066931, 43.2905509512354, 41.5777886205734, 
    45.6550365094507, 44.0100754561533, 42.3176287205335, 46.3454815789384, 
    44.7208760649052, 43.0487719903617, 41.3292461440167, 45.4229504848084, 
    43.7712030066013, 42.0719807371405, 46.0012276067282, 44.2479785386593, 
    42.5623103404995, 44.9558704066931, 43.2905509512355, 41.5777886205734, 
    45.6550365094507, 44.0100754561533, 42.3176287205335, 46.3454815789384, 
    44.7208760649052, 43.0487719903617, 45.4229504848083, 43.7712030066013, 
    42.0719807371405, 46.0012276067282, 44.2479785386593, 42.5623103404995, 
    46.6873156862054, 44.9558704066931, 43.2905509512355, 41.5777886205734, 
    45.6550365094507, 44.0100754561533, 42.3176287205335, 46.3454815789384, 
    44.7208760649052, 43.0487719903617, 45.4229504848084, 43.7712030066013, 
    42.0719807371405, 46.0012276067282, 44.2479785386593, 42.5623103404995, 
    46.6873156862054, 44.9558704066931, 43.2905509512355, 45.6550365094507, 
    44.0100754561533, 42.3176287205335, 46.3454815789384, 44.7208760649052, 
    43.0487719903617, 45.4229504848083, 43.7712030066013, 42.0719807371405, 
    46.0012276067282, 44.2479785386593, 42.5623103404995, 46.6873156862054, 
    44.9558704066931, 43.2905509512355, 45.6550365094507, 44.0100754561533, 
    42.3176287205335, 46.3454815789384, 44.7208760649052, 43.0487719903617, 
    45.4229504848084, 43.7712030066013, 42.0719807371405, 46.0012276067282, 
    44.2479785386593, 42.5623103404995, 46.6873156862054, 44.9558704066931, 
    43.2905509512354, 45.6550365094507, 44.0100754561533, 42.3176287205335, 
    46.3454815789384, 44.7208760649052, 43.0487719903617, 45.4229504848083, 
    43.7712030066013, 46.0012276067282, 44.2479785386593, 42.5623103404995, 
    46.6873156862054, 44.9558704066931, 43.2905509512355, 45.6550365094507, 
    44.0100754561533, 42.3176287205335, 46.3454815789384, 44.7208760649052, 
    43.0487719903616, 45.4229504848083, 43.7712030066013, 46.0012276067282, 
    44.2479785386593, 42.5623103404995, 46.6873156862054, 44.9558704066931, 
    43.2905509512355, 45.6550365094507, 44.0100754561533, 46.3454815789384, 
    44.7208760649052, 43.0487719903617, 45.4229504848084, 43.7712030066013, 
    46.0012276067282, 44.2479785386593, 42.5623103404995, 46.6873156862054, 
    44.9558704066931, 43.2905509512355, 45.6550365094507, 44.0100754561533, 
    46.3454815789384, 44.7208760649052, 43.0487719903617, 45.4229504848083, 
    43.7712030066013, 46.0012276067282, 44.2479785386593, 46.6873156862054, 
    44.9558704066931, 43.2905509512355, 45.6550365094507, 44.0100754561533, 
    46.3454815789384, 44.7208760649052, 43.0487719903617, 45.4229504848083, 
    43.7712030066013, 46.0012276067282, 44.2479785386593, 46.6873156862054, 
    44.9558704066931, 43.2905509512355, 45.6550365094507, 44.0100754561533, 
    46.3454815789384, 44.7208760649052, 45.4229504848084, 43.7712030066013, 
    46.0012276067282, 44.2479785386593, 46.6873156862054, 44.9558704066931, 
    43.2905509512355, 45.6550365094507, 44.0100754561533, 46.3454815789384, 
    44.7208760649052, 45.4229504848083, 43.7712030066013, 46.0012276067282, 
    44.2479785386593, 46.6873156862054, 44.9558704066931, 43.2905509512355, 
    45.6550365094507, 44.0100754561533, 46.3454815789384, 44.7208760649052, 
    45.4229504848083, 43.7712030066013, 46.0012276067282, 44.2479785386593, 
    46.6873156862054, 44.9558704066931, 45.6550365094507, 44.0100754561533, 
    46.3454815789384, 44.7208760649052, 45.4229504848084, 43.7712030066013, 
    46.0012276067282, 44.2479785386593, 46.6873156862054, 44.9558704066931, 
    45.6550365094507, 44.0100754561533, 46.3454815789384, 44.7208760649052, 
    45.4229504848084, 46.0012276067282, 44.2479785386593, 46.6873156862054, 
    44.9558704066931, 45.6550365094507, 44.0100754561533, 46.3454815789384, 
    44.7208760649052, 45.4229504848083, 46.0012276067282, 44.2479785386593, 
    46.6873156862054, 44.9558704066931, 45.6550365094507, 46.3454815789384, 
    44.7208760649052, 45.4229504848083, 46.0012276067282, 44.2479785386593, 
    46.6873156862054, 44.9558704066931, 45.6550365094507, 46.3454815789384, 
    44.7208760649052, 45.4229504848084, 46.0012276067282, 46.6873156862054, 
    44.9558704066931, 45.6550365094507, 46.3454815789384, 44.7208760649052, 
    45.4229504848083, 46.0012276067282, 46.6873156862054, 44.9558704066931, 
    45.6550365094507, 46.3454815789384, 45.4229504848083, 46.0012276067282, 
    46.6873156862054, 44.9558704066931, 45.6550365094507, 46.3454815789384, 
    45.4229504848083, 46.0012276067282, 46.6873156862054, 44.9558704066931, 
    45.6550365094507, 46.3454815789384, 45.4229504848083, 46.0012276067282, 
    46.6873156862054, 45.6550365094507, 46.3454815789384, 45.4229504848084, 
    46.0012276067282, 46.6873156862054, 45.6550365094507, 46.3454815789384, 
    46.0012276067282, 46.6873156862054, 45.6550365094507, 46.3454815789384, 
    46.0012276067282, 46.6873156862054, 46.3454815789384, 46.6873156862054, 
    46.3454815789384, 46.6873156862054, 46.3454815789384, 46.6873156862054 ;
}
