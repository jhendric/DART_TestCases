netcdf True_State {
dimensions:
	metadatalength = 64 ;
	locationrank = 1 ;
	copy = 1 ;
	time = UNLIMITED ; // (200 currently)
	NMLlinelen = 129 ;
	NMLnlines = 200 ;
	StateVariable = 1 ;
variables:
	int copy(copy) ;
		copy:long_name = "ensemble member or copy" ;
		copy:units = "nondimensional" ;
		copy:valid_range = 1, 1 ;
	char CopyMetaData(copy, metadatalength) ;
		CopyMetaData:long_name = "Metadata for each copy/member" ;
	char inputnml(NMLnlines, NMLlinelen) ;
		inputnml:long_name = "input.nml contents" ;
	double time(time) ;
		time:long_name = "time" ;
		time:axis = "T" ;
		time:cartesian_axis = "T" ;
		time:calendar = "no calendar" ;
		time:units = "days since 0000-00-00 00:00:00" ;
	double loc1d(StateVariable) ;
		loc1d:long_name = "location on unit circle" ;
		loc1d:dimension = 1 ;
		loc1d:units = "nondimensional" ;
		loc1d:valid_range = 0., 1. ;
	int StateVariable(StateVariable) ;
		StateVariable:long_name = "State Variable ID" ;
		StateVariable:units = "indexical" ;
		StateVariable:valid_range = 1, 1 ;
	double state(time, copy, StateVariable) ;
		state:long_name = "model state or fcopy" ;

// global attributes:
		:title = "true state from control" ;
		:assim_model_source = "$URL: https://proxy.subversion.ucar.edu/DAReS/DART/releases/Kodiak/assim_model/assim_model_mod.f90 $" ;
		:assim_model_revision = "$Revision: 4933 $" ;
		:assim_model_revdate = "$Date: 2011-06-01 11:55:44 -0600 (Wed, 01 Jun 2011) $" ;
		:creation_date = "YYYY MM DD HH MM SS = 2012 06 03 13 03 33" ;
		:model_source = "$URL: https://proxy.subversion.ucar.edu/DAReS/DART/releases/Kodiak/models/lorenz_63/model_mod.f90 $" ;
		:model_revision = "$Revision: 4933 $" ;
		:model_revdate = "$Date: 2011-06-01 11:55:44 -0600 (Wed, 01 Jun 2011) $" ;
		:model = "Lorenz_63" ;
		:model_r = 28. ;
		:model_b = 2.6666666666667 ;
		:model_sigma = 10. ;
		:model_deltat = 0.01 ;
data:

 copy = 1 ;

 CopyMetaData =
  "true state                                                      " ;

 inputnml =
  "&perfect_model_obs_nml                                                                                                           ",
  "   start_from_restart    = .false.,                                                                                              ",
  "   output_restart        = .true.,                                                                                               ",
  "   async                 = 2,                                                                                                    ",
  "   init_time_days        = 0,                                                                                                    ",
  "   init_time_seconds     = 0,                                                                                                    ",
  "   first_obs_days        = -1,                                                                                                   ",
  "   first_obs_seconds     = -1,                                                                                                   ",
  "   last_obs_days         = -1,                                                                                                   ",
  "   last_obs_seconds      = -1,                                                                                                   ",
  "   output_interval       = 1,                                                                                                    ",
  "   restart_in_file_name  = \"perfect_ics\",                                                                                        ",
  "   restart_out_file_name = \"perfect_restart\",                                                                                    ",
  "   obs_seq_in_file_name  = \"obs_seq.in\",                                                                                         ",
  "   obs_seq_out_file_name = \"obs_seq.out\",                                                                                        ",
  "   adv_ens_command       = \"./advance_model.ksh\",                                                                                ",
  "   output_timestamps     = .false.,                                                                                              ",
  "   trace_execution       = .false.,                                                                                              ",
  "   output_forward_op_errors = .false.,                                                                                           ",
  "   print_every_nth_obs   = -1,                                                                                                   ",
  "   silence               = .false.,                                                                                              ",
  "  /                                                                                                                              ",
  "                                                                                                                                 ",
  "&filter_nml                                                                                                                      ",
  "   async                    = 2,                                                                                                 ",
  "   adv_ens_command          = \"./advance_model.ksh\",                                                                             ",
  "   ens_size                 = 20,                                                                                                ",
  "   start_from_restart       = .false.,                                                                                           ",
  "   output_restart           = .true.,                                                                                            ",
  "   obs_sequence_in_name     = \"obs_seq.out\",                                                                                     ",
  "   obs_sequence_out_name    = \"obs_seq.final\",                                                                                   ",
  "   restart_in_file_name     = \"perfect_ics\",                                                                                     ",
  "   restart_out_file_name    = \"filter_restart\",                                                                                  ",
  "   init_time_days           = 0,                                                                                                 ",
  "   init_time_seconds        = 0,                                                                                                 ",
  "   first_obs_days           = -1,                                                                                                ",
  "   first_obs_seconds        = -1,                                                                                                ",
  "   last_obs_days            = -1,                                                                                                ",
  "   last_obs_seconds         = -1,                                                                                                ",
  "   num_output_state_members = 20,                                                                                                ",
  "   num_output_obs_members   = 0,                                                                                                 ",
  "   output_interval          = 1,                                                                                                 ",
  "   num_groups               = 1,                                                                                                 ",
  "   input_qc_threshold       =  3.0,                                                                                              ",
  "   outlier_threshold        = -1.0,                                                                                              ",
  "   output_forward_op_errors = .false.,                                                                                           ",
  "   output_timestamps        = .false.,                                                                                           ",
  "   output_inflation         = .true.,                                                                                            ",
  "   trace_execution          = .false.,                                                                                           ",
  "   silence                  = .false.,                                                                                           ",
  "                                                                                                                                 ",
  "   inf_flavor                  = 0,                       0,                                                                     ",
  "   inf_initial_from_restart    = .false.,                 .false.,                                                               ",
  "   inf_sd_initial_from_restart = .false.,                 .false.,                                                               ",
  "   inf_output_restart          = .true.,                  .true.,                                                                ",
  "   inf_deterministic           = .true.,                  .true.,                                                                ",
  "   inf_in_file_name            = \'prior_inflate_ics\',     \'post_inflate_ics\',                                                    ",
  "   inf_out_file_name           = \'prior_inflate_restart\', \'post_inflate_restart\',                                                ",
  "   inf_diag_file_name          = \'prior_inflate_diag\',    \'post_inflate_diag\',                                                   ",
  "   inf_initial                 = 1.0,                     1.0,                                                                   ",
  "   inf_sd_initial              = 0.0,                     0.0,                                                                   ",
  "   inf_damping                 = 1.0,                     1.0,                                                                   ",
  "   inf_lower_bound             = 1.0,                     1.0,                                                                   ",
  "   inf_upper_bound             = 1000000.0,               1000000.0,                                                             ",
  "   inf_sd_lower_bound          = 0.0,                     0.0                                                                    ",
  "/                                                                                                                                ",
  "                                                                                                                                 ",
  "&smoother_nml                                                                                                                    ",
  "   num_lags              = 0,                                                                                                    ",
  "   start_from_restart    = .false.,                                                                                              ",
  "   output_restart        = .false.,                                                                                              ",
  "   restart_in_file_name  = \'smoother_ics\',                                                                                       ",
  "   restart_out_file_name = \'smoother_restart\'  /                                                                                 ",
  "                                                                                                                                 ",
  "&ensemble_manager_nml                                                                                                            ",
  "   single_restart_file_in  = .true.,                                                                                             ",
  "   single_restart_file_out = .true.,                                                                                             ",
  "   perturbation_amplitude  = 0.5  /                                                                                              ",
  "                                                                                                                                 ",
  "&assim_tools_nml                                                                                                                 ",
  "   filter_kind                     = 1,                                                                                          ",
  "   cutoff                          = 0.00001,                                                                                    ",
  "   sort_obs_inc                    = .true.,                                                                                     ",
  "   spread_restoration              = .false.,                                                                                    ",
  "   sampling_error_correction       = .false.,                                                                                    ",
  "   adaptive_localization_threshold = -1,                                                                                         ",
  "   output_localization_diagnostics = .false.,                                                                                    ",
  "   localization_diagnostics_file   = \'localization_diagnostics\',                                                                 ",
  "   print_every_nth_obs             = 0  /                                                                                        ",
  "                                                                                                                                 ",
  "&cov_cutoff_nml                                                                                                                  ",
  "   select_localization = 1  /                                                                                                    ",
  "                                                                                                                                 ",
  "&reg_factor_nml                                                                                                                  ",
  "   select_regression    = 1,                                                                                                     ",
  "   input_reg_file       = \"time_mean_reg\",                                                                                       ",
  "   save_reg_diagnostics = .false.,                                                                                               ",
  "   reg_diagnostics_file = \"reg_diagnostics\"  /                                                                                   ",
  "                                                                                                                                 ",
  "&obs_sequence_nml                                                                                                                ",
  "   write_binary_obs_sequence = .false.  /                                                                                        ",
  "                                                                                                                                 ",
  "&obs_kind_nml                                                                                                                    ",
  "   assimilate_these_obs_types = \'RAW_STATE_VARIABLE\'  /                                                                          ",
  "                                                                                                                                 ",
  "&assim_model_nml                                                                                                                 ",
  "   write_binary_restart_files = .false.,                                                                                         ",
  "   netCDF_large_file_support  = .false.                                                                                          ",
  "  /                                                                                                                              ",
  "                                                                                                                                 ",
  "&model_nml                                                                                                                       ",
  "   sigma  = 10.0,                                                                                                                ",
  "   r      = 28.0,                                                                                                                ",
  "   b      = 2.6666666666667,                                                                                                     ",
  "   deltat = 0.01,                                                                                                                ",
  "   time_step_days = 1,                                                                                                           ",
  "   time_step_seconds = 0  /                                                                                                      ",
  "                                                                                                                                 ",
  "&utilities_nml                                                                                                                   ",
  "   TERMLEVEL = 1,                                                                                                                ",
  "   module_details = .false.,                                                                                                     ",
  "   logfilename = \'dart_log.out\',                                                                                                 ",
  "   nmlfilename = \'dart_log.nml\',                                                                                                 ",
  "   write_nml   = \'terminal\'  /                                                                                                   ",
  "                                                                                                                                 ",
  "&preprocess_nml                                                                                                                  ",
  "    input_obs_def_mod_file = \'../../../obs_def/DEFAULT_obs_def_mod.F90\',                                                         ",
  "   output_obs_def_mod_file = \'../../../obs_def/obs_def_mod.f90\',                                                                 ",
  "   input_obs_kind_mod_file = \'../../../obs_kind/DEFAULT_obs_kind_mod.F90\',                                                       ",
  "  output_obs_kind_mod_file = \'../../../obs_kind/obs_kind_mod.f90\',                                                               ",
  "               input_files = \'../../../obs_def/obs_def_1d_state_mod.f90\'  /                                                      ",
  "                                                                                                                                 ",
  "                                                                                                                                 ",
  "&obs_sequence_tool_nml                                                                                                           ",
  "   num_input_files   = 2,                                                                                                        ",
  "   filename_seq      = \'obs_seq.one\', \'obs_seq.two\',                                                                             ",
  "   filename_out      = \'obs_seq.processed\',                                                                                      ",
  "   first_obs_days    = -1,                                                                                                       ",
  "   first_obs_seconds = -1,                                                                                                       ",
  "   last_obs_days     = -1,                                                                                                       ",
  "   last_obs_seconds  = -1,                                                                                                       ",
  "   print_only        = .false.,                                                                                                  ",
  "   gregorian_cal     = .false.                                                                                                   ",
  "   /                                                                                                                             ",
  "                                                                                                                                 ",
  "# other possible obs tool namelist items:                                                                                        ",
  "#                                                                                                                                ",
  "# keep only the U and V radiosonde winds:                                                                                        ",
  "#   obs_types          = \'RADIOSONDE_U_WIND_COMPONENT\',                                                                          ",
  "#                        \'RADIOSONDE_V_WIND_COMPONENT\',                                                                          ",
  "#   keep_types         = .true.,                                                                                                 ",
  "#                                                                                                                                ",
  "# remove the U and V radiosonde winds:                                                                                           ",
  "#   obs_types          = \'RADIOSONDE_U_WIND_COMPONENT\',                                                                          ",
  "#                        \'RADIOSONDE_V_WIND_COMPONENT\',                                                                          ",
  "#   keep_types         = .false.,                                                                                                ",
  "#                                                                                                                                ",
  "# keep only observations with a DART QC of 0:                                                                                    ",
  "#   qc_metadata        = \'Dart quality control\',                                                                                 ",
  "#   min_qc             = 0,                                                                                                      ",
  "#   max_qc             = 0,                                                                                                      ",
  "#                                                                                                                                ",
  "# keep only radiosonde temp obs between 250 and 300 K:                                                                           ",
  "#   copy_metadata      = \'NCEP BUFR observation\',                                                                                ",
  "#   copy_type          = \'RADIOSONDE_TEMPERATURE\',                                                                               ",
  "#   min_copy           = 250.0,                                                                                                  ",
  "#   max_copy           = 300.0,                                                                                                  ",
  "#                                                                                                                                ",
  "                                                                                                                                 ",
  "                                                                                                                                 ",
  "&restart_file_tool_nml                                                                                                           ",
  "   input_file_name              = \"filter_restart\",                                                                              ",
  "   output_file_name             = \"filter_updated_restart\",                                                                      ",
  "   ens_size                     = 1,                                                                                             ",
  "   single_restart_file_in       = .true.,                                                                                        ",
  "   single_restart_file_out      = .true.,                                                                                        ",
  "   write_binary_restart_files   = .true.,                                                                                        ",
  "   overwrite_data_time          = .false.,                                                                                       ",
  "   new_data_days                = -1,                                                                                            ",
  "   new_data_secs                = -1,                                                                                            ",
  "   input_is_model_advance_file  = .false.,                                                                                       ",
  "   output_is_model_advance_file = .false.,                                                                                       ",
  "   overwrite_advance_time       = .false.,                                                                                       ",
  "   new_advance_days             = -1,                                                                                            ",
  "   new_advance_secs             = -1,                                                                                            ",
  "   gregorian_cal                = .false.                                                                                        ",
  "/                                                                                                                                ",
  "                                                                                                                                 ",
  "&obs_diag_nml                                                                                                                    ",
  "   obs_sequence_name  = \'obs_seq.final\',                                                                                         ",
  "   iskip_days         = 0,                                                                                                       ",
  "   obs_select         = 1,                                                                                                       ",
  "   rat_cri            = 4.0,                                                                                                     ",
  "   input_qc_threshold = 3.0,                                                                                                     ",
  "   bin_width_seconds = 0,                                                                                                        ",
  "   lonlim1   = 0.0, 0.0, 0.5, -1.0,                                                                                              ",
  "   lonlim2   = 1.0, 0.5, 1.5, -1.0,                                                                                              ",
  "   reg_names = \'whole\', \'yin\', \'yang\', \'bogus\',                                                                                  ",
  "   verbose   = .false.  /                                                                                                        ",
  "                                                                                                                                 " ;

 time = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 18, 19, 
    20, 21, 22, 23, 24, 25, 26, 27, 28, 29, 30, 31, 32, 33, 34, 35, 36, 37, 
    38, 39, 40, 41, 42, 43, 44, 45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 
    56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 67, 68, 69, 70, 71, 72, 73, 
    74, 75, 76, 77, 78, 79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 
    92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 106, 107, 
    108, 109, 110, 111, 112, 113, 114, 115, 116, 117, 118, 119, 120, 121, 
    122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 
    136, 137, 138, 139, 140, 141, 142, 143, 144, 145, 146, 147, 148, 149, 
    150, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 
    164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 177, 
    178, 179, 180, 181, 182, 183, 184, 185, 186, 187, 188, 189, 190, 191, 
    192, 193, 194, 195, 196, 197, 198, 199, 200 ;

 loc1d = 0 ;

 StateVariable = 1 ;

 state =
  -77.64109263,
  -78.26319591,
  -78.88378501,
  -79.50144611,
  -80.11477639,
  -80.72238923,
  -81.32291942,
  -81.91502833,
  -82.49740887,
  -83.06879045,
  -83.62794375,
  -84.17368535,
  -84.7048822,
  -85.22045591,
  -85.71938687,
  -86.2007181,
  -86.66355892,
  -87.10708838,
  -87.53055842,
  -87.93329679,
  -88.31470966,
  -88.67428402,
  -89.0115897,
  -89.32628117,
  -89.61809898,
  -89.88687091,
  -90.13251283,
  -90.35502918,
  -90.55451321,
  -90.73114684,
  -90.8852002,
  -91.0170309,
  -91.12708291,
  -91.21588521,
  -91.28405006,
  -91.33227097,
  -91.36132045,
  -91.37204739,
  -91.36537416,
  -91.34229351,
  -91.30386515,
  -91.25121207,
  -91.18551671,
  -91.10801678,
  -91.02000102,
  -90.92280463,
  -90.8178046,
  -90.70641488,
  -90.59008135,
  -90.47027675,
  -90.3484954,
  -90.22624793,
  -90.10505584,
  -89.98644611,
  -89.87194565,
  -89.7630759,
  -89.66134723,
  -89.56825358,
  -89.48526695,
  -89.4138321,
  -89.35536122,
  -89.31122878,
  -89.28276644,
  -89.27125815,
  -89.27793533,
  -89.30397228,
  -89.35048178,
  -89.41851082,
  -89.50903664,
  -89.62296292,
  -89.76111628,
  -89.92424296,
  -90.11300587,
  -90.32798182,
  -90.56965912,
  -90.83843539,
  -91.13461579,
  -91.45841145,
  -91.80993829,
  -92.18921613,
  -92.59616817,
  -93.03062072,
  -93.49230336,
  -93.98084932,
  -94.49579631,
  -95.03658756,
  -95.6025733,
  -96.19301244,
  -96.80707464,
  -97.4438427,
  -98.1023152,
  -98.78140944,
  -99.4799647,
  -100.1967457,
  -100.93044643,
  -101.6796941,
  -102.4430534,
  -103.21903097,
  -104.00608008,
  -104.80260543,
  -105.60696823,
  -106.41749136,
  -107.23246468,
  -108.05015049,
  -108.86878902,
  -109.68660411,
  -110.50180888,
  -111.31261141,
  -112.11722057,
  -112.91385169,
  -113.7007324,
  -114.47610825,
  -115.23824845,
  -115.98545137,
  -116.7160501,
  -117.4284178,
  -118.12097298,
  -118.79218455,
  -119.44057686,
  -120.06473436,
  -120.66330625,
  -121.2350108,
  -121.77863947,
  -122.29306082,
  -122.77722414,
  -123.23016281,
  -123.65099739,
  -124.03893845,
  -124.39328903,
  -124.71344686,
  -124.99890626,
  -125.24925969,
  -125.46419898,
  -125.64351626,
  -125.78710455,
  -125.89495795,
  -125.96717164,
  -126.00394136,
  -126.00556272,
  -125.9724301,
  -125.90503523,
  -125.80396544,
  -125.66990166,
  -125.50361601,
  -125.30596919,
  -125.07790752,
  -124.82045968,
  -124.53473326,
  -124.22191102,
  -123.88324682,
  -123.52006148,
  -123.13373828,
  -122.72571835,
  -122.29749582,
  -121.85061286,
  -121.3866545,
  -120.90724338,
  -120.41403434,
  -119.90870896,
  -119.39296997,
  -118.86853561,
  -118.33713404,
  -117.80049757,
  -117.26035705,
  -116.71843616,
  -116.17644583,
  -115.63607861,
  -115.09900327,
  -114.56685934,
  -114.04125183,
  -113.52374612,
  -113.01586297,
  -112.51907361,
  -112.0347952,
  -111.56438628,
  -111.1091426,
  -110.67029307,
  -110.24899603,
  -109.84633568,
  -109.46331889,
  -109.10087218,
  -108.75983905,
  -108.4409776,
  -108.14495841,
  -107.87236277,
  -107.62368122,
  -107.39931241,
  -107.19956224,
  -107.0246434,
  -106.87467518,
  -106.7496836,
  -106.64960194,
  -106.57427149,
  -106.5234427,
  -106.49677661,
  -106.49384657,
  -106.51414034,
  -106.55706238,
  -106.6219365,
  -106.70800878 ;
}
