netcdf wc13_mod_003 {
dimensions:
	xi_rho = 56 ;
	eta_rho = 55 ;
	record = 2 ;
	state_var = 12 ;
	datum = 6815 ;
	Ninner = 50 ;
	Minner = 51 ;
	Nouter = 1 ;
	Mouter = 2 ;
	three = 3 ;
	iteration = UNLIMITED ; // (52 currently)
variables:
	int outer ;
		outer:long_name = "outer loop counter" ;
	int inner ;
		inner:long_name = "inner loop counter" ;
	int Nobs(state_var) ;
		Nobs:long_name = "Number of usable observations" ;
	double obs_mean(state_var) ;
		obs_mean:long_name = "observations mean" ;
	double obs_std(state_var) ;
		obs_std:long_name = "observations standard deviation" ;
	double model_mean(state_var) ;
		model_mean:long_name = "model mean" ;
	double model_std(state_var) ;
		model_std:long_name = "model standard deviation" ;
	double model_bias(state_var) ;
		model_bias:long_name = "model bias" ;
	double SDE(state_var) ;
		SDE:long_name = "model-observations standard deviation error" ;
	double CC(state_var) ;
		CC:long_name = "model-observations cross-correlation" ;
	double MSE(state_var) ;
		MSE:long_name = "model-observations mean squared error" ;
	int nConvRitz ;
		nConvRitz:long_name = "number of converged Ritz eigenvalues" ;
	double Ritz(Ninner) ;
		Ritz:long_name = "converged Ritz eigenvalues to approximate Hessian" ;
	double cg_beta(Nouter, Minner) ;
		cg_beta:long_name = "conjugate gradient beta coefficient" ;
	double cg_delta(Nouter, Ninner) ;
		cg_delta:long_name = "Lanczos algorithm delta coefficient" ;
	double cg_gamma(Nouter, Ninner) ;
		cg_gamma:long_name = "Lanczos algorithm gamma coefficient" ;
	double cg_Gnorm(Nouter) ;
		cg_Gnorm:long_name = "initial gradient normalization factor" ;
	double cg_QG(Nouter, Minner) ;
		cg_QG:long_name = "Lanczos vector normalization factor" ;
	double cg_Greduc(Nouter, Ninner) ;
		cg_Greduc:long_name = "reduction in the gradient norm" ;
	double cg_Tmatrix(three, Ninner) ;
		cg_Tmatrix:long_name = "Lanczos recurrence tridiagonal matrix" ;
	double cg_zu(Nouter, Ninner) ;
		cg_zu:long_name = "tridiagonal matrix, upper diagonal elements" ;
	double cg_Ritz(Nouter, Ninner) ;
		cg_Ritz:long_name = "Lanczos recurrence eigenvalues" ;
	double cg_RitzErr(Nouter, Ninner) ;
		cg_RitzErr:long_name = "Ritz eigenvalues relative error" ;
	double cg_zv(Ninner, Ninner) ;
		cg_zv:long_name = "Lanczos recurrence eigenvectors" ;
	double obs_scale(datum) ;
		obs_scale:long_name = "observation screening/normalization scale" ;
	double NLmodel_initial(datum) ;
		NLmodel_initial:long_name = "initial nonlinear model at observation locations" ;
	double NLmodel_value(datum) ;
		NLmodel_value:long_name = "nonlinear model at observation locations" ;
	double TLmodel_value(datum) ;
		TLmodel_value:long_name = "tangent linear model at observation locations" ;
	double misfit_initial(datum) ;
		misfit_initial:long_name = "initial model-observation misfit" ;
	double misfit_final(datum) ;
		misfit_final:long_name = "final model-observation misfit" ;
	double NLcost_function(Mouter, state_var) ;
		NLcost_function:long_name = "nonlinear model misfit cost function" ;
	double TLcost_function(iteration) ;
		TLcost_function:long_name = "tangent linear model misfit cost function" ;
	double back_function(iteration) ;
		back_function:long_name = "model minus background misfit cost function" ;
	double Jmin(iteration) ;
		Jmin:long_name = "normalized, optimal cost function minimum" ;
	double zeta_ref(eta_rho, xi_rho) ;
		zeta_ref:long_name = "reference free-surface, balance operator" ;
		zeta_ref:units = "meter" ;
	double obs_depth(datum) ;
		obs_depth:long_name = "depth of observation" ;
		obs_depth:units = "meter" ;
		obs_depth:negative = "downwards" ;
	double obs_Xgrid(datum) ;
		obs_Xgrid:long_name = "observation fractional x-grid location" ;
	double obs_Ygrid(datum) ;
		obs_Ygrid:long_name = "observation fractional y-grid location" ;
	double obs_Zgrid(datum) ;
		obs_Zgrid:long_name = "observation fractional z-grid location" ;
	double obs_lon(datum) ;
		obs_lon:long_name = "observation longitude" ;
	double obs_lat(datum) ;
		obs_lat:long_name = "observation latitude" ;
	int obs_type(datum) ;
		obs_type:long_name = "model state variable associated with observation" ;
		obs_type:flag_values = 1, 2, 3, 4, 5, 6, 7 ;
		obs_type:flag_meanings = "zeta ubar vbar u v temperature salinity" ;
	double obs_error(datum) ;
		obs_error:long_name = "observation error covariance" ;
	double obs_value(datum) ;
		obs_value:long_name = "observation value" ;
	double obs_time(datum) ;
		obs_time:long_name = "time of observation" ;
		obs_time:units = "days since 1968-05-23 00:00:00 GMT" ;
		obs_time:calendar = "gregorian" ;
	int obs_provenance(datum) ;
		obs_provenance:long_name = "observation origin" ;
		obs_provenance:flag_values = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11 ;
		obs_provenance:flag_meanings = "gridded_AVISO_SLA blended_SST XBT_Met_Office CTD_temperature_Met_Office CTD_salinity_Met_Office ARGO_temperature_Met_Office ARGO_salinity_Met_Office CTD_temperature_CalCOFI CTD_salinity_CalCOFI CTD_temperature_GLOBEC CTD_salinity_GLOBEC" ;

// global attributes:
		:type = "ROMS observations" ;
		:obs_file = "wc13_obs.nc" ;
		:svn_url = "https:://myroms.org/svn/src" ;
		:svn_rev = "670" ;
		:code_dir = "/Users/arango/ocean/repository/trunk" ;
		:header_dir = "/Users/arango/ocean/repository/Projects/wc13/I4DVAR" ;
		:header_file = "wc13.h" ;
		:os = "Darwin" ;
		:cpu = "x86_64" ;
		:compiler_system = "ifort" ;
		:compiler_command = "/opt/intelsoft/openmpi/bin/mpif90" ;
		:compiler_flags = "-heap-arrays -fp-model source -ip -O3 -free -free" ;
		:history = "Mon Sep 12 12:04:05 2016: ncks -a -v obs_provenance wc13_obs.nc wc13_mod_003.nc\n",
			"4D-Var observations, Monday - June 21, 2010 - 11:00:00 AM" ;
		:title = "California Current System, 1/3 degree resolution (WC13)" ;
		:Conventions = "CF-1.4" ;
		:grd_file = "wc13_grd.nc" ;
		:state_variables = "\n",
			"1: free-surface (m) \n",
			"2: vertically integrated u-momentum component (m/s) \n",
			"3: vertically integrated v-momentum component (m/s) \n",
			"4: u-momentum component (m/s) \n",
			"5: v-momentum component (m/s) \n",
			"6: potential temperature (Celsius) \n",
			"7: salinity (nondimensional)" ;
		:obs_provenance = "\n",
			" 1: gridded AVISO sea level anomaly \n",
			" 2: blended satellite SST \n",
			" 3: XBT temperature from Met Office \n",
			" 4: CTD temperature from Met Office \n",
			" 5: CTD salinity from Met Office \n",
			" 6: ARGO floats temperature from Met Office \n",
			" 7: ARGO floats salinity from Met Office \n",
			" 8: CTD temperature from CalCOFI \n",
			" 9: CTD salinity from CalCOFI \n",
			"10: CTD temperature from GLOBEC \n",
			"11: CTD salinity from GLOBEC " ;
		:variance_units = "squared state variable units" ;
		:obs_sources = "\n",
			"http://opendap.aviso.oceanobs.com/thredds/dodsC \n",
			"http://hadobs.metoffice.com/en3" ;
		:grid_Lm_Mm_N = 54, 53, 30 ;
		:NCO = "\"4.5.5\"" ;
data:

 outer = 1 ;

 inner = 50 ;

 Nobs = 0, 1570, 0, 0, 0, 0, 5120, 125, 0, 0, 0, 0 ;

 obs_mean = 0, 0.00258845199373017, 0, 0, 0, 0, 13.2088473930503, 
    33.677364956665, 0, 0, 0, 0 ;

 obs_std = 0, 0.105560808827345, 0, 0, 0, 0, 2.61113085351517, 
    0.675098577590138, 0, 0, 0, 0 ;

 model_mean = 0, 0.00137164941748997, 0, 0, 0, 0, 13.3050108564258, 
    33.6603444833008, 0, 0, 0, 0 ;

 model_std = 0, 0.103785555259157, 0, 0, 0, 0, 2.67971230432661, 
    0.67065635001406, 0, 0, 0, 0 ;

 model_bias = 0, -0.0012168025762402, 0, 0, 0, 0, 0.0961634633754809, 
    -0.0170204733641981, 0, 0, 0, 0 ;

 SDE = 0, -0.00177525356818758, 0, 0, 0, 0, 0.0685814508114366, 
    -0.00444222757607815, 0, 0, 0, 0 ;

 CC = 0, 0.989843420607303, 0, 0, 0, 0, 0.996752811419038, 0.986571659914458, 
    0, 0, 0, 0 ;

 MSE = 0, 0.000227176746579411, 0, 0, 0, 0, 0.0593925002352884, 
    0.0124690375303049, 0, 0, 0, 0 ;

 nConvRitz = 50 ;

 Ritz = 1505.24607252525, 546.151572927295, 516.357734165814, 
    461.351128003063, 333.85113022939, 262.703265545834, 245.926411213377, 
    236.12879548758, 220.670394450501, 175.937851990562, 170.645230681192, 
    154.759555304143, 139.749552457334, 133.035656878016, 126.432911762351, 
    114.704238057692, 112.012250636493, 110.422359462562, 108.980613214424, 
    100.177016394331, 95.0554514279069, 91.5251303367642, 89.4948199641041, 
    85.2102229400014, 80.0849482850984, 76.8186118922852, 73.2715327224884, 
    69.7571527665927, 64.4434435599309, 59.8955030097135, 54.6543085077524, 
    50.7587073215926, 46.3374115756665, 41.2391098020417, 37.5941435527002, 
    33.4319883394266, 29.9114835046698, 26.4276184285484, 22.7732931831815, 
    19.3141616473858, 15.8811832634076, 13.3891650050172, 10.7025920656435, 
    8.5733680364005, 6.43241429571385, 4.81573277963173, 3.48622962181792, 
    2.39966044479215, 1.60583364004856, 1.15928814696021 ;

 cg_beta =
  0, 576.837751159746, 275.801247344185, 158.284392743192, 105.936785250829, 
    179.076602914418, 105.905861433906, 146.599033398814, 150.903151472083, 
    114.942531598984, 69.8235908459163, 80.7945683150605, 59.8215760011393, 
    53.4609376048075, 71.8816636833254, 68.6314588970497, 41.6363677723498, 
    58.088430512528, 64.725164630219, 55.3914187593564, 41.2396586414287, 
    37.5208128922219, 52.3670201707217, 46.7400455627169, 40.8691375091857, 
    29.8597836877664, 32.8029387993208, 31.4466906806959, 34.1459872768881, 
    36.0188495846866, 35.1637390441155, 28.8568714435612, 30.437706157788, 
    27.5882280133829, 28.9358784329294, 27.9925918178509, 31.7671032336367, 
    24.0859695854857, 22.5581006777668, 29.7623453066221, 31.4196038214026, 
    27.1921229016679, 23.5007829190996, 25.001159678048, 22.9284246074192, 
    22.3901459707751, 23.5218961790355, 25.7892733638672, 24.7741854591191, 
    23.0646233208797, 21.6211096382363 ;

 cg_delta =
  648.455702585648, 1048.87486669404, 366.755691632265, 247.900653431853, 
    295.710672020189, 267.578261566505, 265.214755844329, 284.328324005431, 
    319.121939435475, 152.404740319681, 153.6411558921, 151.676715312983, 
    96.0900471720125, 142.304001036243, 146.378388825422, 109.116176923155, 
    88.729079180642, 133.491492765953, 122.710297487985, 103.6605733136, 
    67.6540200024351, 101.238075961611, 95.7005496379107, 90.1769862502786, 
    73.5840240759833, 59.427086735909, 66.2296147845909, 67.0645127805779, 
    70.1836655430713, 73.8857972575818, 66.9394829730371, 58.5492234266743, 
    59.3628675534845, 53.8491702769334, 60.9057752082868, 65.170579664961, 
    53.2644297874145, 48.3078879204786, 52.5200830738014, 62.7179106214527, 
    61.4138096008519, 47.2904879848836, 54.1703261477972, 47.1970368567157, 
    44.353082809126, 49.1940450656104, 53.8576353178948, 45.9693120557287, 
    53.5310509107858, 43.8361857231055 ;

 cg_gamma =
  0, 0.889556139085009, 0.51479918785962, 0.704195288056908, 
    0.776449011770444, 0.838938558064992, 0.90252476792022, 
    0.864217560198006, 0.957295528748782, 0.658081640997541, 
    0.909597537294562, 0.896424685572296, 0.754841909967597, 
    1.04960757997866, 0.833981126508448, 0.794065846567615, 
    0.762315624364336, 1.01929152178252, 0.871338604825092, 
    0.835305548817532, 0.718563430265042, 0.986851993521043, 
    0.815551183218814, 0.882011393731575, 0.834886419132214, 
    0.756653877208857, 0.890571907252746, 0.849537703392981, 
    0.846258389210621, 0.872394586201918, 0.828100148029078, 
    0.762997814234327, 0.833190848962617, 0.811360021574699, 
    0.919615709623364, 0.816208426302611, 0.750590945718469, 
    0.818684556146157, 0.789046144881428, 0.85719310694088, 
    0.844480581902345, 0.779578067641029, 0.900685575062822, 
    0.757530326346009, 0.811398739454877, 0.869554406714387, 
    0.791327727189469, 0.731732927760743, 0.914228822678169, 0.746868410132881 ;

 cg_Gnorm = 1618.27470777448 ;

 cg_QG =
  1618.27470777447, -4.96323413504364e-12, -2.47038803101719e-12, 
    -2.13351693587849e-12, -5.38993752221933e-13, 5.21027293814536e-12, 
    -8.75864847360642e-13, 4.94077606203439e-13, -6.17597007754299e-13, 
    -2.24580730092472e-13, 1.32502630754559e-12, 5.83909898240428e-13, 
    3.12167214828536e-12, -8.53406774351395e-13, 1.89770716928139e-12, 
    -6.73742190277417e-13, 1.34748438055483e-13, 5.44608270474245e-13, 
    -8.49195885662161e-13, 4.88463087951127e-13, 2.08860078985999e-12, 
    -1.45977474560107e-13, 5.7548812086196e-13, 5.22150197464998e-13, 
    1.12290365046236e-13, -4.32317905428009e-13, -1.15659075997623e-12, 
    -6.59705894646637e-13, 1.17904883298548e-12, 3.93016277661826e-14, 
    1.03868587667768e-13, -4.63197755815724e-14, -2.21773470966316e-13, 
    -9.1797373425298e-13, -4.37581516289551e-13, 3.565219090218e-13, 
    -1.66751192093661e-12, -8.02876110080588e-13, -1.62821029317042e-12, 
    -1.79664584073978e-13, -6.17597007754299e-13, 2.97569467372526e-13, 
    1.03868587667768e-12, 1.56645059239499e-12, -1.31379727104096e-12, 
    -2.89147689994058e-13, 2.10544434461693e-13, -1.13693994609314e-13, 
    -1.29695371628403e-12, -7.01814781538976e-14, _ ;

 cg_Greduc =
  0, 0.457942777956499, 0.322481146436659, 0.250390167465343, 
    0.210061966047025, 0.189586127155454, 0.163843660257676, 
    0.156846803378509, 0.103218001752547, 0.0938868401985816, 
    0.0841624812043912, 0.0635293680599342, 0.0666809062669636, 
    0.055610617325127, 0.0441584919244249, 0.0336627083423559, 
    0.0343121132136013, 0.0298974688561397, 0.0249735216311328, 
    0.0179450593690645, 0.0177091176122163, 0.0144426918224042, 
    0.0127386187435146, 0.0106352997874632, 0.00804724081946265, 
    0.00716664660471112, 0.00608833649759486, 0.00515230583742715, 
    0.00449484371902864, 0.0037221807490952, 0.00284001577574476, 
    0.00236627515526001, 0.00191990106102333, 0.00176557117664016, 
    0.00144107407161048, 0.00108165715026031, 0.000885536003962333, 
    0.000698728770080577, 0.000598945485333489, 0.000505797831982301, 
    0.000394308896473489, 0.000355148335172443, 0.000269035634244906, 
    0.000218295174493976, 0.000189819530945018, 0.000150209457999034, 
    0.000109913206479081, 0.000100485821356217, 7.5049685636619e-05, 
    6.09793574901997e-05 ;

 cg_Tmatrix =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -10.5596904652389, 9.06531651480074, -12.3899169528596, 12.9124983426287, 
    -11.7040203987472, 11.6882671404991, -9.74082052460109, 9.17845981501693, 
    -7.83085847584655, 9.69127978142432, -8.26222589896967, 7.33635930594332, 
    -7.44232995540063, 5.16753489686511, -4.69503537682502, 4.60139873878265, 
    -4.31977910209719, 3.30021813545707, -2.92964657930371, 2.63381304208387, 
    -2.68540752034428, 1.94721429743659, -1.8403482866321, 1.58648823022219, 
    -1.39583969790655, 1.26836472411655, -1.02721738551218, 
    0.840346654928525, -0.704470818209913, 0.576028339104788, 
    -0.488744516567275, 0.431820721487277, -0.367278998008152, 
    0.313869461868315, -0.233932188061603, 0.184539277436195, 
    -0.172447685510225, 0.137966186002716, -0.11132521207438, 
    0.0918796635213896, -0.0779513686899032, 0.069890383131717, 
    -0.0504445800832075, 0.043602802726826, -0.0347494474411256, 
    0.0241848153040863, -0.0175029976422037, 0.0144942955165003, 
    -0.00867448106814825, 0.00456412060129481 ;

 cg_zu =
  -10.5596904652389, 9.06531651480074, -12.3899169528596, 12.9124983426287, 
    -11.7040203987472, 11.6882671404991, -9.74082052460109, 9.17845981501693, 
    -7.83085847584655, 9.69127978142432, -8.26222589896967, 7.33635930594332, 
    -7.44232995540063, 5.16753489686511, -4.69503537682502, 4.60139873878265, 
    -4.31977910209719, 3.30021813545707, -2.92964657930371, 2.63381304208387, 
    -2.68540752034428, 1.94721429743659, -1.8403482866321, 1.58648823022219, 
    -1.39583969790655, 1.26836472411655, -1.02721738551218, 
    0.840346654928525, -0.704470818209913, 0.576028339104788, 
    -0.488744516567275, 0.431820721487277, -0.367278998008152, 
    0.313869461868315, -0.233932188061603, 0.184539277436195, 
    -0.172447685510225, 0.137966186002716, -0.11132521207438, 
    0.0918796635213896, -0.0779513686899032, 0.069890383131717, 
    -0.0504445800832075, 0.043602802726826, -0.0347494474411256, 
    0.0241848153040863, -0.0175029976422037, 0.0144942955165003, 
    -0.00867448106814825, 0.00456412060129481 ;

 cg_Ritz =
  1.15928814696021, 1.60583364004856, 2.39966044479215, 3.48622962181792, 
    4.81573277963173, 6.43241429571385, 8.5733680364005, 10.7025920656435, 
    13.3891650050172, 15.8811832634076, 19.3141616473858, 22.7732931831815, 
    26.4276184285484, 29.9114835046698, 33.4319883394266, 37.5941435527002, 
    41.2391098020417, 46.3374115756665, 50.7587073215926, 54.6543085077524, 
    59.8955030097135, 64.4434435599309, 69.7571527665927, 73.2715327224884, 
    76.8186118922852, 80.0849482850984, 85.2102229400014, 89.4948199641041, 
    91.5251303367642, 95.0554514279069, 100.177016394331, 108.980613214424, 
    110.422359462562, 112.012250636493, 114.704238057692, 126.432911762351, 
    133.035656878016, 139.749552457334, 154.759555304143, 170.645230681192, 
    175.937851990562, 220.670394450501, 236.12879548758, 245.926411213377, 
    262.703265545834, 333.85113022939, 461.351128003063, 516.357734165814, 
    546.151572927295, 1505.24607252525 ;

 cg_RitzErr =
  0.000269181084218068, 0.000552403979973174, 0.00074122397342458, 
    0.00109105844780257, 0.00164507539687702, 0.00159617122611334, 
    0.0020304800349127, 0.00206578233886586, 0.0022677116062269, 
    0.00175390784701051, 0.00191072785996881, 0.00345499525056285, 
    0.00337664950458708, 0.00498414690698201, 0.00378427380658216, 
    0.00287174725948031, 0.00508369845495238, 0.00284582259659401, 
    0.00258781636701397, 0.00255744910207239, 0.0038371607059645, 
    0.00197617980918838, 0.0024448709569464, 0.00230379356997206, 
    0.00337727880883166, 0.00303022078304318, 0.000934833588558271, 
    0.00186351465168619, 0.000761511715807037, 0.00230875194343324, 
    3.37106362059995e-05, 8.61261185027899e-06, 6.19942999606347e-06, 
    2.40840556255953e-06, 4.2420425061803e-07, 2.95843229762714e-10, 
    5.05938474400834e-11, 3.2490551875589e-13, 4.58433337157568e-16, 
    2.77365345298856e-18, 1.97817224807635e-18, 3.53825767912769e-24, 
    1.74679564923476e-26, 2.25586114945351e-27, 2.00788680917567e-29, 
    2.05829888617399e-36, 2.49786867747715e-44, 1.04498045623343e-46, 
    3.79187648920381e-48, 0 ;

 cg_zv =
  -0.00854294546546421, 0.00958643562669468, -0.0185494610612244, 
    0.0261407032963783, -0.0331698062457375, 0.0390947234152111, 
    -0.0422605490950909, 0.047877319058097, -0.0487863809145711, 
    0.0721004538283593, -0.0758659866540688, 0.080870222982627, 
    -0.10101402637839, 0.0888789875145329, -0.0993924492994279, 
    0.117219023779258, -0.140097530738366, 0.127180869614152, 
    -0.134292113921806, 0.14607929263011, -0.182704822511036, 
    0.163233350954291, -0.181048346909502, 0.183322348589075, 
    -0.192241040000491, 0.215365936706274, -0.20756137717565, 
    0.204837165040577, -0.204203231655576, 0.1971366042465, 
    -0.198553730315815, 0.212387644580201, -0.212212893863322, 
    0.213386568319268, -0.186230234622776, 0.176906609271286, 
    -0.192367354072018, 0.18282501336969, -0.176725390203877, 
    0.166403938116994, -0.15862183194438, 0.159212900796559, 
    -0.128992204418796, 0.123849568203639, -0.108023147742634, 
    0.0815650857087457, -0.0637408229114025, 0.0558554138593565, 
    -0.0346753246595929, 0.0187401931074241,
  -0.0154317539978226, 0.0173047412916771, -0.0334338640453009, 
    0.046976845576454, -0.0592626520930049, 0.0695392726438352, 
    -0.0744337910864916, 0.0836076104111285, -0.0843311082591823, 
    0.123190545717056, -0.127231619341167, 0.132955645546154, 
    -0.161699972425094, 0.137006173031405, -0.147908169986249, 
    0.168505991788206, -0.191298712150169, 0.166136133119293, 
    -0.166839768348059, 0.170637480296256, -0.198179917708956, 
    0.161307611235873, -0.164904693287079, 0.15125063027156, 
    -0.139195249157223, 0.128518658568476, -0.0998315996765723, 
    0.0710951044075452, -0.0443512785384524, 0.0170439089760952, 
    0.0103956211657058, -0.044305268430308, 0.0730313596809792, 
    -0.104012623598841, 0.118163362970954, -0.142801492400172, 
    0.181616868446976, -0.201182796169352, 0.222591058045665, 
    -0.22830038461133, 0.233200863676684, -0.249122293119539, 
    0.214454102326581, -0.216714032223401, 0.197076436976791, 
    -0.154334152716432, 0.124646247735634, -0.111781323142422, 
    0.0704149148616435, -0.0384579670153214,
  0.0253086642447348, -0.0283456057114005, 0.0546189720328165, 
    -0.0763372702518428, 0.0952978212843987, -0.110930043530298, 
    0.116619264484125, -0.128931009049854, 0.127585643083527, 
    -0.182292139944421, 0.181596650180933, -0.182396632038605, 
    0.209884291405688, -0.163724895897283, 0.16256179939468, 
    -0.169552322559434, 0.166613471398412, -0.126085370460591, 
    0.10583900753178, -0.0825518132963771, 0.0605412185345025, 
    -0.0145564501308535, -0.0159035068961719, 0.0480549221824009, 
    -0.0850226389839241, 0.136917241946544, -0.160634397628289, 
    0.183230674934184, -0.199061877109917, 0.200911996948676, 
    -0.204541464788851, 0.212644423966949, -0.198354787009594, 
    0.174948398943515, -0.121950757022095, 0.0740402816377607, 
    -0.0388407707637166, -0.0156281200518909, 0.0732764223931499, 
    -0.11155386174533, 0.144745795672021, -0.185240109899858, 
    0.186361295991096, -0.211780605869898, 0.210566887245078, 
    -0.177676639836421, 0.153033822325062, -0.143296751952826, 
    0.0927077294022395, -0.0516034788929513,
  -0.0308865826538425, 0.0345346726975672, -0.0662999450512769, 
    0.0919865775213242, -0.113167487321778, 0.130254556942559, 
    -0.133453816736021, 0.144161589775975, -0.13864814658522, 
    0.191468446337477, -0.180120024648292, 0.169279876718456, 
    -0.176072718513654, 0.115568809060187, -0.0922348142858177, 
    0.0709930049600992, -0.0280710727111246, -0.00969268115433617, 
    0.04466120923985, -0.0848024976284051, 0.146004768186825, 
    -0.156488542034333, 0.187500191806939, -0.194594676656033, 
    0.198335290175521, -0.199262990888902, 0.159275169554604, 
    -0.109933717675874, 0.058007402888408, -0.00319692920163267, 
    -0.0530176123631192, 0.120475845080502, -0.167681436328917, 
    0.206699267933227, -0.199888497552609, 0.196354872893061, 
    -0.205137545693452, 0.164982035673622, -0.108778295523141, 
    0.0541670225945215, 0.000925962987063615, -0.0645607991492231, 
    0.119266623429553, -0.181099268459819, 0.215199753227165, 
    -0.207332984956823, 0.198044574669025, -0.19771470866878, 
    0.132884473551495, -0.0759587029032932,
  -0.0303688063643807, 0.0338857461601913, -0.0647598551181621, 
    0.0890387737814856, -0.10755007234882, 0.12203319667944, 
    -0.120919178434717, 0.126625699269222, -0.117074046951757, 
    0.153893274074447, -0.132565056228479, 0.111191504176207, 
    -0.0939319462417746, 0.0359500424255403, 0.00109876199636037, 
    -0.0399189026377915, 0.0981869902390422, -0.113226003090015, 
    0.136977849167912, -0.159237160005484, 0.197682874989139, 
    -0.156051180787558, 0.145694720045436, -0.108461653289967, 
    0.0599142769922409, 0.0104666454732763, -0.0719638275678536, 
    0.129623855348493, -0.170031769228337, 0.185694180135597, 
    -0.190581560916617, 0.184009538246008, -0.144159588658809, 
    0.0820155703749938, -0.00153434918715133, -0.0817048624097747, 
    0.156584465207511, -0.207207208096389, 0.232306764170405, 
    -0.215300310720708, 0.176716510494759, -0.11904786480986, 
    0.010690360582632, 0.0907997731944095, -0.179492672535955, 
    0.223972138201789, -0.251707528536315, 0.274376350237146, 
    -0.193758726305054, 0.114528963665116,
  0.0384211360860856, -0.0427629157076312, 0.0812727179478381, 
    -0.110499754863087, 0.130436074608882, -0.145336304031382, 
    0.137819785604024, -0.138291228013225, 0.120781568065525, 
    -0.147017372949997, 0.108523904309356, -0.0706778513641783, 
    0.0250313217796981, 0.0371076806230267, -0.0887580650115327, 
    0.142121007531384, -0.204194668410792, 0.187423512112112, 
    -0.18466559326496, 0.168645375321538, -0.149569379708994, 
    0.0586874246821962, 0.000917840691470845, -0.0675056996881896, 
    0.137275615563975, -0.216323698558282, 0.224522058979511, 
    -0.201284694615224, 0.150642523409069, -0.075809882006466, 
    -0.00888237135592622, 0.111003203093446, -0.181643625559469, 
    0.226031064803835, -0.197209637097883, 0.150120587303437, 
    -0.103799171875349, 0.00382912677034972, 0.103721374114473, 
    -0.163517159432546, 0.194676328801987, -0.204689124242741, 
    0.130614400099738, -0.0569935179885239, -0.0410927588812747, 
    0.127959704768761, -0.193508752202977, 0.23914363019327, 
    -0.180209644244967, 0.111124290537612,
  0.0391660366796678, -0.0434466276439782, 0.0819617153554837, 
    -0.109768267443853, 0.125520904709179, -0.136328456084863, 
    0.121163076996711, -0.113626108342592, 0.0899290200318348, 
    -0.0937928781437675, 0.0451665276582698, -4.02589531075943e-05, 
    -0.0609052645724882, 0.099748247789869, -0.140276994879701, 
    0.177189941615959, -0.196649229179354, 0.144349109834297, 
    -0.102105186755568, 0.0417204081583539, 0.040947820566623, 
    -0.110332346433626, 0.165896763169421, -0.185629712083827, 
    0.180919743734081, -0.139826364630762, 0.0520827176922717, 
    0.0503652888316379, -0.134239858846168, 0.18187102599493, 
    -0.200299325955965, 0.183506662981895, -0.111404273877058, 
    0.00263320385801926, 0.102095607676074, -0.193590611878764, 
    0.254941978756116, -0.217712421511137, 0.111275937235076, 
    0.000704474692536396, -0.106620578265107, 0.206373887759218, 
    -0.216629493413141, 0.201098591633195, -0.102544195160924, 
    -0.0420663556053946, 0.170255973943151, -0.260590381369494, 
    0.216121957618056, -0.141360556836925,
  0.0472432247050738, -0.0522322151178216, 0.0978036261296416, 
    -0.128992971432094, 0.142689766805329, -0.150788184014107, 
    0.124463526690829, -0.107150290171475, 0.0733771545619173, 
    -0.0562160721878104, -0.00670572375020258, 0.06044607512021, 
    -0.133389103423567, 0.145410405274774, -0.167012101037979, 
    0.17786534375069, -0.145115490999519, 0.0674348590199332, 
    0.00230635036823577, -0.0834616889776982, 0.185032523334062, 
    -0.189119965922064, 0.194387553635164, -0.141610815450537, 
    0.0530657309247953, 0.0820723540342798, -0.170212347665711, 
    0.214940597661231, -0.198027657595393, 0.123255983746212, 
    -0.0186265658157996, -0.113894574633397, 0.19669603585273, 
    -0.221275309648057, 0.142410653855738, -0.0266739386497983, 
    -0.0797544404871029, 0.176112873566639, -0.208431275026312, 
    0.159372555751151, -0.0664047417108327, -0.0603100120343153, 
    0.170730581822158, -0.240146421485477, 0.196068760047248, 
    -0.0487549691149668, -0.106851868422209, 0.223271367278848, 
    -0.206602826796966, 0.143818277798786,
  0.0521904317766691, -0.0574587858312147, 0.106570728557456, 
    -0.137798319905992, 0.145811542358786, -0.148360103568806, 
    0.109532039714721, -0.080974381419166, 0.0389775799678852, 
    0.00263232135467151, -0.0694051297839652, 0.118206083650226, 
    -0.179515033832232, 0.145429126229643, -0.127305483350293, 
    0.0943673642017876, -0.00711744961336181, -0.0584089845199233, 
    0.114769835236837, -0.158259842776783, 0.192268198690754, 
    -0.104124184116962, 0.0369151627191377, 0.0516502511601693, 
    -0.139262215639572, 0.210047343037358, -0.168027734873959, 
    0.063233710909658, 0.055345442637805, -0.147214425807692, 
    0.196580283971484, -0.185409117227067, 0.088718728309538, 
    0.0567162125306612, -0.16389102458551, 0.219572826270455, 
    -0.213493089421937, 0.0638504846158885, 0.129115953502178, 
    -0.218153891814146, 0.220195782261807, -0.136823275813426, 
    -0.0574066282737012, 0.222252212818102, -0.265113811949152, 
    0.139037466774845, 0.0407159830703481, -0.190704807430003, 
    0.208408670395531, -0.157876447879269,
  0.0709925877162254, -0.077852224407547, 0.14310903879824, 
    -0.181581851079803, 0.183870008244824, -0.179900960355839, 
    0.116648214592605, -0.068429850236443, 0.00841123673046339, 
    0.0676481556547051, -0.146116456606605, 0.190675713010037, 
    -0.235491854337055, 0.139952884740122, -0.0710003421124664, 
    -0.0115792373577378, 0.142962691067268, -0.170987815751431, 
    0.182393535083158, -0.151968038687008, 0.0784833136088946, 
    0.058735568016046, -0.151970520297888, 0.19371791049276, 
    -0.17835753613462, 0.079526784862523, 0.0567830755151576, 
    -0.173870475001861, 0.208329896746559, -0.149251060518315, 
    0.032802169792903, 0.123831938424103, -0.204688030256326, 
    0.185985854269875, -0.0488849319910961, -0.113624346575048, 
    0.21937446909217, -0.190626061174156, 0.0397874009017797, 
    0.0955030678910924, -0.180053750814965, 0.191145487920977, 
    -0.047134734148712, -0.107487815827922, 0.198203574653596, 
    -0.14196897107602, 0.0123963537213825, 0.111232675115354, 
    -0.147995824753605, 0.12210580041715,
  0.0655060932074122, -0.071445747679478, 0.129699728354759, 
    -0.160206861152163, 0.151898904340766, -0.13967501525371, 
    0.070579211255931, -0.0174835202874377, -0.0378617915423852, 
    0.12170932465979, -0.16966234670132, 0.176893710552208, 
    -0.162254287563991, 0.0350752557284324, 0.0606603416167105, 
    -0.149042834410745, 0.221468385536575, -0.157821572557523, 
    0.0796428259864688, 0.0357504258947172, -0.180092404006767, 
    0.192727859097708, -0.172471284239425, 0.0659364943530451, 
    0.0829200138755042, -0.240953701320247, 0.219168902430815, 
    -0.075633359242717, -0.0960762151565427, 0.207389331134396, 
    -0.223440978670153, 0.116050837059389, 0.0622433840882614, 
    -0.218393448785742, 0.201308385345984, -0.0733527748565708, 
    -0.0715031501998471, 0.197532271914476, -0.177540386853481, 
    0.0483644431945046, 0.101364109039158, -0.212818431676197, 
    0.136062385470492, 0.0103509947962491, -0.160950130011376, 
    0.169390839053908, -0.0619712631575721, -0.0714906157564379, 
    0.14142894699119, -0.133023496712505,
  -0.0444324586023138, 0.0481948480280239, -0.0863755698257805, 
    0.103734020706802, -0.0913890449767703, 0.0779232880703256, 
    -0.0255922412381225, -0.013969481945571, 0.0490750924458509, 
    -0.108187093045765, 0.120068790035936, -0.100986177419694, 
    0.0554408295441355, 0.0369692473701567, -0.102708794672489, 
    0.146258283650393, -0.1340008233141, 0.0473152039729345, 
    0.0393238600700202, -0.126236036129307, 0.19478059424339, 
    -0.0942400584941163, 0.00164606439022587, 0.103017188497676, 
    -0.171784297555901, 0.151315967973733, -0.0127080774047862, 
    -0.140280647746261, 0.193663398872208, -0.12192595517384, 
    -0.0211465553337853, 0.180939061842622, -0.192624233760247, 
    0.0558451499354815, 0.12367774748912, -0.226205132909422, 
    0.192917279114909, 0.0541234054820051, -0.267248516538609, 
    0.226086491868972, -0.0342778285774787, -0.212526069659285, 
    0.261379801639104, -0.128474889245064, -0.148154984572706, 
    0.27435641639559, -0.167141757796018, -0.0487757658167641, 
    0.219658808791403, -0.240534279623928,
  0.0596650532494762, -0.0643393028443193, 0.113728593729297, 
    -0.132420972346581, 0.10691482869609, -0.0824345514437717, 
    0.00692313686376483, 0.0482755307784416, -0.0892308642385465, 
    0.163842202061563, -0.148716894990294, 0.092565027182356, 
    0.00705149048924581, -0.112766629851195, 0.176540291399719, 
    -0.190441689683812, 0.0872105622712378, 0.0429681915371264, 
    -0.149343239231789, 0.209383405612599, -0.191538084368487, 
    -0.0196817214993833, 0.165353369114805, -0.223017314845927, 
    0.158765005180121, 0.0545127298140329, -0.19935957115668, 
    0.195465120551461, -0.049021768542892, -0.125749455011779, 
    0.219929621859095, -0.155524067738249, -0.0443791048519432, 
    0.224567984051596, -0.170503265207885, -0.0221284824635361, 
    0.17723212606049, -0.168288319579871, -0.0260045746533278, 
    0.150350661368615, -0.149025185953801, 0.0180149756071444, 
    0.156440195988505, -0.190528788473358, 0.00200562451317899, 
    0.193503571479063, -0.189197803435024, 0.0247439319457884, 
    0.177432091265573, -0.235079905246189,
  0.0501674914843055, -0.0537946966560756, 0.0938223571588715, 
    -0.105928783457509, 0.0777889637594721, -0.0527957784760385, 
    -0.0130529206778161, 0.0590916402913252, -0.0869455855662132, 
    0.141187578448143, -0.104560371375234, 0.0381089576822819, 
    0.0636486742157325, -0.121432882364167, 0.142531892476561, 
    -0.11469158520825, -0.0167656285423597, 0.0991842081486424, 
    -0.14367846266838, 0.124811331507285, -0.0302177138509634, 
    -0.106785627207831, 0.167098453779061, -0.115558426772388, 
    -0.0207002816483014, 0.188440987485594, -0.1507134320214, 
    -0.0225075502271313, 0.163288948288649, -0.161233903736867, 
    0.0343726303327674, 0.152367077871853, -0.175944116672189, 
    0.0197219410610163, 0.15143444740628, -0.188059582340361, 
    0.0752907247036823, 0.175033348843358, -0.223132011367374, 
    0.0368345430976766, 0.172902314384449, -0.242870035027306, 
    -0.0204564059644503, 0.248143877482356, -0.164767986720996, 
    -0.147834451304637, 0.278030569148254, -0.123323195554827, 
    -0.209488365591347, 0.346992716014716,
  0.0665668789164214, -0.0709735259778762, 0.122085280956178, 
    -0.133426490172103, 0.0877089733669755, -0.0495286402645584, 
    -0.0388050142274977, 0.0971337025452712, -0.12379935262623, 
    0.180180903284194, -0.10321449856021, -0.00214802457013021, 
    0.14364655711664, -0.165955118060643, 0.14452069639356, 
    -0.0640225712965161, -0.121844679209888, 0.161879457510788, 
    -0.140900562646103, 0.0379425098789914, 0.124638114356879, 
    -0.155383244709925, 0.111891158188768, 0.0250247096124817, 
    -0.162710185038613, 0.184542759040475, 0.0018682396052637, 
    -0.194450306947551, 0.189805750686421, -0.00932794849026976, 
    -0.183690185231876, 0.224660648161821, -0.0112403428918101, 
    -0.237299866339362, 0.178155838586123, 0.0704423712751926, 
    -0.227366821906673, 0.0943075633428838, 0.180575509142265, 
    -0.187291756625742, 0.00352204223272315, 0.212785138434675, 
    -0.129555452739324, -0.0925498109982085, 0.196829449777967, 
    -0.00123141901695482, -0.186533873888436, 0.148861905245449, 
    0.118843187603513, -0.263458415411035,
  -0.0863559102718785, 0.091449468891956, -0.154704651854307, 
    0.162371947509744, -0.091191607210618, 0.0353865264436878, 
    0.0773511876391478, -0.145665116358487, 0.163024784606072, 
    -0.208057738364443, 0.0737394279674236, 0.0738923199065707, 
    -0.240508059139542, 0.180475346078395, -0.0840236732785922, 
    -0.0558405184572036, 0.234422338588341, -0.166335615287449, 
    0.0360589095984917, 0.138954815666733, -0.271040137066798, 
    0.0644171509666174, 0.115910461341568, -0.216270105399934, 
    0.145695188375206, 0.120403425954758, -0.212761058082712, 
    0.0681447522389741, 0.137128270301006, -0.188673838886407, 
    0.0542628040738814, 0.174728478153541, -0.171737776499792, 
    -0.0572643454134225, 0.195908149627053, -0.103954092709403, 
    -0.0823900577538445, 0.190708377599382, -0.00260466880733227, 
    -0.143239439263583, 0.117004510319955, 0.0630152370783706, 
    -0.161382643332062, 0.047765814536429, 0.155966372564493, 
    -0.0959958956241043, -0.101121393244139, 0.151326188285034, 
    0.0541073259386066, -0.19992897478182,
  -0.0423157728070973, 0.0445443096143945, -0.0742386196801624, 
    0.0750580986441309, -0.0355004891326733, 0.00604462690314818, 
    0.0471094914118779, -0.0763411595114512, 0.077211817370685, 
    -0.0864407334393765, 0.0105167446754644, 0.0600720925376651, 
    -0.125103924107295, 0.0611373537968674, 0.00708571620202378, 
    -0.0748875498139951, 0.110404544174423, -0.0365832376210904, 
    -0.0469421107357709, 0.111791424205285, -0.106159806796366, 
    -0.0481343092175485, 0.131212564987238, -0.0989595713135738, 
    -0.0315644045901469, 0.169637541296594, -0.0653251651638555, 
    -0.125040216779313, 0.15473192227769, -0.00580321416279598, 
    -0.153106872642433, 0.143430880180041, 0.0635849658886212, 
    -0.200016670175239, 0.0265423346838413, 0.188109013687845, 
    -0.165098904175761, -0.165669531836327, 0.228195113571073, 
    0.039073768867341, -0.242870009104105, 0.135044520042364, 
    0.246244803601337, -0.254304074738542, -0.202424746017054, 
    0.288570561732764, 0.0950926514103354, -0.30972783641073, 
    -0.039851767232696, 0.353923423046108,
  0.0656508767421972, -0.0685280975938962, 0.111790939167788, 
    -0.106894466133406, 0.0363540785276098, 0.0126109216594293, 
    -0.0878158752120855, 0.122001725485981, -0.107099019374963, 
    0.0939992396485289, 0.0335128018609458, -0.125743769452959, 
    0.176158995943143, -0.02323535513649, -0.0999950047755372, 
    0.170093921489178, -0.091638236670936, -0.0550435839614333, 
    0.156359499223341, -0.151267495027559, 0.00024628197730195, 
    0.166120333797457, -0.174334101190437, -0.00200146498770781, 
    0.201524370430192, -0.181148609087057, -0.111157652138625, 
    0.259276164376762, -0.0550138726471714, -0.209372756711823, 
    0.220380939791712, 0.0977938696255591, -0.248170632342384, 
    0.00927622385689427, 0.234204302859629, -0.131477255059896, 
    -0.12843009881845, 0.210341923327341, 0.118755107445885, 
    -0.184096315152213, -0.0165132890597565, 0.221872864706064, 
    0.0101090075698641, -0.211724939561405, -0.0030849394572999, 
    0.216541588717836, -0.0233615396205537, -0.190691094470503, 
    0.0214854220746271, 0.198124118433368,
  -0.0842895491674107, 0.0873375748522593, -0.13978055271205, 
    0.126875560438863, -0.0272560186584499, -0.0377736318952527, 
    0.123420716125562, -0.153260697153835, 0.11731819003659, 
    -0.0727003864487867, -0.0872934750508564, 0.173986553655245, 
    -0.175614527081651, -0.0457774992826611, 0.188910929385088, 
    -0.215251727562063, -0.0096955272279368, 0.160624805736655, 
    -0.196611931434917, 0.0677013552174558, 0.177234391524853, 
    -0.154218706773828, 0.0216717411884863, 0.151946924047924, 
    -0.171337709377311, -0.0769966141933401, 0.176311727445873, 
    -0.00642316226112243, -0.159306728430432, 0.0920032649353727, 
    0.10267046124048, -0.1696811280576, -0.0539082916334238, 
    0.204019623610852, 0.0296075045535156, -0.221627079970478, 
    0.0744565967271396, 0.284559138768238, -0.0485837119802985, 
    -0.212803778184407, 0.127020343133741, 0.19611545865321, 
    -0.118029316943386, -0.168240027075777, 0.102565017196415, 
    0.201627616493639, -0.0842179801387409, -0.173780716591456, 
    0.0540730581362501, 0.180161910653079,
  0.0764715232673198, -0.0787203976024438, 0.12383474137463, 
    -0.107008719673233, 0.0101752862361658, 0.0496063813676802, 
    -0.11693916033467, 0.132123349730255, -0.0874874531991639, 
    0.0278379950539355, 0.105048354398518, -0.152759702277399, 
    0.105877811240669, 0.0888723811375759, -0.187112585494795, 
    0.156989744671843, 0.103079474345294, -0.172993005773753, 
    0.118200650898288, 0.0569174549814159, -0.22639890653824, 
    0.0158808940320104, 0.148087080597612, -0.147840102280218, 
    -0.0408601865719445, 0.228252463266384, 0.00398372676541525, 
    -0.239563028022497, 0.0833992898648708, 0.191149324241396, 
    -0.189969347327307, -0.152051076974607, 0.199559947477634, 
    0.133696379639802, -0.186545616000334, -0.0965412027299309, 
    0.196339864670244, 0.138658439363508, -0.170628338337174, 
    -0.117330483819065, 0.191740350904974, 0.0879081127604204, 
    -0.194312148572457, -0.0863941175073156, 0.183779074345015, 
    0.173023915894084, -0.134771623607943, -0.161975076478326, 
    0.0835106882444596, 0.178047763550943,
  -0.043392629136436, 0.0442744505076482, -0.0680055346491968, 
    0.0546942270447863, 0.00454439287738146, -0.038339834727681, 
    0.0675007794967767, -0.0668407980652008, 0.0338344149189536, 
    0.0114466964373749, -0.0708634202731582, 0.0723302107094263, 
    -0.0152649768830257, -0.07060104978151, 0.0922934460379178, 
    -0.0423549591669289, -0.10206207798145, 0.0810199434719357, 
    -0.00052710572799448, -0.094074484067978, 0.100543352678999, 
    0.0826083461589731, -0.137256423556385, 0.0125913380869376, 
    0.147644101767229, -0.0849177794308585, -0.135609734194209, 
    0.115895181874557, 0.10055716489902, -0.138591429756222, 
    -0.0478623309235273, 0.180564763575041, 0.0533630154863428, 
    -0.198184319028969, -0.0922895560325716, 0.208193473949671, 
    0.0467523691392512, -0.2617160656156, -0.184356884986277, 
    0.152679765841041, 0.160917647659912, -0.18540148915822, 
    -0.285636484188163, 0.108865380424002, 0.371751083886236, 
    0.146573402989762, -0.287179735586463, -0.200922202881278, 
    0.186003118003069, 0.267140363234958,
  0.0866150037525887, -0.0876922911258312, 0.131849450717589, 
    -0.0990246751869817, -0.0255144576615223, 0.0915307381986504, 
    -0.132419842045411, 0.115229025674307, -0.0392602780642503, 
    -0.0642901669856466, 0.145620156250357, -0.105205271458564, 
    -0.0432606059588176, 0.143330752029067, -0.123078115436329, 
    -0.00318300477196261, 0.206291389083908, -0.083964891229479, 
    -0.0955660926361592, 0.198640461185766, -0.0605380201119772, 
    -0.213148443595887, 0.193139772353186, 0.109648127876695, 
    -0.289925289877457, -0.0613245889253682, 0.254534524247889, 
    0.0495118710686476, -0.23821371533169, -0.00897397106957762, 
    0.24641632619279, -0.0103790352296418, -0.235628155675563, 
    -0.03194162123134, 0.212959320900066, 0.0599315107923186, 
    -0.189027676364589, -0.166777321273982, 0.082536652509598, 
    0.159473113303374, -0.0694250715265487, -0.192000992837001, 
    -0.0598094722175711, 0.155902525029167, 0.182483733161875, 
    0.00408951059352906, -0.17105231718882, -0.0739423730872763, 
    0.122922057251224, 0.137580214251536,
  -0.0980331661964184, 0.0983494076072126, -0.144112531750373, 
    0.0990389626973315, 0.0487801951456008, -0.12013811818867, 
    0.141922872913141, -0.102432965044439, 0.00777588330897229, 
    0.117610301158975, -0.152011479881571, 0.056183949005186, 
    0.128367353130002, -0.12609760757221, 0.0317931560070419, 
    0.0965748800014467, -0.143698983237729, -0.0222898204363024, 
    0.150913102385178, -0.118224288171581, -0.105507252801756, 
    0.124028057186974, 0.0010350054030174, -0.139534124322344, 
    0.0685330681037733, 0.182197303871019, -0.00500785647415402, 
    -0.190616954676346, -0.0104194474675119, 0.180828877426877, 
    -0.0105586506897503, -0.22138124921417, -0.0715078778118373, 
    0.217305153943067, 0.187644630670211, -0.165293806111374, 
    -0.189214346487054, 0.0884434232453408, 0.286125924159586, 
    0.0986769295074655, -0.248926364556651, -0.190395877977439, 
    0.106008210055284, 0.24505998386624, 0.125532107129045, 
    -0.108521531575967, -0.214362911303233, -0.0331779278007287, 
    0.191289132991003, 0.170210154212734,
  0.136943535924702, -0.13655096926408, 0.196610349280779, 
    -0.126614475345347, -0.0850485997188493, 0.180544344029652, 
    -0.187437846315987, 0.114985206140953, 0.0212705858548998, 
    -0.196454800922335, 0.187632910301158, -0.0168675529088815, 
    -0.231308122399539, 0.117602713555714, 0.0590907789871578, 
    -0.186116104564284, 0.0628243845181467, 0.116685675198947, 
    -0.164946302627331, 0.0108724768344944, 0.213537305397142, 
    0.0200201231831168, -0.163690561235355, 0.0561194183855148, 
    0.163991228571875, -0.0785269609595838, -0.182419780067581, 
    0.0410640975255744, 0.175463782068439, -0.0238865290740825, 
    -0.179313437581143, -0.0102395692151211, 0.165047743259581, 
    0.0945063523320401, -0.0939262359716884, -0.139183016914588, 
    0.0472729190026494, 0.22283659390056, 0.196124645106704, 
    -0.032151351388568, -0.19657926492344, -0.0485728818136678, 
    0.173757330993586, 0.178410741016548, 0.0134259268534171, 
    -0.165359361039152, -0.182045121014813, 0.0137793886315559, 
    0.204689647934095, 0.160388448194015,
  -0.0830615798205929, 0.082312712268877, -0.11638646383319, 
    0.0697655816700454, 0.0612301250665563, -0.116115278727528, 
    0.105614806843569, -0.0518430003123939, -0.031312152727554, 
    0.134069701727986, -0.093588878909646, -0.0268767105963303, 
    0.160032772320162, -0.0276136950630579, -0.0938655025925727, 
    0.124056546377725, 0.058492182176148, -0.100913954125854, 
    0.035864960005311, 0.0882044355469941, -0.105582616782595, 
    -0.122735677910846, 0.13288296838455, 0.0838299093884266, 
    -0.179372204934899, -0.134168796557129, 0.0921446476768818, 
    0.170983022810814, -0.0360176694405627, -0.168727194119147, 
    0.0228209358731373, 0.213416412906891, 0.10646158822948, 
    -0.16809850190534, -0.234940691765837, 0.0402072435706848, 
    0.221768226806033, 0.163842336842928, -0.0297116825049603, 
    -0.148439985419858, -0.0384733857107194, 0.149721691370456, 
    0.232637938315596, 0.070007693936674, -0.163224475648307, 
    -0.308364898675595, -0.206778691550853, 0.097152269618977, 
    0.336227066324776, 0.235123716954211,
  0.0536865971940169, -0.0528985692799132, 0.0735281106198691, 
    -0.0409949877289268, -0.0449206529586529, 0.0783403598680427, 
    -0.0627354861461601, 0.0226297889119163, 0.0303173068620094, 
    -0.0927582168907775, 0.0461664448076101, 0.0381323057884125, 
    -0.107987076953455, -0.0103400877058627, 0.089263944610748, 
    -0.075393287286523, -0.0945700884880315, 0.0681130274275263, 
    0.028671175967939, -0.101653756619999, 0.0196028231338517, 
    0.118223651600625, -0.0618006112455012, -0.111809190096833, 
    0.098288004630118, 0.174432209157552, 0.0203804260718334, 
    -0.172975641117523, -0.084727822047885, 0.140690498920118, 
    0.111591100252463, -0.120605141112291, -0.19112771309306, 
    -0.0104979578365148, 0.172707832206771, 0.12918278739234, 
    -0.0915368366696026, -0.272309086040295, -0.285858676360851, 
    -0.0583583076906418, 0.238523494748542, 0.231210346465556, 
    0.0466562474875999, -0.168973967262031, -0.293245666789357, 
    -0.294947065408369, -0.108212703105101, 0.158964766538406, 
    0.331551208570933, 0.210961787293921,
  -0.0793257646266844, 0.0774565781375864, -0.104727844341598, 
    0.0513192047184727, 0.0776655598646381, -0.121653116289491, 
    0.0781595605232532, -0.00808529960776405, -0.0652616358443905, 
    0.143424354968855, -0.0305912750476055, -0.0980389418765719, 
    0.150245346996571, 0.0791269520338531, -0.174591309090142, 
    0.0727312705050064, 0.246028805965538, -0.0670358261049257, 
    -0.170796821520491, 0.193961423285015, 0.142630231161255, 
    -0.146448255755136, -0.0573710531526706, 0.176955322873462, 
    0.0441073764457486, -0.225025417592772, -0.217020119887232, 
    0.103741318197598, 0.254994075952371, 0.00803283253765238, 
    -0.258608051897269, -0.173526257221297, 0.0931816554716651, 
    0.278750798663553, 0.213271621708234, -0.102971895546543, 
    -0.252888828038019, -0.199602317774639, -0.0565082583311839, 
    0.0892196594077993, 0.117397239075645, -0.000353526121857814, 
    -0.136407615913793, -0.169022966670588, -0.131485392008132, 
    -0.0668457785029179, 0.0228063106515857, 0.0886948725821047, 
    0.116746902369161, 0.0650824407806302,
  0.0412569859224389, -0.0399783842495507, 0.0527766908618346, 
    -0.0227869785944975, -0.0447827080683517, 0.0650497238053017, 
    -0.0336595483203724, -0.00664733825613916, 0.041281983793104, 
    -0.0737443191376246, -0.00151534004054371, 0.0649337794281415, 
    -0.0654491990065098, -0.0645852623947947, 0.0961256321391017, 
    -0.0120276170436447, -0.152780959148699, 0.0066070932182404, 
    0.132624089250204, -0.0872484901115982, -0.148165529868407, 
    0.00964915795272815, 0.103996342994421, -0.0246185220184443, 
    -0.118524641805569, -0.0294604820662762, 0.0808863579776703, 
    0.0905732222736251, -0.0149951172083752, -0.0939031967526352, 
    -0.0263234310188807, 0.0938512566728799, 0.120373558027056, 
    0.0279276127646266, -0.0803637349325971, -0.11094479720993, 
    -0.0141359655945082, 0.125062155646191, 0.243433834330392, 
    0.207636098998671, -0.0536387679197573, -0.295308858246371, 
    -0.468272106429378, -0.384041615661889, -0.197866331225949, 
    -0.00565251719983096, 0.178661413330955, 0.2520407460514, 
    0.256825939566225, 0.1297365471744,
  -0.0699305873031767, 0.0675172211356762, -0.0881032677355775, 
    0.0355523240596959, 0.0791590847341674, -0.111290024438393, 
    0.0511531393980977, 0.0197920560203374, -0.0749816838859021, 
    0.122486499730298, 0.0166369879230446, -0.118644990724228, 
    0.0968297121449214, 0.124492967105066, -0.159960397265555, 
    -0.00254129193860447, 0.264744981484397, 0.0145648741042707, 
    -0.247042326384858, 0.12206479846445, 0.295897564451863, 
    0.0540897872791466, -0.222042198999618, -0.0407659358300881, 
    0.252594127792601, 0.207566363826209, -0.0268247862152109, 
    -0.238096071930249, -0.145856851701036, 0.13929447039985, 
    0.21927865953371, 0.0170840900484376, -0.189381311966076, 
    -0.239628729737765, -0.131447456955923, 0.103921474881276, 
    0.202044194477031, 0.183885817266163, 0.136563253379176, 
    0.0395984039965077, -0.0930540943667824, -0.148798527479073, 
    -0.172407501866901, -0.117729202080337, -0.0396156127964867, 
    0.03709647830802, 0.104470044466122, 0.118752681588558, 
    0.109616885376234, 0.0530158968979732,
  0.00430248001786901, -0.00412766591247335, 0.00527631764955713, 
    -0.00186475343768001, -0.00519309810948118, 0.00692199992078775, 
    -0.00249505085449126, -0.00210454488968757, 0.0050635476650744, 
    -0.00710780313029961, -0.00249757324534046, 0.00795368350885489, 
    -0.0041549768032856, -0.008819582714427, 0.00888740485823656, 
    0.00259121047691597, -0.0155246457611291, -0.00354809518290925, 
    0.0160397744150947, -0.00386208644302321, -0.0207380993206783, 
    -0.0109001497662382, 0.0161456938920876, 0.0119895647874689, 
    -0.0170338753464224, -0.0286587738861417, -0.0156216922382283, 
    0.0155750461081113, 0.0271543088283659, 0.00398543624908954, 
    -0.0254152909345831, -0.0296192315961797, -0.0114292659528309, 
    0.0178917411462621, 0.0363757856366919, 0.0258821355192849, 
    -0.00770508461650904, -0.0475049935124036, -0.090218511588614, 
    -0.0929313590020056, -0.0101865421599864, 0.0947765089524154, 
    0.204418304201369, 0.245202458327659, 0.288912402552184, 
    0.403143287462294, 0.511010131629722, 0.448628649478795, 
    0.356938816533663, 0.160733646581306,
  -0.0318193038990164, 0.0302439396558212, -0.0374827341465706, 
    0.0104292110093827, 0.0414614321230054, -0.0514413515088494, 
    0.011204043509026, 0.0245489383388328, -0.0408422288336503, 
    0.0455678713120931, 0.0331492973576601, -0.0613161399796039, 
    0.00801516124942491, 0.0692241103697346, -0.0465306574508197, 
    -0.0411788417650447, 0.0855399107023603, 0.0463740008704997, 
    -0.10063790107532, -0.0132486717931469, 0.136291831915782, 
    0.132699402706055, -0.100341441573979, -0.158284985317798, 
    0.0760258012728881, 0.284353177793358, 0.284037295241465, 
    0.0100076745230136, -0.251878902685959, -0.219230050883728, 
    0.094090193198908, 0.375517985799744, 0.424369572802296, 
    0.213510516017365, -0.0627636797038212, -0.30875747395035, 
    -0.284935672071074, -0.147751529439816, -0.0354990494473404, 
    0.0551441100166982, 0.0993705724401437, 0.077938598855962, 
    0.0604152256916053, 0.0379137005659627, 0.0217292022548121, 
    0.0153508654640211, 0.012588811771621, 0.00860918037176103, 
    0.00573288660972843, 0.00234691020028275,
  0.067941821694873, -0.0635411261783642, 0.0744395897995344, 
    -0.010512402464212, -0.097437749030436, 0.107820934809132, 
    0.00329230491519459, -0.0814005327361751, 0.0913880738719121, 
    -0.0602110813687434, -0.112995662679423, 0.114495339455184, 
    0.0708930016218497, -0.111023880193032, -0.0012564333453039, 
    0.116966317752518, 0.0016902162563434, -0.0832493339588269, 
    0.0300089215523634, 0.0898390750588349, -0.0287172424620359, 
    -0.130373470306682, 0.00129991797029275, 0.146438307026949, 
    0.0658886689945737, -0.122324166826218, -0.244765119752145, 
    -0.205152305456542, -0.0264198431917315, 0.166027477476428, 
    0.192764373415581, 0.0785215140512208, -0.0526527082035273, 
    -0.181328190173404, -0.295283582624501, -0.319685293575326, 
    -0.180679698607431, 0.00368233023875865, 0.20282127479378, 
    0.381970244793494, 0.370295535374597, 0.206398789365058, 
    0.113342839022872, 0.0544702892863231, 0.0231881112495557, 
    0.0111509966885522, 0.00627052456402963, 0.00323225084187689, 
    0.00169353939690891, 0.000599603830641989,
  -0.120146523747658, 0.112064156180145, -0.130027830240464, 
    0.0153080976670145, 0.174413872899787, -0.189519693243292, 
    -0.0136848469225982, 0.151362230066836, -0.161140500028376, 
    0.0938635767938369, 0.208830288018195, -0.192825904172362, 
    -0.149067361639956, 0.175804426992281, 0.0328922157607373, 
    -0.201362296429276, -0.0605349795036754, 0.121724623819124, 
    0.0109431993156707, -0.144663484899121, -0.0384179437101665, 
    0.115210752218509, 0.0477323452859597, -0.114046471528863, 
    -0.111084442927297, 0.0190495339320411, 0.130731994511235, 
    0.163849513173466, 0.0876552039147947, -0.0574052890419506, 
    -0.149433241797915, -0.155221351755521, -0.122862164052223, 
    -0.0561361815791772, 0.00738690466744474, 0.0710946676948524, 
    0.0947641218029091, 0.131115724883143, 0.259848924790497, 
    0.406154905322588, 0.370522892062297, 0.198497316105245, 
    0.104515795862478, 0.0485730946324161, 0.0199766658505842, 
    0.00920669855105746, 0.00494986323177033, 0.0024594970123562, 
    0.00124600268240569, 0.000431599848925747,
  0.118599392175193, -0.110294215677838, 0.126605376520028, 
    -0.0115779387513873, -0.174314781142208, 0.185662890571531, 
    0.022027709790399, -0.157146252277771, 0.158045633515481, 
    -0.0784645782307321, -0.21478107006625, 0.178474614364367, 
    0.171744786545712, -0.148558510717426, -0.0651284312461781, 
    0.188205901207724, 0.12044560281299, -0.0866240394828362, 
    -0.0793490034455677, 0.116545752348158, 0.130180670059267, 
    0.0258064010078862, -0.0879645600660756, -0.0596117502847668, 
    0.0687518599277595, 0.170071321427298, 0.210051687399771, 
    0.128403996687658, -0.0244234044570947, -0.150090237504459, 
    -0.137718730800551, -0.0322152182512663, 0.0739808909538359, 
    0.176727755520459, 0.284699459770275, 0.337096798935605, 
    0.246188691353676, 0.155877483357006, 0.177336845151228, 
    0.236333974065094, 0.202802266060147, 0.104293389550023, 
    0.052569646951635, 0.0235890354390037, 0.00936070579885667, 
    0.00413030554259081, 0.00212018678424362, 0.00101383347688187, 
    0.000495615305043041, 0.000167671459733018,
  -0.0505570276269597, 0.0467807238410043, -0.0527117850878148, 
    0.00242538167047382, 0.0757093084297678, -0.0779599838650464, 
    -0.0154827063797058, 0.0722155471090221, -0.0661334523670798, 
    0.0228052630871986, 0.0965544235719161, -0.0662405546277881, 
    -0.089465974148638, 0.0429711440796208, 0.050039763771263, 
    -0.0681000291120509, -0.0916230046118664, 0.00784176387297796, 
    0.079952076616051, -0.0207191034340381, -0.112936768685196, 
    -0.118847394189662, 0.050357287526337, 0.153629676739369, 
    0.0346083117796243, -0.162613743254226, -0.305528149709907, 
    -0.301340239099808, -0.139047582633395, 0.113803800842278, 
    0.274533594376395, 0.315739797388368, 0.322238221606936, 
    0.298051387474071, 0.319601697111097, 0.306141759565749, 
    0.195732089288278, 0.0955122503910602, 0.0721367323030371, 
    0.0783267164353209, 0.0612662082711073, 0.0295640061855885, 
    0.0139170792839115, 0.00590684439164454, 0.00221608820712615, 
    0.000914229377029885, 0.000436733688831888, 0.000196568267185904, 
    9.07420675675182e-05, 2.95327942402218e-05,
  0.0540446597686605, -0.0489089766833216, 0.0505461530597313, 
    0.00847692395497177, -0.0852427221601747, 0.0755636347391343, 
    0.0434302822111853, -0.0957029944817333, 0.0579459493648195, 
    0.0285041123275096, -0.105992229055929, 0.0110601861741901, 
    0.13848507140889, 0.0662239788592648, -0.11761815196129, 
    -0.0351783229263744, 0.179245502693218, 0.141558997944916, 
    -0.176303847921513, -0.177261043094574, 0.138921416682697, 
    0.412459929011249, 0.0989060612359498, -0.397083064607573, 
    -0.465375316932979, -0.280180378199145, -0.148697381355074, 
    0.0075895804657375, 0.150138338544004, 0.227270297304986, 
    0.185833141774505, 0.106185362676542, 0.060638307434773, 
    0.0302656296950024, 0.018105176624709, 0.0110964287084711, 
    0.00544532752374563, 0.0019067097257232, 0.00078932840650271, 
    0.00051507181892983, 0.00029680631840898, 0.000114545225458524, 
    4.23216915870123e-05, 1.46542155826801e-05, 4.49434382439476e-06, 
    1.46925773676941e-06, 5.46503058452158e-07, 1.97868413288487e-07, 
    7.37577441580223e-08, 2.05963924671092e-08,
  -0.0203667021652573, 0.0181981961822461, -0.0178329104144336, 
    -0.00537751543216146, 0.032475590789639, -0.0263199683779357, 
    -0.02147625584237, 0.03837781832495, -0.017613178515279, 
    -0.0218697359711802, 0.035061216979321, 0.0099582142864169, 
    -0.0504565032657856, -0.0460123308674765, 0.0434590677340653, 
    0.0397424190753911, -0.0488044787089373, -0.0657116980266826, 
    0.0442629900869271, 0.0850354054604809, 0.00111863976107243, 
    -0.0915143444475988, -0.0563695821555198, 0.0575046321496422, 
    0.1247711412071, 0.169716010189061, 0.267260003957383, 0.390737432549997, 
    0.508784609165724, 0.517396048487458, 0.349168423535754, 
    0.169287832266615, 0.0832434129231713, 0.0355238882268261, 
    0.017848901458181, 0.00927117576698763, 0.00407818255928771, 
    0.0012788868331605, 0.000449073580285104, 0.000245550509671593, 
    0.00012416055561697, 4.33032986971833e-05, 1.43339723490626e-05, 
    4.51147263069673e-06, 1.2601237921022e-06, 3.71148158594189e-07, 
    1.2342985315596e-07, 4.04363126536736e-08, 1.36220711313555e-08, 
    3.52230720011e-09,
  0.117202803988099, -0.103359717842943, 0.0955758334492814, 
    0.0430265930737008, -0.186729624876855, 0.137172930472455, 
    0.150173635756132, -0.227620758111195, 0.0721908034156859, 
    0.186176976574369, -0.152583076692039, -0.134661545595115, 
    0.232926227118425, 0.340905164494851, -0.185350178679555, 
    -0.339147305782618, 0.0559997548996402, 0.292278441698701, 
    -0.0219982744684635, -0.348295907497537, -0.275247867766231, 
    -0.146066591574644, 0.089794752916485, 0.248276212227361, 
    0.198454839519071, 0.0999349054245886, 0.0640552192096275, 
    0.0455112161683057, 0.0378861468397782, 0.0300275553190989, 
    0.0174359196457925, 0.00740306869291246, 0.00321921505760703, 
    0.00121245905741276, 0.000530077474994157, 0.000239697078306914, 
    9.56372845761114e-05, 2.7265684890754e-05, 8.40952375907403e-06, 
    3.98141440929978e-06, 1.79530394833201e-06, 5.71562768855619e-07, 
    1.71399961467094e-07, 4.94418479878834e-08, 1.26816214698749e-08, 
    3.40141746725179e-09, 1.02346037743755e-09, 3.06297323567797e-10, 
    9.40631203224704e-11, 2.26196880841024e-11,
  -0.114916960704746, 0.0983535849433709, -0.0785022013257877, 
    -0.0662344394929959, 0.175527524741096, -0.0989751689803541, 
    -0.191364501055474, 0.215685288904789, 0.000714190327719276, 
    -0.284185282788531, -0.0107598964402073, 0.245447230693458, 
    0.027181091425466, -0.244820601492675, -0.0626377116194067, 
    0.248765439707876, 0.375955287663377, 0.249048169853944, 
    -0.255571085006604, -0.438886526701878, -0.200540208233905, 
    0.016827150243017, 0.16088457157139, 0.18443488884248, 0.10745337451859, 
    0.0396817986895088, 0.0175115196283818, 0.00790589317563058, 
    0.00417701488507158, 0.0023132394183426, 0.00104167233519912, 
    0.000351306016979871, 0.000122869437060811, 3.72763341159233e-05, 
    1.28497630853997e-05, 4.55032414740893e-06, 1.5097601387883e-06, 
    3.60486955628098e-07, 8.91210098383686e-08, 3.2920254178072e-08, 
    1.20174675398149e-08, 3.2155681742984e-09, 7.99703497053183e-10, 
    1.94918506149937e-10, 4.24107022277848e-11, 9.52391093988376e-12, 
    2.37288285804688e-12, 5.97457389189053e-13, 1.5349081890538e-13, 
    3.19157985791226e-14,
  0.132043346281473, -0.109375111930082, 0.0721130814531381, 
    0.101233371001693, -0.18157245506664, 0.0669216477689041, 
    0.24576978019606, -0.206888991454821, -0.0828997378121664, 
    0.378701255634617, 0.235398983884816, -0.277735744703887, 
    -0.405993884648436, -0.255408139574127, 0.201250670296041, 
    0.338662190106702, 0.16873318616253, -0.00479768956662743, 
    -0.154185750122563, -0.127823994095278, -0.000525683208326517, 
    0.139050215878871, 0.184673557461708, 0.140321972785055, 
    0.0650811951808068, 0.0194918133477319, 0.00684490172652098, 
    0.00239535122973072, 0.000962417410850588, 0.000413514783728603, 
    0.000152039810671107, 4.25089845077709e-05, 1.24087591544446e-05, 
    3.1535212277308e-06, 8.97957148403653e-07, 2.60476831512589e-07, 
    7.35841401473471e-08, 1.50615031567251e-08, 3.11368911842619e-09, 
    9.4233441151134e-10, 2.87493660510934e-10, 6.60326234450508e-11, 
    1.39516341090188e-11, 2.92774026143696e-12, 5.50287049736069e-13, 
    1.05781427507393e-13, 2.23737241869499e-14, 4.83897664954409e-15, 
    1.06166032410874e-15, 1.930997546617e-16,
  -0.0258947587097487, 0.0212117457683873, -0.012978344663839, 
    -0.021314332966886, 0.0338702793989972, -0.0100446788427811, 
    -0.0485797105246547, 0.0368408739553722, 0.0207320977575759, 
    -0.074192819337242, -0.0591345654703707, 0.0477990501891349, 
    0.0992519986310838, 0.0947540377671689, -0.0294812559114359, 
    -0.111938870265267, -0.131053727904261, -0.116517295313223, 
    0.0412045362768269, 0.175745955598946, 0.252670900505743, 
    0.536035031541384, 0.583597827773957, 0.401278129379265, 
    0.17462004712348, 0.0493352269422484, 0.0162780601355663, 
    0.00532637453871802, 0.00199171455775664, 0.000798410715271668, 
    0.0002769952003857, 7.33592700797672e-05, 2.03145800768537e-05, 
    4.90368390465682e-06, 1.32157855142243e-06, 3.61935905338695e-07, 
    9.7466993546683e-08, 1.90548435154641e-08, 3.74064963584374e-09, 
    1.06918838573905e-09, 3.09454577088379e-10, 6.79061954989998e-11, 
    1.3668742825953e-11, 2.7422822339563e-12, 4.93240522644281e-13, 
    9.05187876931236e-14, 1.82369842331614e-14, 3.76906549087733e-15, 
    7.88779396150248e-16, 1.37718926411136e-16,
  0.0277480971624542, -0.0205781058381479, 0.0037589725546418, 
    0.0323868736933282, -0.0139412352651495, -0.0133172456961026, 
    0.0294717648382994, 0.00066558033323586, -0.0289119323304873, 
    0.0238900796632415, 0.070951415573366, 0.0382170271744044, 
    -0.0517498181939061, -0.163356901489536, -0.139605803390254, 
    0.0199729212301122, 0.283632175152675, 0.629922379135002, 
    0.593898732921678, 0.314246288667432, 0.0939146622834692, 
    0.0376076994974383, 0.0184814845198962, 0.00727909205275401, 
    0.00210545431797018, 0.000408355924512683, 9.07311845569652e-05, 
    1.96306978412422e-05, 4.75005020439507e-06, 1.23574070785748e-06, 
    2.9281181369877e-07, 5.40932941065154e-08, 1.05144362181604e-08, 
    1.7972126344215e-09, 3.36556153917716e-10, 6.30823857981116e-11, 
    1.22208268275747e-11, 1.73937951840714e-12, 2.41746873953792e-13, 
    4.74664822965363e-14, 9.62758281981323e-15, 1.54007437518799e-15, 
    2.22270715653265e-16, 3.26039182940127e-17, 4.31279187592175e-18, 
    5.74511070064087e-19, 8.29449002531982e-20, 1.25120983018031e-20, 
    1.88859527444729e-21, 2.46330949900485e-22,
  -0.367278476709736, 0.262532745197317, -0.00548353817145204, 
    -0.452922488316329, 0.0585226150397099, 0.248464983321362, 
    -0.17273946797706, -0.145223363917183, 0.214197890438535, 
    0.0359980493766655, -0.309444771551474, -0.347039193922453, 
    -0.0719928390708123, 0.199746673400753, 0.314266449803412, 
    0.201764885861522, 0.0974657918627203, 0.102699849630692, 
    0.0753833645062184, 0.0343483403064959, 0.00908038709610053, 
    0.00301971997567549, 0.00127234077568019, 0.00043942717916452, 
    0.000114167469266074, 2.00374989384569e-05, 4.01318814377557e-06, 
    7.80639416529427e-07, 1.69178204184583e-07, 3.93848084793148e-08, 
    8.42643959149612e-09, 1.41201702482381e-09, 2.4918747006984e-10, 
    3.87591071287695e-11, 6.57850353525063e-12, 1.11373918215668e-12, 
    1.96854563436138e-13, 2.56338986406086e-14, 3.24269673764635e-15, 
    5.75737774444614e-16, 1.05950950423499e-16, 1.55105958952302e-17, 
    2.04092824968178e-18, 2.7410861547965e-19, 3.32447488111116e-20, 
    4.04895403166302e-21, 5.32926114502059e-22, 7.35959009689259e-23, 
    1.0138830264667e-23, 1.21610654333156e-24,
  0.268617763340798, -0.187447020778693, -0.0160933670572683, 
    0.338900577454874, 0.0177299792468559, -0.205413275701481, 
    0.0120158887858944, 0.146813405315062, -0.0490343190110386, 
    -0.161519956112845, -0.135620172226399, -0.0153208181857994, 
    0.159029424679618, 0.462859563781018, 0.548968393333866, 
    0.311484015597406, 0.11859102253263, 0.0976636701402696, 
    0.0632217845884089, 0.026513952963142, 0.00654916646703186, 
    0.00197514902713568, 0.000764812946589671, 0.00024522900573404, 
    5.98712085921077e-05, 9.91464158196835e-06, 1.86972942159389e-06, 
    3.42007568547194e-07, 6.95636706010515e-08, 1.51899461651374e-08, 
    3.06236706320266e-09, 4.84750080040342e-10, 8.08462408023308e-11, 
    1.18993028212035e-11, 1.90700032875623e-12, 3.04281713992709e-13, 
    5.09587678310775e-14, 6.29696721605371e-15, 7.53876871554535e-16, 
    1.26231220479126e-16, 2.1944543473765e-17, 3.04903999209929e-18, 
    3.79993750096277e-19, 4.84492286545847e-20, 5.58261101504988e-21, 
    6.44971096411305e-22, 8.04022921662617e-23, 1.0540299583633e-23, 
    1.37607096285085e-24, 1.57051427618319e-25,
  -0.189576900783103, 0.126776985966171, 0.0351218392486172, 
    -0.243989712296532, -0.0865697788233302, 0.160294137625027, 
    0.139002586111467, -0.118180809059881, -0.118102091873484, 
    0.213124068149267, 0.531084457056465, 0.532710359800162, 
    0.271411339528869, 0.249773836841099, 0.216504192643318, 
    0.10535495963778, 0.0317550015773866, 0.0195900062420543, 
    0.0106088758008497, 0.00392121445629832, 0.000872941801283634, 
    0.000228062599034582, 7.77337489350396e-05, 2.22248064484922e-05, 
    4.92019675219421e-06, 7.43314386702065e-07, 1.27491548457103e-07, 
    2.11734086008992e-08, 3.89949075584985e-09, 7.70192833916107e-10, 
    1.41358403204103e-10, 2.04455942275616e-11, 3.11749630097194e-12, 
    4.2032236553222e-13, 6.15100936558622e-14, 8.93756677219491e-15, 
    1.37357898339222e-15, 1.56114819489332e-16, 1.71252919561122e-17, 
    2.61385814743934e-18, 4.15170628415988e-19, 5.3069871944885e-20, 
    6.06608587859122e-21, 7.1177413414217e-22, 7.55646184024924e-23, 
    8.02534582215533e-24, 9.17549084929629e-25, 1.10695855494825e-25, 
    1.326486478793e-26, 1.39787632742123e-27,
  0.171426863470507, -0.0934953979070935, -0.116149067371474, 
    0.187055596384452, 0.325308175171415, -0.0413714888675296, 
    -0.575953864424755, -0.23976898813676, 0.48083983641914, 
    0.376399205978723, 0.186574893101834, 0.0908614613330319, 
    0.0247134179509984, 0.00823803739893362, 0.00357211986638003, 
    0.0011293839807384, 0.000207805311898621, 6.73837708930013e-05, 
    2.20919250627318e-05, 5.47163797100293e-06, 8.68492141219382e-07, 
    1.47694457731957e-07, 3.37832432822937e-08, 6.65768188802214e-09, 
    1.05885779137227e-09, 1.16951169203754e-10, 1.45397990289922e-11, 
    1.7432996386995e-12, 2.30201315323958e-13, 3.24804903425942e-14, 
    4.32874717783822e-15, 4.59424487062559e-16, 5.14603988062198e-17, 
    5.12711167811271e-18, 5.49494389048027e-19, 5.80318136121988e-20, 
    6.61840304452076e-21, 5.61873108545103e-22, 4.5589598168428e-23, 
    5.0728274227268e-24, 5.906716286411e-25, 5.64416396396566e-26, 
    4.78013793508695e-27, 4.19584558136766e-28, 3.34361963715916e-29, 
    2.6485157862547e-30, 2.24363980603876e-31, 2.02542235814347e-32, 
    1.80182236845492e-33, 1.43297285215064e-34,
  -0.311549456929375, 0.101054982069062, 0.43633336828762, 
    0.0846833666858283, -0.481315883853674, -0.495299020981681, 
    -0.09237541243815, 0.234223176074691, 0.364505240789476, 
    0.143534938539624, 0.0350518439553528, 0.00945208472773854, 
    0.00158922903899911, 0.000281418774853916, 6.7112763544785e-05, 
    1.32569124113234e-05, 1.52513356421922e-06, 2.81100945566048e-07, 
    5.51414342629889e-08, 8.64459018857599e-09, 9.14798633279309e-10, 
    9.73760313660525e-11, 1.41766992882109e-11, 1.80628183682323e-12, 
    1.91477979803988e-13, 1.43229746537798e-14, 1.1967463688781e-15, 
    9.61810337492252e-17, 8.46897053762253e-18, 7.93733295229885e-19, 
    7.11402682473783e-20, 5.12598060137888e-21, 3.89949680191023e-22, 
    2.6536763695435e-23, 1.92710468005973e-24, 1.37020009060255e-25, 
    1.0703135917066e-26, 6.26033509022655e-28, 3.47326581438716e-29, 
    2.60940450562769e-30, 2.05920751593331e-31, 1.35678049240076e-32, 
    7.85999564792761e-34, 4.75935859670043e-35, 2.62459001568838e-36, 
    1.4305214180275e-37, 8.29014409341561e-39, 5.16576936011791e-40, 
    3.14792794067776e-41, 1.7389981732515e-42,
  -0.285506413822269, 0.0653820197463286, 0.470896463548721, 
    0.33114212500934, 0.13557035336042, -0.0288531942057562, 
    -0.297014351680953, -0.487979660161099, -0.461777074737449, 
    -0.151739304058101, -0.0307653611817138, -0.00698219530290038, 
    -0.00101301278248699, -0.00015058867996703, -3.02113868827481e-05, 
    -5.14376786493852e-06, -5.11679560104663e-07, -7.98959701585612e-08, 
    -1.33921208348462e-08, -1.81425604838908e-09, -1.68035992987112e-10, 
    -1.54334087696548e-11, -1.94519988008888e-12, -2.15247470077824e-13, 
    -1.99562998011495e-14, -1.31100914575756e-15, -9.60115953712798e-17, 
    -6.75956945003553e-18, -5.20757881115833e-19, -4.26579461690561e-20, 
    -3.35130106187532e-21, -2.12184304658919e-22, -1.41836117569189e-23, 
    -8.49429199299726e-25, -5.41737101174286e-26, -3.37740603934904e-27, 
    -2.32305283168407e-28, -1.19826977313141e-29, -5.85237471566221e-31, 
    -3.8581379129978e-32, -2.67381810319875e-33, -1.55399941009481e-34, 
    -7.92449799449533e-36, -4.2329670908641e-37, -2.06093302513441e-38, 
    -9.90304357685205e-40, -5.05199228700904e-41, -2.77762901953666e-42, 
    -1.49043466832557e-43, -7.27507863347263e-45,
  0.210905335612749, -0.0374047758781134, -0.372927636697893, 
    -0.357491962537865, -0.449264926385863, -0.416820301652928, 
    -0.336734665723288, -0.344186799259696, -0.270048233676705, 
    -0.081519683645468, -0.0151537551295286, -0.00316864999875375, 
    -0.000428134040552309, -5.86039627746293e-05, -1.08319813617107e-05, 
    -1.71620038856938e-06, -1.59130903955119e-07, -2.29598967990304e-08, 
    -3.5684481933861e-09, -4.5034329676227e-10, -3.90751865032839e-11, 
    -3.34153986301772e-12, -3.92678905922406e-13, -4.05675597050735e-14, 
    -3.52212753823434e-15, -2.17081327652498e-16, -1.49020566112701e-17, 
    -9.83209460350545e-19, -7.09472854689216e-20, -5.4408532712082e-21, 
    -4.00673735737965e-22, -2.38055496773525e-23, -1.49326202813507e-24, 
    -8.3976522694292e-26, -5.02457781064329e-27, -2.93678273099941e-28, 
    -1.89728279715992e-29, -9.19828329324268e-31, -4.21918309285531e-32, 
    -2.60854112636688e-33, -1.69599489892421e-34, -9.26550127720028e-36, 
    -4.43723364469199e-37, -2.22805634538118e-38, -1.02010992525941e-39, 
    -4.606494703217e-41, -2.20696771199352e-42, -1.14075471965199e-43, 
    -5.74928479282863e-45, -2.6398770869655e-46,
  0.546969126219743, 0.8124258148104, 0.200344663278698, 0.0254126059872762, 
    0.00227485059461268, 0.000331604134429685, 2.8735392944219e-05, 
    3.50592786489041e-06, 4.49750218399525e-07, 3.83150102022746e-08, 
    1.98644551031961e-09, 1.18794165228273e-10, 5.05059395525891e-12, 
    1.98663445839617e-13, 1.05351194859532e-14, 5.18344353642473e-16, 
    1.52625054183007e-17, 6.47740019078699e-19, 3.03728479673799e-20, 
    1.20136000807672e-21, 3.44865809836861e-23, 9.22866413124132e-25, 
    3.43200926031974e-26, 1.13422497357183e-27, 3.23702234606323e-29, 
    6.67785329567701e-31, 1.51714037242784e-32, 3.2905217040106e-34, 
    7.68824213208244e-36, 1.86180025151198e-37, 4.22177363236416e-39, 
    7.33128736011347e-41, 1.20684238301875e-42, 1.50539306122237e-44, 
    1.45977486065955e-46, 7.52489643149132e-49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0 ;

 obs_scale = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1 ;

 NLmodel_initial = 17.7537797833681, 17.6128448875051, 17.3864659361365, 
    17.1345272907666, 17.418381759779, 17.1207431184336, 16.8590772750634, 
    16.4974815056981, 16.4861379993712, 16.5543740624218, 16.4610111479159, 
    16.390141729834, 16.1503622931495, 15.6786201376981, 14.842076447458, 
    14.9081996219385, 14.6818498371035, 14.6575606456933, 14.4105201636211, 
    13.5999557170209, 13.2098864041791, 13.3550665798365, 13.1907037692145, 
    13.1080469623982, 13.2820554045892, 13.5184947825299, 13.7771438883842, 
    13.6220601640567, 12.8953146434843, 12.4432877790404, 12.6614103868119, 
    12.8887228673124, 12.323317469353, 11.3390329870824, 11.1062612764637, 
    11.0916940765239, 10.8865965068421, 10.957313183357, 11.0779284719594, 
    11.0903069221219, 10.8165942985575, 10.706517795932, 10.4962396796461, 
    10.4190119235619, 10.3398849474556, 10.0695518143835, 10.0743225734044, 
    9.86439754301222, 9.70421428013077, 9.61147890905523, 9.21116938375195, 
    17.7278526369271, 17.6894537918638, 17.4883591008051, 17.4137565234566, 
    17.2516728956583, 17.1622576366573, 16.8347739310962, 16.4287496640414, 
    16.3605071474149, 16.540823419583, 16.4184119585769, 16.3173946810696, 
    16.1115550015357, 15.5923842760269, 14.9414319588734, 14.9186724661149, 
    14.5979920623309, 14.7162613198676, 14.4842005738101, 13.7820047019333, 
    13.5292939305537, 13.6012222039863, 13.2381665797561, 12.989170861375, 
    13.3936698987732, 13.639192832316, 13.73418234602, 13.0277016589256, 
    12.4179070648414, 12.3957611970871, 12.4517252388761, 12.292080019991, 
    11.5703737825703, 11.2177851887946, 11.122120098356, 10.9478417142391, 
    10.8626701853369, 10.9795224928024, 11.1752661268791, 11.0641074074609, 
    10.7264946326577, 10.6999695875331, 10.4702741923128, 10.2470465103751, 
    10.1245755897274, 10.1279020000071, 10.0960513757605, 9.9342095496119, 
    9.75210413725438, 9.51916910596143, 9.28583055958591, 17.5759766493908, 
    17.5308647968256, 17.446880473973, 17.0695282737136, 16.8513995067693, 
    16.7712183224452, 16.6472073985642, 16.3394029868642, 16.2210850113693, 
    16.4841891197151, 16.3208725830661, 16.3609866748677, 16.1042533864607, 
    15.6212398855305, 15.3078202689421, 15.0828390257111, 15.0201714958667, 
    15.0132515771677, 14.3685934187337, 14.1306786817201, 13.5146637540786, 
    13.4309708712878, 13.5822474454241, 13.489979957779, 13.5569213685135, 
    13.5957340681602, 13.3897897945846, 12.6242228439315, 12.2395229085007, 
    12.1680263005458, 12.1187007833761, 11.9523134059249, 11.5773653942261, 
    11.4350899510696, 11.183059053567, 10.9914490881191, 10.9654584024814, 
    11.0943343090585, 11.3637463661935, 10.6942159810167, 10.4676583512504, 
    10.510451338114, 10.2002822982206, 9.79697669168673, 9.77857289109458, 
    10.0016710295989, 9.93580281738239, 9.9347555663498, 9.79323902422911, 
    9.53746673073291, 9.24668438583931, 17.5520506172291, 17.3918350595156, 
    17.1550565314307, 16.7252435967647, 16.5777388356364, 16.3869071534416, 
    16.3975295255228, 16.2871971736119, 16.2601065184296, 16.4024450800418, 
    16.1811384590682, 16.3113422657153, 16.1180514858214, 15.7697501328357, 
    15.5391569327823, 15.2071836874677, 15.2809336708045, 14.9462388839762, 
    14.1823571607038, 13.8960255628585, 13.5552036222961, 13.7371752924337, 
    13.7486495602256, 13.8258068685126, 13.5606004344484, 13.6364821450545, 
    13.4114071980589, 12.5190764741473, 12.1408471354666, 11.9232461452229, 
    11.9533298918555, 11.7579929829919, 11.5134305394477, 11.4872191630919, 
    11.3733883306148, 11.175436789319, 11.1368256669298, 11.4512629971678, 
    11.4540610979103, 10.4508645059479, 10.2506367531331, 10.3342681081302, 
    9.83600094635087, 9.34581468628399, 9.36876477674341, 9.52216361244451, 
    9.5574452641359, 9.57136099927503, 9.74300398935355, 9.38107790220169, 
    8.88290902864179, 17.5780320209499, 17.4693089124186, 17.0919836198028, 
    16.8451758629628, 16.7861732675779, 16.4141706913854, 16.3454896075671, 
    16.2537159064991, 16.2444931297322, 16.1166388933459, 16.0208530008347, 
    16.2662653635957, 16.1626401350816, 15.9166499310407, 15.7032890164091, 
    15.2875400767, 15.2585148450236, 14.0862698099653, 13.0287069415335, 
    13.1643615259436, 13.1738226752261, 13.3613448588691, 13.5163433614096, 
    13.7430940941262, 13.7552802806147, 13.3724149757173, 13.1215470611253, 
    12.0460863888764, 11.4369765389548, 11.4261197018678, 11.8388640132243, 
    11.7976028606874, 11.3335677863964, 11.3517235043126, 11.2064244075004, 
    11.1434005522748, 11.2597469797137, 11.4100063449116, 11.3990405250299, 
    10.4111079017337, 10.1145141558681, 9.98310914164656, 9.64011287945406, 
    9.3427161873037, 9.43617495750297, 9.39138261940255, 9.52525708427922, 
    9.57470463362313, 9.6082219547562, 9.36511325581372, 8.92029081414435, 
    17.6192232438717, 17.4995658003344, 17.2553001851915, 17.0727677685526, 
    17.0819199914851, 16.4761457972023, 16.1810400486006, 16.2034168538604, 
    16.0874851856225, 15.8113054638311, 15.9290142910094, 16.0505828797184, 
    16.12422186107, 15.9657102648792, 15.605833655553, 15.1118006528425, 
    14.4565342325828, 13.4528002584243, 12.7258791580845, 13.1109641695218, 
    13.1477451835754, 13.4816578544592, 13.4879061391502, 13.6798745248051, 
    13.7140511669554, 13.18636483182, 12.6736783413687, 11.5225011257983, 
    10.987126773006, 11.2179155557669, 11.4955360264755, 11.400707487424, 
    11.0718909410303, 10.8416711425735, 10.6582931049215, 10.6125062128378, 
    10.7428985632104, 11.0184303234895, 11.2573377720405, 10.4652163967639, 
    10.1385672266782, 9.89087957618312, 9.67883208101568, 9.57188265087556, 
    9.74025909286184, 9.48804633494063, 9.5155964884655, 9.53099715652797, 
    9.55892778500034, 9.4282090261298, 9.02484893220252, 17.7571637636958, 
    17.4586035369934, 17.2942684653617, 17.0593751807953, 17.1064405568828, 
    16.4782068704873, 16.1705148622131, 16.2207249971469, 15.9665530700481, 
    15.7142085798115, 15.8402829303981, 15.9094273241645, 15.9060455584418, 
    15.6470921374822, 15.0493847648545, 14.2379251261637, 13.5726962088134, 
    12.8056419486342, 12.7958345033328, 12.9890558708791, 13.2269783739779, 
    13.5376869829605, 13.4516069355937, 13.6756663819794, 13.6155503565305, 
    12.8376613404171, 12.0855767850114, 11.0955564285549, 11.2482688396142, 
    11.2061380337813, 11.2716551833136, 11.0743340633233, 10.9954368403663, 
    10.6811955509935, 10.5122978795224, 10.5828237997697, 10.6828818324684, 
    10.7389829927323, 11.1698757225206, 10.6611362189615, 10.3390366501642, 
    9.94789180898925, 9.76378695728107, 9.62509118100597, 9.91493179270365, 
    9.6961945769281, 9.49920890588736, 9.52077308899604, 9.48887191307827, 
    9.53416979530493, 9.40492184369244, 17.6456336575767, 17.5784977564498, 
    17.2953806711945, 17.3048719548974, 16.9750526271214, 16.5904564146484, 
    16.2001765345704, 16.2135594136309, 15.9168653254978, 15.7142109140028, 
    15.7074295070364, 15.6730900530987, 15.7036228526008, 15.6049277435495, 
    14.9577702937068, 13.9561991289017, 13.166554796106, 12.7895981525346, 
    12.7469951749935, 12.9648371682777, 13.2979879922219, 13.542983140916, 
    13.6043242751829, 13.7680305370157, 13.3547946426573, 12.4266162184916, 
    11.5915094188308, 11.1281903109677, 11.3814437158845, 11.4470048303212, 
    11.382656103523, 11.2801793511173, 11.0452304480389, 10.58030974211, 
    10.5237214732418, 10.5923566613671, 10.7744316585273, 10.9253107617298, 
    11.1777046575018, 10.8935212000699, 10.5219561542699, 10.2246880051837, 
    9.91816157612402, 9.83242373520534, 9.98131947891523, 9.90665961042119, 
    9.52667576151452, 9.50593563805962, 9.55935177406745, 9.48874994192647, 
    9.44535009116277, 17.7936042990752, 17.4921648335217, 17.5657398102161, 
    17.3243557477129, 17.0738983563605, 16.5534784900331, 16.3918215956852, 
    16.2924149695267, 15.9570587902205, 15.5512812820772, 15.2649375502921, 
    14.9682448379985, 14.954357128174, 15.1482514055768, 15.0305895183466, 
    14.176120582381, 13.1544557068157, 12.8084675696312, 12.7298661969984, 
    13.0835646256795, 13.4525618730732, 13.6217205093811, 13.7567462673495, 
    13.7759221430537, 13.0854323830487, 12.1028918974464, 11.413147460746, 
    11.3622709473274, 11.4342853530263, 11.5361338913703, 11.5063460700342, 
    11.3750216534911, 11.2171239485463, 10.8143879368725, 10.7503276400142, 
    10.5683852712921, 10.677564615275, 10.8744248423392, 11.0951851884143, 
    11.0119070888052, 10.6552181621949, 9.9892881292007, 9.99593742726899, 
    10.0227182122853, 9.97026201129322, 9.97151632921441, 9.57591902562365, 
    9.5175250721672, 9.46393219519053, 9.43638358966768, 9.4887762223327, 
    17.5603565769974, 17.7426906805316, 17.6473054297576, 17.5282104012193, 
    17.2740238490724, 16.8113907616845, 16.4062343237547, 16.0907672232321, 
    15.7698916639951, 15.2382279513468, 14.7139606301977, 14.1651386700824, 
    14.063019329026, 14.2737175522222, 14.3636038567766, 13.6928347076201, 
    12.9380871651644, 12.7288417195991, 12.7485421472043, 13.05267468618, 
    13.3892993243639, 13.6310777209177, 13.6323677911198, 13.4605547113012, 
    12.773714785709, 11.9406875897048, 11.3218705052562, 11.438608971643, 
    11.6345440143018, 11.5175096525585, 11.4442670070131, 11.491482853582, 
    11.3140984656469, 11.0637720140331, 10.9391228319547, 10.5429139062815, 
    10.643948470696, 10.7365941443523, 10.4518330468416, 10.7555930345548, 
    10.416313982468, 10.282701907598, 10.2172609378593, 10.1762549726414, 
    10.0581843297523, 10.0100858797213, 9.84038784330582, 9.50513978723419, 
    9.57720260707159, 9.38190430691448, 9.40998683599558, 17.4202101093716, 
    17.4710431188295, 17.4813932182629, 17.5544128459168, 17.3246331465772, 
    17.1467601706147, 16.6203513352048, 16.3229395680876, 15.7009096813619, 
    15.0958372383109, 14.6400171494821, 14.1502179133351, 13.8846029062237, 
    13.8453619550585, 13.7344160540681, 13.2856209111493, 12.7650481667963, 
    12.7456298782823, 12.7015896321226, 12.941528186568, 13.3827323279464, 
    13.2552923193853, 13.1560020877215, 12.9704623955824, 12.5710328394124, 
    11.9776330485438, 11.3569214609714, 11.572629085903, 11.9650451849942, 
    11.6847739391635, 11.3644485043987, 11.2415270416763, 11.0046231578608, 
    10.8525573272115, 10.551419879177, 10.3825508575367, 10.9463824965925, 
    10.8743058475793, 10.7497327468795, 10.550503718079, 10.2817616587052, 
    10.2886347421469, 10.0828784356274, 9.98806954017758, 9.8647507633472, 
    9.55235653989843, 9.7730588000405, 9.53485605095148, 9.59154063548007, 
    9.48783013565395, 9.39675647697101, 17.2643752606844, 17.3741307948362, 
    17.4696487323383, 17.5306899650498, 17.5629570981632, 17.2316443384781, 
    16.8652618282918, 16.302960930947, 15.5998977759886, 14.8527992744139, 
    14.4707074559283, 14.2190107170424, 14.0806505171923, 14.0318025948289, 
    13.7719199211099, 13.2425982071477, 12.7835998079123, 12.8353180686578, 
    12.5816541799919, 12.7360834288358, 13.1635677547383, 13.2279336294449, 
    13.1095234220489, 12.8825377012912, 12.4470591151684, 12.0898843724922, 
    11.5502701959285, 11.6987058703403, 12.0719290512762, 11.676342852792, 
    11.3452655308382, 11.3339549998513, 10.9282921726699, 10.4937970238154, 
    10.4009287048308, 10.5120696469325, 10.9506285002575, 10.8975895130367, 
    10.7485722469457, 10.48952336722, 10.3070491353886, 10.2610399218146, 
    9.94958522284063, 9.67502476051182, 9.74159115439995, 9.72813828513842, 
    9.69697429805031, 9.55076112434237, 9.73321153727514, 9.55507733138544, 
    9.42500775115694, 17.076888950623, 17.2545157908218, 17.2894199104215, 
    17.3492336888295, 17.514469699294, 17.43686653614, 16.7500578917171, 
    16.1851465844498, 15.3889151004912, 14.6100804857022, 14.3654813852804, 
    14.1977692815269, 14.1250640496913, 14.0809918228521, 13.8735524012563, 
    13.4593422135153, 13.0024638384934, 12.9726115472597, 12.4998114299264, 
    12.2823833237221, 12.5240841594476, 12.9487855137617, 13.0602562814339, 
    12.750002802925, 12.3254399830871, 11.6467152003307, 11.4298068390885, 
    11.8563235245806, 11.9073986285033, 11.430533722875, 11.3940100068746, 
    11.4959436982707, 11.4465668973604, 11.0152444816992, 11.1312090259604, 
    11.0753349833713, 10.9363644027814, 10.9563377723288, 10.7664167682877, 
    10.5450132314249, 10.4230975971258, 10.2260190109893, 10.059198713701, 
    9.85721495712447, 9.81899838406241, 9.81201736189396, 9.95174668926385, 
    9.87006113409127, 9.7924790312023, 9.60190943764371, 9.4494039693916, 
    16.8498477761548, 16.9972572031885, 17.1188322368153, 17.2127849459617, 
    17.3639030966896, 16.9474124641567, 16.6791805869692, 16.0166079437303, 
    15.3005897653935, 14.571281596082, 14.4266280973565, 14.444684453304, 
    14.0465820423932, 14.0701972705177, 13.956710149456, 13.5176074551393, 
    13.1416632327615, 13.1272954260051, 12.5152781577732, 12.071757380637, 
    12.0695932926091, 12.5209905265477, 13.1299153655296, 12.8572222857585, 
    12.5587126259456, 12.055084162032, 12.2296421080792, 11.6995120817589, 
    11.5296222005492, 11.3042942446991, 11.3625836857673, 11.5096892915944, 
    11.4071828430594, 11.456142980229, 11.4238853192332, 11.0017556110604, 
    10.7531083524444, 10.7723812445596, 10.8346541189536, 10.6484403183141, 
    10.5217526288586, 10.3110499712216, 10.1107397063421, 10.0961194359727, 
    9.96347279877204, 9.80600427183173, 9.81859829304815, 9.92444939753934, 
    9.81975798401888, 9.71799629852526, 9.51923227324718, 16.595454633755, 
    16.5510899676896, 16.4963874450148, 16.7278954885397, 16.9630093283267, 
    17.0763058847409, 16.6594390525623, 16.0124505796897, 15.3914293058262, 
    14.9645898002077, 14.7125309926502, 14.4418543354804, 14.0546901241387, 
    14.0700567974855, 14.1713825755306, 13.5309844753491, 13.2039918961678, 
    13.0660383137931, 12.4500463493652, 12.3863541797655, 12.1531396344946, 
    12.2542972616177, 12.8628799321312, 12.6955783410287, 12.2163487472153, 
    12.0216259604027, 11.8718192862037, 11.3980437204871, 11.5414081176667, 
    11.3868483799413, 11.4090825045161, 11.3737900771854, 11.2737861997608, 
    11.3435229136571, 11.1006631084111, 10.8286328217526, 10.5912910043014, 
    10.6577247626404, 10.7372699651785, 10.6373539632077, 10.5003605876131, 
    10.4011373032887, 10.1142685286414, 10.0303666989351, 9.8571687763391, 
    9.82336627477529, 9.82168908917645, 9.83524944107073, 9.78903222162201, 
    16.4783972654872, 16.3565933058254, 16.136867909863, 16.3417473275331, 
    16.5769885436203, 16.6807389882897, 16.435221094116, 16.1750505153208, 
    15.6740189060021, 15.5024550356693, 15.2625398563914, 14.526984758344, 
    14.0024219855165, 13.8826635769441, 14.0201102836504, 13.4263542788573, 
    13.1327346203569, 12.8485038509532, 12.6192365546387, 12.7250243159195, 
    12.3976197153637, 12.0299519780436, 12.0950564368237, 12.5920133727539, 
    12.5402694797385, 11.9913930332071, 11.4951165144751, 11.3229966156614, 
    11.3591546987314, 11.3619552132802, 11.3007714685267, 11.2513413816965, 
    10.8839935270302, 11.0739073471378, 10.5550690404606, 10.6452711829384, 
    10.6414688141313, 10.7916525576013, 10.7665044236196, 10.5720587911759, 
    10.4468741962972, 10.4109526621156, 10.3010813556808, 10.2073417833287, 
    9.86293463994062, 10.1993021803036, 9.91743473514918, 9.90624190480227, 
    9.92093991541031, 9.8449542606181, 9.78517238070612, 16.2429291083023, 
    16.0780523411531, 16.0934808165837, 16.0159633252339, 16.0605708416515, 
    16.3804780658112, 16.569524471618, 16.3097798660322, 16.0092118335631, 
    15.9003458931985, 15.7665333754242, 14.7315592171058, 13.6778848334661, 
    13.7195010026689, 13.8065628784527, 13.3892201790594, 13.1822373471738, 
    12.8639528399532, 12.8984779733832, 13.0788891256862, 12.7238759818099, 
    12.1903384248954, 11.9051617890993, 12.0454244943336, 12.3061176246087, 
    12.1362334755852, 11.6492554221029, 11.3202763071695, 11.4136247760247, 
    11.3841240990038, 11.2403269995997, 11.0218586970291, 10.8299685677634, 
    10.7790749531124, 10.6804223450354, 10.7443859634595, 10.2457829242402, 
    10.4728242023009, 10.4066704927409, 10.2435262518944, 10.2303932263459, 
    10.2329540998739, 10.1904569500649, 10.0047240353471, 9.88375261942033, 
    9.84678217720741, 9.60595214543235, 9.3459082060531, 16.3858791774233, 
    16.5363822379334, 16.3532619011012, 16.153835883561, 15.9823009404615, 
    15.9868652883885, 16.3437298206259, 16.5285740673638, 16.3614196580632, 
    16.1077892331531, 15.3982962425593, 14.1566332120803, 13.4402373450748, 
    13.4795322754475, 13.5893044250819, 13.499646958047, 13.1981059785916, 
    12.9881973725514, 13.0941544174431, 13.1246752986124, 12.7785704435919, 
    12.3863322783566, 12.0601257839486, 11.9840063658904, 12.2381254567239, 
    12.0408423244924, 11.7242442499229, 11.5703866065894, 11.5343924987472, 
    11.0865796603903, 10.9080192440392, 10.8270044394372, 10.7909521973134, 
    10.6185364798737, 9.82283732960778, 10.1152168101094, 10.027235448453, 
    10.1742104139306, 10.0097947260226, 9.93007361798728, 9.68588458601979, 
    9.38986781582929, 9.04784075272255, 8.90748941171513, 16.6754731397834, 
    16.5360272328101, 16.5091414066185, 16.429894009947, 16.2112698760754, 
    16.1730187817779, 16.3932174562584, 16.5144881953504, 16.4583360081264, 
    15.9272000338887, 14.9055618418622, 13.8027985267868, 13.2727326887681, 
    13.3030270331279, 13.3413287867579, 13.3760226172904, 13.2185114994201, 
    13.2176689078487, 13.0803870031304, 12.9081434547236, 12.6452662525272, 
    12.3315679766749, 11.8046701786111, 11.8781756111259, 12.0346659548377, 
    12.1690618913694, 11.9715309539705, 11.8380156896662, 9.8634204623732, 
    9.6628609473464, 9.49684298429912, 8.76991317849824, 16.6866311674386, 
    16.4883329012023, 16.4345095289295, 16.3546037651826, 16.1657445476969, 
    16.0757340007177, 16.2245737653534, 16.0957060495771, 15.7148150553623, 
    14.9725219596127, 14.4692878673885, 13.6886665269464, 13.3929781041333, 
    13.354129692385, 13.1653583784506, 13.1180595712946, 13.2487767030733, 
    13.2187346780419, 13.0427517328519, 12.7494571860074, 12.7266041433038, 
    12.2878065124034, 11.9729323881387, 11.8230765193232, 11.7185483915482, 
    16.6362916811415, 16.3403436404168, 16.2052568441374, 16.1509821328953, 
    15.828361365386, 15.5353168064013, 15.0551710879584, 14.4283841744058, 
    13.8766590449267, 13.7764553874226, 14.0029084802899, 13.6416495717376, 
    13.5829799370059, 13.480424459476, 13.1708651701833, 12.9636386740451, 
    13.0976356871188, 13.1430603931375, 12.7953115663409, 12.6982612163861, 
    12.6869299308085, 12.3829604390326, 12.064700424688, 12.032126064156, 
    16.599839753818, 16.2932434078296, 16.177721838006, 15.7969183722763, 
    15.2836251489947, 14.9093639295333, 14.2754845869247, 13.6832371598593, 
    13.4764184938837, 13.701913395141, 13.7415449512542, 13.4864546015892, 
    13.7115378322053, 13.441547666169, 13.0967374535624, 12.9286753748168, 
    13.1033750374573, 12.926715970417, 12.4997884953005, 12.4567732999038, 
    12.6043591852848, 12.4249195735458, 16.3495460498458, 16.2068516882272, 
    16.2664324414935, 15.5277716701979, 14.9762550562352, 14.4145622436438, 
    13.8956115532902, 13.5587403027113, 13.5627268882371, 13.7673984882492, 
    13.6907108926756, 13.6926024255343, 13.4216195172909, 13.2864995181179, 
    12.9902010721397, 12.8333388158758, 12.9208464648711, 12.5625979737977, 
    12.2806904378038, 12.4212108797843, 12.3495930964001, 12.1356520680349, 
    16.0458645433269, 16.2371096691375, 16.3488674374741, 15.9193805246194, 
    15.1490220315736, 14.3079824895461, 13.6965040971987, 13.5348710405634, 
    13.6218427271189, 13.8291871537175, 13.69595812518, 13.2927969581881, 
    13.2740564773624, 13.1577833876742, 12.9361602119151, 12.7945199021004, 
    12.883416926562, 12.3709508778389, 12.2037293962206, 12.3311145600151, 
    16.0238019055509, 16.2517632446187, 16.2875756013625, 16.3122995985891, 
    15.5718237318991, 14.5784241723228, 13.7010742144895, 13.6566649183453, 
    13.7013739634431, 13.7987287682334, 13.7034151244929, 13.4902504462733, 
    13.3118797395846, 13.091753017435, 12.8749312317479, 12.8554357667255, 
    12.8771040071868, 12.7381476025169, 12.3882646651594, 16.0421621021165, 
    16.230028537928, 16.123736737303, 16.1848766176304, 15.9104115918868, 
    14.9351442235869, 13.9772765326784, 13.9244467234406, 13.8456674107053, 
    13.7784269455732, 13.945148866856, 13.742428383227, 13.3847532097465, 
    13.302214915048, 12.9366983654067, 12.7316143228278, 12.8460645693864, 
    15.7777694865521, 15.8411505384898, 15.8854520556104, 15.9907830075667, 
    16.2973496705103, 15.4271291705912, 14.3664564054934, 14.1980014369123, 
    14.3564564146259, 14.3035743964499, 14.1269220336557, 14.0130482723677, 
    13.8611957858388, 13.5798915354705, 13.3601395465763, 12.9396772535591, 
    15.7581300178104, 15.6023722458135, 15.6235942520917, 15.7638893679516, 
    16.140844503488, 15.7261249344292, 14.717883674119, 14.5162724984865, 
    14.8491418962931, 14.4657289989278, 14.3076235721774, 14.1601936277164, 
    13.4571941824864, 13.4419036498682, 13.362252908521, 15.7532242517714, 
    15.6113138984563, 15.6613449223337, 15.6382884608572, 16.0655645169972, 
    15.7605691342392, 15.0557681414851, 14.7677628254106, 14.7798860568887, 
    14.0740266497678, 13.9702765008677, 13.7218200253012, 13.3341627220993, 
    13.2558648029076, 16.1046132963634, 16.0587015775681, 15.859718064158, 
    15.5921656027558, 16.045667833077, 15.9658173276441, 15.2605745793514, 
    15.0737420268304, 14.5318375212358, 13.7540298786381, 13.4940451517382, 
    13.4278537750748, 16.3090341823811, 16.3501313598741, 15.9562924660575, 
    15.4268710149764, 15.7496021139885, 15.8896614075549, 15.3046346333405, 
    14.8663741745206, 14.2327507455465, 13.6968225290846, 13.575463213427, 
    13.5109709332598, 16.2930893309188, 16.3235463412034, 15.7859568910011, 
    15.3349115748339, 15.4637785298152, 15.4659151083743, 14.9971339924135, 
    14.5638114711006, 14.2168129999791, 13.6746055974307, 13.6770914637504, 
    13.7179286080639, 16.4803749127748, 16.0936567279166, 15.5807064297095, 
    15.6733630765052, 15.5380225258205, 14.9889387753678, 14.6823396103953, 
    14.4066910382741, 14.2855541932963, 13.9719286110123, 13.7721826221782, 
    16.3374846993252, 15.765483597213, 15.5447499081975, 15.9657515960408, 
    15.8298358616152, 14.9594828489515, 14.5503686907173, 14.5499448703732, 
    14.6180518993415, 14.2123302489648, 13.8784210321689, 15.8590851760722, 
    15.463058076629, 15.5906422674032, 15.7549675713184, 15.412843922415, 
    14.9231822544076, 14.4933029574651, 14.4689335748436, 14.329427097054, 
    14.0473235892928, 13.734058362603, 15.5706036796874, 15.2987990538596, 
    15.1628833679763, 14.9535960642614, 14.9504506906428, 14.7297703179157, 
    14.6270715057878, 14.2956631462144, 14.2146178056826, 14.0742182810208, 
    15.6474476734682, 15.4045620801293, 15.3211111725307, 15.1063496337754, 
    14.7807261940745, 14.8002465535796, 14.782250481285, 14.5228956980648, 
    14.3708128634878, 15.9192055397658, 15.5510812740254, 15.5224126656366, 
    15.102324324387, 14.7875744373369, 14.5491636424701, 14.5202439689001, 
    14.6509321690057, 14.5356829523937, 16.1648906818186, 15.7617310550611, 
    15.7000168182608, 15.5848114420693, 15.1547037457204, 14.6858792951263, 
    14.2586786395657, 14.3840822659501, 16.0754439053485, 15.8427560985297, 
    15.6134696720077, 15.3948625906094, 15.2440331786457, 16.0080979129131, 
    15.6688659457742, 15.0798307616011, 14.9614987301552, 13.4754975940026, 
    13.4967701858408, 13.4387779613822, 12.8534528079167, 9.97312003611153, 
    8.53539415894808, 7.88309474387969, 7.27760601293366, 5.85047641457708, 
    5.14333016023509, 4.53900047008456, 3.93551214930784, 3.39660876594238, 
    2.98468177046345, 2.6392801989193, 2.34565017369255, 2.13970772541042, 
    11.6954597242306, 6.66734708998324, 32.3522623632796, 32.3514008238056, 
    32.3613573739676, 32.4297467475598, 32.9237525497239, 33.5136765935476, 
    33.8586707231655, 34.0168448269664, 34.1135818379451, 34.2079610459339, 
    34.303153042507, 34.3893840865968, 34.4559506768072, 34.5000670163041, 
    34.5357248263515, 34.565073042324, 34.5847832888809, 32.5769910982372, 
    34.0583413958089, 12.5665905319167, 12.6138845288356, 12.6811343038373, 
    12.3855463704015, 11.1399621594296, 8.93940299971363, 7.9013942176856, 
    7.3876659507936, 6.95298705404669, 6.31874732459739, 5.42408361745676, 
    4.87005946838081, 4.39327208811808, 3.8657686612582, 3.36421996848644, 
    2.99007090238006, 2.6870225113931, 2.41261654025156, 2.14698200554632, 
    2.01953224689918, 32.4764081119144, 32.4778341884801, 32.4915941239632, 
    32.5456733244945, 32.6925528868204, 33.0966287090027, 33.5935541480676, 
    33.8297110845854, 33.9402230282634, 34.0091483221786, 34.0699542193124, 
    34.1477993660771, 34.2515604353705, 34.369914135477, 34.4573565359771, 
    34.5000174907463, 34.5306657130524, 34.5580920210935, 34.581732973612, 
    34.5927782106655, 17.6449306368776, 17.4554283946941, 17.2371170554078, 
    17.0184862335564, 17.2931912347184, 16.9752200988574, 16.72748019298, 
    16.3650963354689, 16.3454183285978, 16.3724356278229, 16.2967737682435, 
    16.2277005391416, 16.0338515645295, 15.6230813667865, 14.7294947052889, 
    14.7552328829298, 14.5618684203666, 14.5527837833449, 14.3091857415309, 
    13.5665961994293, 13.0896932052982, 13.3155367871616, 13.0931846373074, 
    12.9896002287281, 13.0596579016274, 13.2955583129472, 13.5884152331874, 
    13.4208471382869, 12.8293833672674, 12.3567969959774, 12.5734439660965, 
    12.8726839200308, 12.3775004246475, 11.2882209901632, 11.0446191896783, 
    11.0415979355078, 10.7726416772719, 10.8384736617661, 10.9848097963424, 
    11.006187937415, 10.7303782935642, 10.6179993848928, 10.4252855978676, 
    10.2844903078126, 10.1859975784984, 9.94942763211012, 9.93805346386368, 
    9.71488024376766, 9.58793571658805, 9.49922035912191, 9.07052343015194, 
    17.6170090042779, 17.5595670187386, 17.3175798869051, 17.291362846593, 
    17.1140461251531, 17.0121555762669, 16.7410830077041, 16.2990329837383, 
    16.1931659838708, 16.3613165382468, 16.2279577162972, 16.1632129279946, 
    16.0088402282396, 15.5466569684498, 14.785536992815, 14.7412603869493, 
    14.4874650041307, 14.6241314200997, 14.442534495525, 13.7109900130852, 
    13.3539036472218, 13.4623852056311, 13.2852139025491, 12.9575316015902, 
    13.1967194931504, 13.440392593928, 13.5683686657255, 12.839993435203, 
    12.2753681431851, 12.3161761967368, 12.405267914494, 12.2286074430781, 
    11.572952884969, 11.1377775676197, 11.0291987563448, 10.9174798519076, 
    10.7523631710655, 10.8328476975079, 11.0801099618165, 10.9226996599017, 
    10.6528772065034, 10.5890483041966, 10.3668923027989, 10.066070792918, 
    9.96008803154168, 9.99016538893277, 9.92714182129559, 9.77183102486106, 
    9.58508047775104, 9.41987804541286, 9.1779727325129, 17.4729440632671, 
    17.4381762027697, 17.3545323982621, 16.9351439561322, 16.6876404756342, 
    16.6557307131607, 16.5826861052107, 16.2080792128924, 16.0682593653113, 
    16.3167164516728, 16.1289462580164, 16.211423883093, 15.9849769733994, 
    15.4742711748869, 15.0849152339312, 14.9181659707721, 14.905010958715, 
    14.9188126016564, 14.2640318232416, 13.9158770870261, 13.5262217446801, 
    13.3520642235887, 13.4672672824353, 13.3912644858166, 13.452890407039, 
    13.5038786388308, 13.1764242676163, 12.3941701981251, 12.0754460117311, 
    12.0458317062902, 12.038310253003, 11.8288382178965, 11.4397459556109, 
    11.3555094173364, 11.0763789401436, 10.8926498290401, 10.8064757703145, 
    10.923942222868, 11.2460597327393, 10.5370989219283, 10.3266929958781, 
    10.3829389667311, 10.0349153237607, 9.61275233020481, 9.61341703151845, 
    9.84452547836339, 9.7788931233268, 9.80368702716045, 9.62450928830696, 
    9.38162762284223, 9.10970044585114, 17.432287026894, 17.2744416902527, 
    17.0825172869208, 16.6124832233359, 16.4843207475675, 16.256238500248, 
    16.2632876144951, 16.1474870510015, 16.1180361248064, 16.2262817355919, 
    15.978589463597, 16.159370497069, 15.9803794565991, 15.5919866735745, 
    15.3457617954155, 15.0533795407275, 15.1280128996147, 14.6702684029926, 
    13.9859756008143, 13.8521315921156, 13.4914685686075, 13.514123905551, 
    13.5747958869979, 13.6726858652504, 13.4725411734905, 13.511835300626, 
    13.1567544555827, 12.2810059636007, 11.9024642921509, 11.7433765404188, 
    11.8375742476722, 11.6613888151517, 11.4034495908582, 11.3639956502679, 
    11.2205412926235, 11.017954085647, 10.9743577312757, 11.2781895539107, 
    11.3123087815152, 10.3041464157639, 10.1385185947816, 10.2232816979991, 
    9.70488789696469, 9.19000942577757, 9.2683999753068, 9.36229804077171, 
    9.42220782640002, 9.44083531632099, 9.59948108675316, 9.17613961534544, 
    8.73404915142206, 17.4562631213909, 17.3449551964948, 16.9759810023529, 
    16.7660075805825, 16.7105182623027, 16.2727868155892, 16.2073494950229, 
    16.1065854770781, 16.0602336059837, 15.9031652761776, 15.8466800276356, 
    16.1310113684457, 16.0134392596568, 15.7180267139892, 15.5381974975201, 
    15.1555199125215, 15.0475490359556, 13.7289742460446, 12.9741277884154, 
    13.1018647901452, 13.085942752237, 13.2243360401685, 13.3247037380437, 
    13.5929018938533, 13.6299131356132, 13.25976297742, 12.9187244603509, 
    11.7708972419212, 11.2311392401649, 11.299132837497, 11.7338630600031, 
    11.6635353919225, 11.2359341889667, 11.2230384944496, 11.0658054063426, 
    10.9696044520381, 11.1048247842787, 11.2436196111648, 11.2821103652521, 
    10.3043680966186, 9.97945694231469, 9.84110484666558, 9.51307845231747, 
    9.24084902162734, 9.38949147323626, 9.30767029643764, 9.41149159919121, 
    9.46704970797896, 9.41335875950137, 9.10781377031785, 8.7866191245996, 
    17.5341649778878, 17.3889780709429, 17.1372779641784, 16.9686691049332, 
    16.9861336403274, 16.3249031882694, 16.0440823415304, 16.0603656860477, 
    15.9099371928282, 15.6382389424387, 15.7906568289533, 15.9202306820706, 
    16.0280822047013, 15.8210153446275, 15.5082394731785, 15.0822499816846, 
    14.5096784112341, 13.2903662711447, 12.6895899742819, 12.9855348658516, 
    13.1004897083364, 13.3814901343, 13.3539325595153, 13.5451337329288, 
    13.5735891280357, 13.0770769621628, 12.5246977654772, 11.3465752865167, 
    10.9330594023262, 11.0755028361353, 11.354249049193, 11.3373750489679, 
    10.9213726184173, 10.6859091341336, 10.5055280328962, 10.4811247484876, 
    10.6298810428683, 10.8741860962278, 11.1308627299156, 10.3310847636032, 
    10.0006770155593, 9.73602516211026, 9.52405586659371, 9.45818814505458, 
    9.63045851797898, 9.39134865624813, 9.4036409573707, 9.46940309167273, 
    9.36276890268669, 9.17031704494432, 8.84991584927105, 17.6477239915229, 
    17.3627412481234, 17.170312955925, 16.9557420132286, 17.0012950796708, 
    16.3336937550671, 16.0430162064465, 16.0523299116622, 15.7837731775831, 
    15.5828557023896, 15.6928579648028, 15.7567194820583, 15.7647723319728, 
    15.4941863509838, 14.8452750741426, 14.1744718481322, 13.65376679391, 
    12.803541559794, 12.6926310914708, 12.8125265663837, 13.123647509443, 
    13.3823470694235, 13.3176818600555, 13.5061487170851, 13.4594610858309, 
    12.6665920120797, 11.93308501069, 10.9380627991507, 11.2502341962831, 
    11.123910030542, 11.1387838881587, 10.9920405993431, 10.8591839074809, 
    10.532926856411, 10.3988476516015, 10.4972615513708, 10.6336214048065, 
    10.6735002677208, 11.0312584994194, 10.4986541663734, 10.2085872990891, 
    9.81116817790274, 9.59796976286602, 9.48563261274131, 9.75910594418317, 
    9.56673378583383, 9.3516692175608, 9.40197529682259, 9.36850975684515, 
    9.34905861889289, 9.20025680638853, 17.5432259894007, 17.4833672755516, 
    17.1969444744611, 17.2064315693308, 16.8928541674493, 16.4478794974651, 
    16.0892250056173, 16.0441015954246, 15.7564779739653, 15.5838488604397, 
    15.4983837034295, 15.4798417255617, 15.5615662388918, 15.4625028815782, 
    14.6832295152519, 13.6925151329508, 13.0580820593589, 12.6039779835956, 
    12.635562681232, 12.8820185890217, 13.2274830032129, 13.4039349063982, 
    13.4506244674418, 13.5966424390125, 13.1657449124952, 12.1852691405925, 
    11.4833718417736, 11.141304670277, 11.332208393667, 11.3788638815274, 
    11.30976140665, 11.1240701010725, 10.9142359008694, 10.4560013126296, 
    10.4206323814566, 10.4829363271612, 10.6670264607277, 10.8342484233723, 
    11.0409129894102, 10.7533350535012, 10.4230245870583, 10.1123890045365, 
    9.76421743938232, 9.65969275945747, 9.81737035474801, 9.75666256220584, 
    9.36138800686927, 9.37717019060051, 9.39685487057947, 9.30675458516381, 
    9.26869667281649, 17.6604370009696, 17.4285683209705, 17.4409860097011, 
    17.2410168307679, 17.0119884174663, 16.4799594581686, 16.2848262455642, 
    16.1537809224009, 15.8036691332418, 15.3544849140222, 14.925312775247, 
    14.6602164733496, 14.7824464979344, 15.0556279498376, 14.8527752116106, 
    14.059248199856, 13.049204047429, 12.6737799296486, 12.6282630766117, 
    12.9752486162268, 13.3687412945606, 13.520722373642, 13.6217526985317, 
    13.6345610280215, 12.9061511995001, 11.9190278185632, 11.3066018320295, 
    11.2927958409259, 11.4007911497214, 11.423685927315, 11.3878693928336, 
    11.2581070282438, 11.115100967031, 10.7003184991699, 10.6261872570049, 
    10.4527128786228, 10.5398886992838, 10.7460318824002, 11.0206094179213, 
    10.9057005064445, 10.5680364705019, 9.90727632686272, 9.83864670610916, 
    9.86140423890458, 9.81715752011179, 9.82047089181178, 9.45997226969792, 
    9.37819145004051, 9.32181207159284, 9.25835196108855, 9.30987099337354, 
    17.4085172959521, 17.587294847104, 17.5554033318571, 17.4364106340907, 
    17.1997779673057, 16.7121152430586, 16.3033783117331, 15.9610535750502, 
    15.6466127778255, 14.9872079953997, 14.3225608698601, 13.9036587659667, 
    13.9478868601246, 14.1716374162662, 14.2929551591532, 13.6778051747908, 
    12.8556070727193, 12.6335119783734, 12.6284108399405, 12.9642348171202, 
    13.3335343558642, 13.5364835975121, 13.5388843854509, 13.3843386720888, 
    12.6439101658582, 11.7907828828247, 11.2039946161859, 11.3001879507493, 
    11.6619110934808, 11.482336928271, 11.330671365764, 11.3529899037435, 
    11.2008346466769, 10.9463307260694, 10.8271987125528, 10.4188749288387, 
    10.5987312201498, 10.6301219492941, 10.4213503803788, 10.6457780648398, 
    10.3256829487377, 10.1689533046444, 10.0562192143218, 10.0210837864923, 
    9.91506243673416, 9.82609002348442, 9.66308738123443, 9.37182322914273, 
    9.4088642530501, 9.22263520506783, 9.20981689869164, 17.2781101133571, 
    17.3355421858715, 17.3753376541067, 17.4345121482492, 17.2377271514269, 
    17.0433370986338, 16.5277072838403, 16.2030191033993, 15.5754167651111, 
    14.9530429747088, 14.406806001916, 13.9609845332389, 13.7910757255419, 
    13.7295529400338, 13.6183360990646, 13.1802978283309, 12.6742208646909, 
    12.6462551500184, 12.5687303654175, 12.8641675585276, 13.2339803920342, 
    13.0763328804682, 13.0298134869525, 12.8898056299449, 12.4934879880087, 
    11.8140790549571, 11.2639324167119, 11.4234128994772, 11.8795543433169, 
    11.5820683813892, 11.2067011394615, 11.0539560969256, 10.8407773187859, 
    10.7319863463911, 10.4428404112584, 10.2448751850101, 10.7968902176206, 
    10.7832487619822, 10.6345524216859, 10.4141179806707, 10.145957537842, 
    10.1332748562734, 9.89754724935808, 9.7707379075983, 9.70977480700742, 
    9.43289960208984, 9.61679356479426, 9.35476615131042, 9.41663532873484, 
    9.31731220688824, 9.23232333953975, 17.117684604244, 17.3008771636467, 
    17.3426908519937, 17.3855933079504, 17.4944535961666, 17.1507241482521, 
    16.7441243944054, 16.2546728594123, 15.4780743466585, 14.7829896969145, 
    14.4053024839539, 14.1171930921436, 14.003160289934, 13.950728700078, 
    13.6659431438972, 13.0880959351891, 12.6585872723247, 12.7150441062522, 
    12.4529534946178, 12.6165062369908, 13.0008160687238, 13.0355810888628, 
    12.9060715101467, 12.7070658862238, 12.3853181862034, 12.0125881964129, 
    11.4959891106188, 11.5407828099101, 11.8702236609294, 11.5249020284835, 
    11.2052635959784, 11.1848140239654, 10.7375396626547, 10.3577070138248, 
    10.2853253935721, 10.4024784131372, 10.7934029255279, 10.7820726237084, 
    10.603863796609, 10.3151554117879, 10.1614345237889, 10.0801134113838, 
    9.76056594986296, 9.55051308005385, 9.62220408282935, 9.55237311294674, 
    9.51332574591703, 9.37850265130981, 9.54139439565009, 9.36304800547011, 
    9.2579756331346, 16.9575188950537, 17.164085553736, 17.1561242061527, 
    17.2220686774401, 17.4198589599655, 17.3143015812708, 16.6352325511929, 
    16.0767648769666, 15.2118081267214, 14.4904113436919, 14.2708069558917, 
    14.1253329321628, 13.9982063292732, 13.9813593028568, 13.7882979600085, 
    13.3165545156544, 12.9067714830068, 12.8545728435956, 12.3483149519359, 
    12.1358004988893, 12.4258686982291, 12.7767435868542, 12.8769699854575, 
    12.6002516609738, 12.2092006007172, 11.7824294293452, 11.3594897708579, 
    11.6712604749151, 11.7287365347043, 11.2836169171146, 11.2726144972655, 
    11.34005534708, 11.3353582718913, 10.8482611921364, 10.9930850514633, 
    10.9443991172715, 10.8105157611935, 10.8335810168345, 10.6626266269667, 
    10.4064559674661, 10.2765510261738, 10.0753019257684, 9.92032160619785, 
    9.76265620608726, 9.70325369504203, 9.68623461851669, 9.78271805308506, 
    9.64227512109723, 9.60531665277975, 9.45092282987618, 9.27731426939823, 
    16.7280445866022, 16.8920349192481, 16.9224347049519, 17.0503018415276, 
    17.2670786838124, 16.8537083284216, 16.4923707190739, 15.8272850425421, 
    15.0507438282019, 14.4331540731405, 14.2740164017154, 14.290916487311, 
    13.9456757762913, 13.9536122612442, 13.8578422418414, 13.446648735468, 
    13.0669125031041, 13.0101573365716, 12.42538254091, 11.9451191769475, 
    11.9518155288035, 12.4305985233182, 13.0270298777985, 12.706102066935, 
    12.3259412977732, 11.7970597650325, 12.0304945599909, 11.5597117191702, 
    11.4141485531531, 11.182645627076, 11.2649995326213, 11.4358056600942, 
    11.2816705888198, 11.3161980630224, 11.2876991154072, 10.8540205661176, 
    10.6009405172033, 10.6312279058295, 10.720578140797, 10.5261717909434, 
    10.3701070117811, 10.1630209492041, 9.97196461887966, 9.9401961726262, 
    9.79145613370742, 9.63863263502883, 9.62809790855399, 9.72082314265375, 
    9.63110624976146, 9.50771079787995, 9.36024852485785, 16.4456665973945, 
    16.3796059776458, 16.3091952174318, 16.5460434335139, 16.8475143138318, 
    16.9364423736106, 16.5309566485133, 15.8059213885124, 15.1975442048548, 
    14.9086186813697, 14.6269869203543, 14.3243070261306, 13.9381480422972, 
    13.9278724137831, 14.0492373580196, 13.440184168303, 13.0839606611569, 
    12.9486446821555, 12.3660429457293, 12.2451134753804, 12.0479110036638, 
    12.1469115138668, 12.6956834564894, 12.5111227604366, 12.1159169776259, 
    11.8657024578749, 11.7823035162764, 11.2603678980172, 11.4330419152695, 
    11.266645687127, 11.2942816234492, 11.3059309672217, 11.098894307919, 
    11.1942645954073, 10.9517649080651, 10.6753523313334, 10.4881839374953, 
    10.5388858436147, 10.6234615259914, 10.5122268153891, 10.3567651281277, 
    10.2457557793557, 9.91082352418514, 9.81937975666681, 9.70114874754052, 
    9.60679449454909, 9.59735185038634, 9.64693287075104, 9.62662882513267, 
    16.3260677180524, 16.1551299870347, 16.0237722899532, 16.1822958466869, 
    16.4090017461837, 16.5487256778326, 16.378192563719, 16.0246129117596, 
    15.5218733422843, 15.4437823153683, 15.2649964659507, 14.4906981739699, 
    13.8488172184073, 13.7285976838661, 13.8440233640615, 13.3019766697862, 
    12.9862983778083, 12.742372633185, 12.5004736569668, 12.6451952441619, 
    12.3239810616037, 11.9152554594682, 12.0603647981535, 12.4674585250494, 
    12.3909706305055, 11.8994521497813, 11.4541747739571, 11.1954683320665, 
    11.2259390057689, 11.2590141781063, 11.1670823468905, 11.112936477431, 
    10.7377230514722, 10.9483348613483, 10.439223003847, 10.5047702787238, 
    10.5575025716414, 10.6473346846776, 10.5933182013135, 10.4332547070218, 
    10.3134855109376, 10.2601578520719, 10.1389181992917, 9.99896183736892, 
    9.74846257512394, 9.99581951270767, 9.7060271851585, 9.67884681234942, 
    9.70225072248525, 9.61661915769505, 9.53323911124125, 16.0825317531522, 
    16.0191145418696, 15.9836072689609, 15.8822039534452, 15.9582056623458, 
    16.2668862292989, 16.4620163349211, 16.2312493047277, 15.882302118677, 
    15.7978496108211, 15.6915311898067, 14.6915092319276, 13.5226405554203, 
    13.6067631315755, 13.6377552949383, 13.2508731869707, 12.9856548367711, 
    12.7107577494864, 12.7559310532963, 12.9093653668128, 12.5839411962656, 
    12.1093626806253, 11.8296691721153, 11.8821653673236, 12.1631751681176, 
    11.9803671116894, 11.5710741225233, 11.3152937940576, 11.350154565058, 
    11.2987212825037, 11.0920815306505, 10.825378970201, 10.6991329182773, 
    10.646654421912, 10.651163402558, 10.6988014732446, 10.214116719204, 
    10.3794993887525, 10.2918282745937, 10.1293894895653, 10.0316980505349, 
    10.0245906162237, 9.97396063546777, 9.80538684358117, 9.6574142559845, 
    9.5600778455979, 9.35456341429227, 9.06706429301087, 16.2867626609295, 
    16.4508534684185, 16.2563238672468, 16.0843604663829, 15.9461720663527, 
    15.9622563029964, 16.2421708407996, 16.3961912285755, 16.2222089173104, 
    16.0410122895008, 15.3386648905497, 14.0737053528853, 13.2920751234304, 
    13.3546656148311, 13.4616159644375, 13.3250498328603, 13.066782361039, 
    12.8447785319792, 12.9081349649316, 12.9696278246242, 12.6695084639943, 
    12.2522845002609, 11.897196645696, 11.8595725057573, 12.1413225823548, 
    11.9035114826697, 11.5621454117, 11.5419589725238, 11.4524072814604, 
    11.0181648068339, 10.8332067651259, 10.7729702097459, 10.7573446276107, 
    10.6054937799241, 9.74490181904149, 9.98376552661876, 9.8571597222842, 
    9.96432692359831, 9.74660212656276, 9.59408478973653, 9.42606290951092, 
    9.04252642549548, 8.72168760198169, 8.57997607710683, 16.5587625557699, 
    16.4227159350211, 16.3838056310574, 16.3356660022506, 16.1753112088392, 
    16.107753805274, 16.3181617206431, 16.4512030393249, 16.4018439415654, 
    15.8665841415054, 14.7820103141129, 13.6728831098325, 13.1720675282098, 
    13.1810053659799, 13.1764818243849, 13.2296441270979, 13.0634347013447, 
    13.0859839846188, 12.9632850667893, 12.786689680106, 12.5642609800848, 
    12.2396863841113, 11.699941781852, 11.763981694217, 11.9331773007135, 
    11.9674467349588, 11.9266331900507, 11.7550948301887, 9.75066969941403, 
    9.47514788400987, 9.22826150331098, 8.46844255054616, 16.5800237123914, 
    16.3660540610195, 16.2943338959264, 16.2882838904092, 16.1149610431176, 
    15.9902532934782, 16.1771430913517, 15.9718774351811, 15.449413709711, 
    14.7598398288204, 14.358105034194, 13.5382632648553, 13.2684174072685, 
    13.2548388338707, 13.0122888178767, 12.9582542337086, 13.1078714748098, 
    13.0709644113546, 12.8813409426255, 12.5911777120734, 12.5969920128782, 
    12.1882469589577, 11.8487505704945, 11.7268516386741, 11.5747050868159, 
    16.5350257049102, 16.2423361148076, 16.1010185010852, 16.0216630001076, 
    15.6924178794936, 15.4325643923803, 14.8234919250671, 14.0942076353167, 
    13.648778703474, 13.7204510872563, 13.9159283298611, 13.5036224938753, 
    13.470005189741, 13.3501553884762, 13.0357728539241, 12.8473819820657, 
    12.9725432636094, 12.9924146711808, 12.6636128173205, 12.5484714010504, 
    12.5531516092105, 12.2531349169049, 11.9637251308906, 11.9916121590243, 
    16.4781146943255, 16.2114191859008, 16.0737646116353, 15.6400276928673, 
    15.1842408151013, 14.823701027037, 14.0444487401235, 13.4586767299361, 
    13.4367700422436, 13.6452336371617, 13.6229296208032, 13.392648771423, 
    13.5395009395835, 13.3109172265273, 12.9665879473389, 12.8052181000056, 
    12.9489222336721, 12.7226056938746, 12.3238203438371, 12.3103498110002, 
    12.473581823615, 12.2639720794626, 16.2646511785483, 16.134951590965, 
    16.1715746611419, 15.3555320953927, 14.7707675023425, 14.3595790247207, 
    13.7871782289937, 13.4255840396576, 13.5265487532419, 13.6532080952398, 
    13.5350166870293, 13.510112142847, 13.2517494950487, 13.1403798700734, 
    12.8674607252126, 12.7183165630248, 12.7194087889134, 12.3066324796776, 
    12.1262814748031, 12.2731357772133, 12.2897692025666, 11.9770672104269, 
    15.9780587203902, 16.1515540484796, 16.2655418400614, 15.7699016125285, 
    14.9203304221776, 14.1344663955232, 13.6209695165014, 13.4205027003964, 
    13.5510756515082, 13.6366701846084, 13.4322958611519, 13.1397286023424, 
    13.1580169557819, 13.0042367499408, 12.789567484866, 12.6863113380505, 
    12.7301259003202, 12.2143565509648, 12.1237954267468, 12.111262731398, 
    15.9560361626836, 16.1495340355436, 16.1606896118949, 16.2119873972845, 
    15.435062038405, 14.3630278439039, 13.5735530883646, 13.5446077873605, 
    13.5965328191054, 13.602995292615, 13.5633278040603, 13.322986706391, 
    13.1618208844585, 12.9377443382565, 12.7401428477974, 12.7147061033367, 
    12.7041016280947, 12.5227984899658, 12.4730108523998, 15.9442651902805, 
    16.0842187046259, 15.9612514332229, 16.0239703565314, 15.7398195116788, 
    14.6852642483944, 13.7488254102796, 13.7729883288801, 13.7663501309659, 
    13.7465846306944, 13.8034610186571, 13.589701769748, 13.3351075999267, 
    13.1954407083997, 12.8491867284104, 12.6716783237036, 12.7250105027003, 
    15.6259784045221, 15.6308730718429, 15.6810859041092, 15.8396538206183, 
    16.181887764563, 15.2823729424805, 14.183387721029, 14.070672452121, 
    14.2701816387161, 14.260222552013, 14.0536993100342, 13.9065350261845, 
    13.7329952033599, 13.482523537154, 13.3024707877308, 12.8693905214471, 
    15.5991638149384, 15.4461717536741, 15.5122087103659, 15.627169992725, 
    16.0456935916401, 15.5991522615543, 14.6071857294877, 14.3667536799266, 
    14.6772767349785, 14.358250819993, 14.1845648932614, 14.0409158931746, 
    13.3278392962687, 13.2552952190112, 13.2542539475587, 15.5850662888356, 
    15.5769492057914, 15.6086446544522, 15.5257874978571, 15.9824292353515, 
    15.6437477591047, 14.852967216906, 14.6394804002835, 14.6379570641146, 
    13.9016095752282, 13.8264017379281, 13.6361842533275, 13.2550023866856, 
    13.1245983619084, 15.971012348325, 16.0024985711275, 15.7646493476715, 
    15.4191392815544, 15.8679159951815, 15.7312079969774, 15.0723032035443, 
    14.9121563405421, 14.3042981760056, 13.5887567049996, 13.3656452572882, 
    13.3048939929083, 16.190312293049, 16.278996408163, 15.7823487532561, 
    15.2820920180416, 15.6175251378555, 15.7266593570526, 15.1050370774673, 
    14.6903675296176, 14.05161091204, 13.5913139188284, 13.4511895285182, 
    13.360969771276, 16.2088893526181, 16.1779175881647, 15.6079327704288, 
    15.2732455543901, 15.3404681137098, 15.3454203534552, 14.8339358103639, 
    14.3851198728245, 14.0575689258695, 13.5731391612218, 13.5550507456194, 
    13.6336945723176, 16.35247393507, 15.9227050710971, 15.5003944181448, 
    15.62549465892, 15.4022700608063, 14.8632727865953, 14.5965456898623, 
    14.3110503175352, 14.2578385214299, 13.8730597526968, 13.5941107308173, 
    16.2592249284006, 15.6809720346324, 15.48735293877, 15.8234807276725, 
    15.640389520624, 14.8010514068461, 14.4641142939453, 14.4165465658774, 
    14.4572193426374, 14.0680597219141, 13.6853017127815, 15.7626984304509, 
    15.3757322214921, 15.5111061079146, 15.5332821543447, 15.1884436400797, 
    14.7501297248004, 14.3959592876676, 14.3060660341928, 14.1845518253422, 
    13.8493486229493, 13.5963403283514, 15.3738651526621, 15.1553568888779, 
    15.0276338820324, 14.8395809373933, 14.8033389016791, 14.627865266512, 
    14.5128143621712, 14.2226799149438, 14.1114841544519, 14.0415748230219, 
    15.4612303258942, 15.2928485361249, 15.2172966782025, 14.9705021957922, 
    14.6705766734428, 14.6693362233978, 14.619360680534, 14.4567029969371, 
    14.3008437187928, 15.8022175429719, 15.4809043848858, 15.42742427073, 
    15.0959956008342, 14.7406084721735, 14.4607082095522, 14.3892131130541, 
    14.5201940839027, 14.4485321791731, 16.087745412679, 15.6946908186666, 
    15.5852359952192, 15.4868344154039, 15.0946696355371, 14.6277019274825, 
    14.2049290308372, 14.295255279753, 15.9913297143777, 15.7514589226655, 
    15.4941907412007, 15.28312841489, 15.1069309883809, 15.876875916954, 
    15.4763849062793, 14.8845904782086, 14.8612403216798, 13.2836325389309, 
    13.2901696041177, 13.3215494874029, 13.30596106506, 12.994739602689, 
    12.4842339734821, 11.4932839523579, 10.2457535620789, 9.24982936326835, 
    8.43458162047381, 7.65351006569355, 7.02390906784671, 6.56315604641417, 
    6.1594969258866, 5.77633661863945, 5.45933606792874, 5.27138275669757, 
    5.09504003530588, 4.84209224835656, 4.60924102915853, 4.47008955838973, 
    4.33654547057626, 4.21130429761282, 33.1215360692035, 33.1207717751379, 
    33.1174912802448, 33.1230645148815, 33.1715763098267, 33.2482187944529, 
    33.408596853075, 33.6345163099807, 33.8132887446419, 33.9439481136966, 
    34.0557708210852, 34.1332498478489, 34.1829282938006, 34.227573065371, 
    34.2710825797059, 34.3045129335687, 34.3226561834867, 34.3384684345782, 
    34.3586102370292, 34.376997615444, 34.3884485312239, 34.3993958899198, 
    34.4092633699398, 11.9295135107994, 11.9678538491498, 11.990385878787, 
    11.945788042957, 11.8201855336721, 11.3619527601337, 9.84675904383059, 
    8.13720490089891, 7.39656494329402, 6.66787655756908, 5.99822862506876, 
    5.22970122036829, 4.65183401700823, 4.21881603978893, 3.78722375696716, 
    3.40060992903172, 3.07050439590039, 2.7810962003688, 2.53296927580216, 
    2.3142607961581, 2.15575651399982, 2.02170518539028, 1.92960794933378, 
    32.6499905004991, 32.6539612658927, 32.6554412465048, 32.6560295229312, 
    32.6599913867961, 32.6872481973336, 32.8841745894358, 33.320635562012, 
    33.6726325907358, 33.9228090112393, 33.980000107366, 34.0275302295351, 
    34.1240201392671, 34.2103250106915, 34.2990759046811, 34.3749223745146, 
    34.4317742185738, 34.4768683646941, 34.5119441214494, 34.5423404050731, 
    34.564207205878, 34.5822245972792, 34.5940770854183, 7.60407645282423, 
    6.34456694680316, 5.71132460381734, 9.72621088046892, 9.79939899317099, 
    9.84960750438525, 9.973292284575, 10.0649717192094, 9.93701052402682, 
    9.35570926096186, 8.46225691953717, 6.89983162312238, 5.96860108107276, 
    5.55211542951472, 5.44590702016772, 5.39831469901514, 17.5490322020655, 
    17.3507551413782, 17.1360909162866, 16.9244857757166, 17.1887216685931, 
    16.9001959578325, 16.6502667343571, 16.2954057753179, 16.2255275143984, 
    16.2662221845228, 16.2225809680072, 16.1519128177169, 15.9808608627598, 
    15.6324031576102, 14.7215687733068, 14.6739517312914, 14.5212745831834, 
    14.5119338624951, 14.2058702519688, 13.5511400220063, 12.9835272864452, 
    13.3399911508008, 13.1629188304434, 13.0064108945973, 12.9884062980349, 
    13.133535603073, 13.4390619098344, 13.2885966949351, 12.8759207296761, 
    12.356043397328, 12.5749267466045, 12.9502823691547, 12.5261780325159, 
    11.31714943162, 11.0440379098699, 11.0271619864136, 10.7299734832891, 
    10.7706332165784, 10.9123212838211, 10.9720095713715, 10.7085485326249, 
    10.5852566076638, 10.4012408171596, 10.2354382397903, 10.1373704625117, 
    9.91750770948347, 9.88692603992288, 9.65216975508518, 9.55930732044088, 
    9.44838048315776, 9.03768229075341, 17.5176983304324, 17.459133855379, 
    17.2029045608203, 17.1944634191382, 17.0146868603068, 16.9385853620817, 
    16.6682657838664, 16.2466779650999, 16.100771695927, 16.2785052734265, 
    16.1141551136866, 16.0738453525144, 15.9597092438591, 15.5894758252022, 
    14.7328070784581, 14.6376576939809, 14.4341652889906, 14.5564827722051, 
    14.4721082931936, 13.7549669982929, 13.2403483885716, 13.3379082281289, 
    13.3370500186314, 13.0117581456297, 13.077624524759, 13.3176216258604, 
    13.4869621764698, 12.7585319470501, 12.2499906290201, 12.3224819845046, 
    12.3980542746339, 12.3016561359865, 11.6767218198552, 11.1077203407971, 
    10.9914963012984, 10.9485608749866, 10.7368557583923, 10.7419085569105, 
    11.0081711395393, 10.8945432931019, 10.6594380754782, 10.553486883021, 
    10.3488258315424, 10.0180641591871, 9.86423728264649, 9.93226410494719, 
    9.8477782056348, 9.70846916826152, 9.51474066808639, 9.35830787832804, 
    9.15818145782087, 17.3613743092776, 17.3498287984136, 17.2479205143942, 
    16.8300025275618, 16.5683349232211, 16.5741270566818, 16.4943936857774, 
    16.1353894868762, 15.972509408608, 16.2064000351314, 15.9975650491797, 
    16.1278905017828, 15.9023088236696, 15.4196993805097, 14.8911486124132, 
    14.7879751946304, 14.8050149412837, 14.8349870881176, 14.2383003719828, 
    13.8388093135143, 13.5014573964041, 13.3354153754545, 13.4167925305712, 
    13.3161100420751, 13.3931236365387, 13.4487211549887, 13.0502991503717, 
    12.2670418769364, 11.995245410103, 12.0187584447882, 12.0134928279434, 
    11.7760790558463, 11.3745511796378, 11.2868844436289, 11.0182640799796, 
    10.8646779678978, 10.733778114205, 10.7846229201404, 11.1523357707912, 
    10.5138637331053, 10.2610777240825, 10.3166817231743, 10.0336881576455, 
    9.57854767046189, 9.50685944369389, 9.76059630001698, 9.69163647756828, 
    9.7479782583968, 9.51161095873406, 9.27260370614223, 9.04937368134152, 
    17.327895715746, 17.1730646973719, 16.9870152566317, 16.505547268657, 
    16.3786730966926, 16.1796483582032, 16.1553381305447, 16.0448369844835, 
    15.9911898658802, 16.1258987110498, 15.8228343126503, 16.0148554938878, 
    15.8592197341239, 15.4212934176434, 15.1240049777028, 14.9201165116635, 
    14.9843005731977, 14.4895490009761, 13.8860398082076, 13.8281687455386, 
    13.4862830642639, 13.3749182276517, 13.4327857294088, 13.552033104959, 
    13.3951918660681, 13.3916748918142, 12.9260635934374, 12.1036470850887, 
    11.7816844911011, 11.6566208702918, 11.7816570062026, 11.576474919627, 
    11.331385944092, 11.2803929090949, 11.1200991886111, 10.9144900684141, 
    10.8425232649452, 11.1375693958523, 11.2555110542213, 10.281653139505, 
    10.0523604169584, 10.1854340032555, 9.67272877850269, 9.13851755339341, 
    9.23951721518599, 9.26364734820769, 9.3428597059045, 9.36181055795382, 
    9.51941495692226, 9.00344957249223, 8.79998879788096, 17.3839415445673, 
    17.2443621101345, 16.8789161522721, 16.6455800881745, 16.5767385679366, 
    16.1406764301486, 16.0951978037995, 15.9793841809442, 15.8940925039569, 
    15.7389140418428, 15.6920177747859, 15.9591277963924, 15.8504214009318, 
    15.5083356950343, 15.3449461570343, 15.0075602021721, 14.8511742886303, 
    13.5640528079474, 12.9616573170152, 13.0782457780088, 13.0166046538155, 
    13.1352366324077, 13.210728349569, 13.4894038502995, 13.5472812726151, 
    13.1836095850666, 12.7591548439909, 11.649138312037, 11.1516698368223, 
    11.2470967628457, 11.6874792838783, 11.5934136961892, 11.1868616698435, 
    11.1270889308022, 10.9651204353901, 10.8513818102436, 11.0068701600275, 
    11.1372960876882, 11.238549642109, 10.2486519973695, 9.88435593441409, 
    9.81323374128168, 9.48858618706461, 9.1923772236199, 9.38111918891549, 
    9.26949053498607, 9.33209295488255, 9.41504529733739, 9.27958919286109, 
    8.90632539756079, 8.77322101687147, 17.4808465737447, 17.3018669444747, 
    17.0245585521542, 16.8370513358249, 16.84424195285, 16.1843537847434, 
    15.9177626995472, 15.8986604391268, 15.7478991601732, 15.4952227608794, 
    15.6510450904465, 15.764677470677, 15.8739732386621, 15.6587628945643, 
    15.4057323265632, 15.0848131798555, 14.5291557734461, 13.1711711267928, 
    12.6611498149061, 12.8584381045825, 13.0004426144501, 13.2768118622272, 
    13.2673714392634, 13.4536223869643, 13.4960520333349, 13.0291910640811, 
    12.4933134154189, 11.3353217878986, 10.963367558731, 11.0155311884123, 
    11.3019031175554, 11.3063753607024, 10.861795515486, 10.6026627675831, 
    10.4437928414009, 10.4240358048819, 10.5772550435908, 10.7715410157126, 
    11.0839647942043, 10.2640430076646, 9.89656658309147, 9.64796791523904, 
    9.45286086188571, 9.39022998341614, 9.57215613812367, 9.33898352006154, 
    9.32789823602002, 9.41475248505545, 9.2338055663562, 9.01516366118783, 
    8.76086538358596, 17.5493871774134, 17.3409438412061, 17.0694869526527, 
    16.8180882336991, 16.8393572998883, 16.1808550555182, 15.9100853432851, 
    15.879955123997, 15.6074431950819, 15.4828677526517, 15.5282593401408, 
    15.6032940409137, 15.6400010396876, 15.3583981930635, 14.736973897299, 
    14.278550632321, 13.8021667395684, 12.8075283322452, 12.6238174116171, 
    12.7059641084048, 12.9589806335234, 13.220528630906, 13.2254702747881, 
    13.3797931091236, 13.337926047807, 12.6554883713294, 11.923158868127, 
    10.9070465531008, 11.2334588794533, 11.0740703876992, 11.1024852301288, 
    10.9639289222911, 10.7819267438708, 10.4613320815232, 10.3530190033825, 
    10.4917148613592, 10.6039986361297, 10.6347583424777, 10.9641154055372, 
    10.4101549664972, 10.1438004106878, 9.72162528782854, 9.49699706953168, 
    9.40003384627918, 9.66829211458778, 9.50848856132438, 9.25214891171136, 
    9.32864704391921, 9.24798091856441, 9.25405577684088, 9.08979333730313, 
    17.4497672771657, 17.4293895688247, 17.0784167061714, 17.0819738308607, 
    16.7767184726513, 16.2994167583538, 15.9413277214214, 15.868852233424, 
    15.5958336472159, 15.410310131615, 15.2806562848509, 15.312767022726, 
    15.4306211237578, 15.2316420069215, 14.4238938895957, 13.548425822004, 
    13.101266009385, 12.5440323310685, 12.5360879120446, 12.8003915201849, 
    13.1024334957308, 13.2697130607676, 13.3016345861764, 13.4270958958512, 
    13.0016070665037, 12.1434790512946, 11.4937511208027, 11.1559103233396, 
    11.3279298737731, 11.3244146644764, 11.2623628050238, 11.0291402843458, 
    10.8265780595674, 10.3825698910486, 10.3805377398021, 10.4365620142374, 
    10.6110452695211, 10.7697310445002, 10.9481805840123, 10.6448745148822, 
    10.3871829261588, 10.0711270474642, 9.67060810911934, 9.54944396442651, 
    9.70016541091929, 9.70050676559066, 9.300200551675, 9.2813172073337, 
    9.25506503114516, 9.16152801229596, 9.15586285595143, 17.5328332619739, 
    17.3711112333525, 17.324074705589, 17.1447888834113, 16.8886102406835, 
    16.3653731103719, 16.1476795560047, 16.0194936476571, 15.6389150308638, 
    15.1116322358948, 14.6358376864279, 14.4394147624836, 14.6683265135502, 
    14.9847493705931, 14.6739502012817, 13.9161004003461, 13.0325648525082, 
    12.5948601052053, 12.5309911579408, 12.8534805530092, 13.2541623016923, 
    13.3975301258779, 13.4595964823806, 13.5096670507321, 12.8034768124259, 
    11.8452377289877, 11.2976452936069, 11.2261887654593, 11.4316246990678, 
    11.3716504951068, 11.3139251661385, 11.1680003041985, 11.0619829779332, 
    10.6375885459018, 10.5705616458544, 10.4123971422072, 10.4932407987831, 
    10.6723237294618, 10.9736063593204, 10.8286421364934, 10.5505545319459, 
    9.90280759526977, 9.73991646208232, 9.74412258005025, 9.71861664409989, 
    9.73602807702805, 9.42925012971559, 9.28199333033379, 9.19598801675317, 
    9.11037385863609, 9.22014470358827, 17.2743849358438, 17.4261790142341, 
    17.4350217215478, 17.3445355721611, 17.1043415553599, 16.6078328934327, 
    16.1754139838537, 15.834649049171, 15.4951199897457, 14.7437765422024, 
    14.0078953725726, 13.7156114828462, 13.8438067176725, 14.1033257807733, 
    14.2798437457421, 13.6736533111852, 12.8500381174297, 12.592939439508, 
    12.5264337915624, 12.8551843255927, 13.2384073113753, 13.4359692832766, 
    13.4593006703559, 13.3626360935491, 12.6080172712442, 11.6952403003462, 
    11.206754487778, 11.1915652806293, 11.6356463879125, 11.4762903437551, 
    11.2509757251941, 11.2643476275002, 11.1653375656143, 10.8854041462105, 
    10.8127616009048, 10.3959537467141, 10.5702681918331, 10.5734480061288, 
    10.39445047306, 10.5928380626902, 10.3015532222901, 10.1104592722025, 
    9.97585903594167, 9.91896559903513, 9.84215027449995, 9.71945588434273, 
    9.55425800790278, 9.26660328661773, 9.27348396394248, 9.1157596378807, 
    9.09589238059243, 17.1381563536538, 17.1666058501138, 17.2269006224409, 
    17.2899941679911, 17.1223128689338, 16.9278992664661, 16.4091149085218, 
    16.0560237502362, 15.4659136934534, 14.7795761072649, 14.1588282402015, 
    13.7981132181606, 13.6869485220007, 13.6116737318509, 13.5359113226241, 
    13.138524092838, 12.6605330142561, 12.5926980607463, 12.4832025583476, 
    12.7751525941771, 13.0798767892038, 12.9618204553882, 12.9703572311179, 
    12.8879133246474, 12.4721115024183, 11.7203571203575, 11.217900094222, 
    11.2942636827725, 11.7414584751486, 11.5384584063638, 11.0963071876201, 
    10.9233169496445, 10.7711725693361, 10.7052838107271, 10.453735747966, 
    10.1788398033487, 10.6671867591862, 10.7041463387703, 10.5274996717237, 
    10.3295876967389, 10.0551347378684, 10.0094861104803, 9.77887794017243, 
    9.63046427983172, 9.59979379316735, 9.3338277680332, 9.48365279785212, 
    9.20562426371077, 9.29082168732747, 9.21945252955002, 9.11705030837643, 
    16.9857335308942, 17.1776214260883, 17.1811813077971, 17.1996316842552, 
    17.349948459891, 17.072573494361, 16.6351133122843, 16.1374351787131, 
    15.3678247046435, 14.7061625312062, 14.3065525325548, 14.0027150175437, 
    13.9145977771993, 13.8669239532722, 13.5446438185907, 12.9514809872724, 
    12.568521005806, 12.6401233554096, 12.3634611471124, 12.5408912410125, 
    12.8671952411135, 12.8838359664007, 12.7680541722814, 12.6031052109591, 
    12.3213252641381, 11.8595864991142, 11.4353560591028, 11.4180373534386, 
    11.6959698028821, 11.4395636525395, 11.1160017039642, 11.0534682780208, 
    10.6000757641463, 10.3270750149498, 10.2359863116476, 10.3200385454406, 
    10.6585805610993, 10.676039088139, 10.4710847237615, 10.1898328418737, 
    10.057919722444, 9.93477522292179, 9.61069709118961, 9.44468308176244, 
    9.47760698334842, 9.36952007807336, 9.34236009581103, 9.19803428385436, 
    9.39059223890028, 9.25583816452855, 9.1487153206635, 16.8400884056555, 
    17.026203077381, 16.9889073704613, 17.0614654418857, 17.301675115735, 
    17.2094855086068, 16.5563049415428, 15.9488247332286, 15.0585413553909, 
    14.4125621488271, 14.2191884491406, 14.0445372600694, 13.898613492709, 
    13.8820932995685, 13.7029691845711, 13.175381827029, 12.7936515271168, 
    12.7665199878048, 12.2367340752481, 12.0797998490726, 12.3270024494383, 
    12.6612400228724, 12.7369895855782, 12.4689956882433, 12.1125710980299, 
    11.8313098698425, 11.3309387203504, 11.5095037549305, 11.6281375689807, 
    11.2127409281222, 11.1942416243109, 11.1999530866311, 11.2328125098283, 
    10.726890869957, 10.8859051814495, 10.8525286208333, 10.7183190334851, 
    10.7237484821143, 10.5361223468619, 10.2794970684767, 10.1551949564321, 
    9.94161135749807, 9.79396543140974, 9.68211119296794, 9.62918229784668, 
    9.50175694100289, 9.58164192251262, 9.42921916100224, 9.48650878810354, 
    9.33165634662977, 9.19071975202753, 16.612249154619, 16.7493322645505, 
    16.7121820525367, 16.8510215484592, 17.1395177100583, 16.7856482208939, 
    16.3428269275098, 15.6706299814578, 14.8338756943886, 14.3321871835371, 
    14.1940843652164, 14.186667283915, 13.9173233898348, 13.8547309552855, 
    13.7577434723876, 13.3681663975001, 12.9895281359479, 12.9163586698942, 
    12.3669702328126, 11.8647992104586, 11.8972440316823, 12.3759081502193, 
    12.9319788582799, 12.5394769407534, 12.1235206357112, 11.6929899683882, 
    11.8144445493201, 11.4820633681562, 11.3399554588705, 11.0974096656235, 
    11.182878857183, 11.3617365138547, 11.20915728097, 11.1971038904474, 
    11.1741020366053, 10.7755045167593, 10.5253767350114, 10.617551914662, 
    10.489258227573, 10.3155290698972, 10.0944262711757, 9.84682349959375, 
    9.80733957250043, 9.63826501916716, 9.46311799818488, 9.42487669324252, 
    9.52776247277889, 9.4783909260198, 9.41045710217451, 9.2696662126647, 
    16.32332973892, 16.2216120534903, 16.1389367874931, 16.3677151141521, 
    16.7000605617049, 16.8406107491586, 16.3990742190193, 15.6315709920507, 
    15.0038619047806, 14.8569183974607, 14.5970180373097, 14.2805317399147, 
    13.834109834049, 13.7741009507984, 13.9258697253556, 13.3539794428197, 
    12.9938187696521, 12.8625380528104, 12.3211849490723, 12.1584847233763, 
    12.0087177814937, 12.074624265971, 12.5853318062377, 12.366114619444, 
    11.9844860798507, 11.6929817220801, 11.7210574528781, 11.1605995959339, 
    11.3035954689638, 11.1628064684879, 11.1995619581693, 11.2717100083575, 
    11.0095478661391, 11.0964751623535, 10.8182393955784, 10.584778325157, 
    10.4152510625546, 10.4944095992078, 10.5437993662132, 10.4878586967414, 
    10.3088191016522, 10.1407159172167, 9.75744353418658, 9.6482716818535, 
    9.57137779465879, 9.43952738237303, 9.4049507612829, 9.4922678769349, 
    9.48842713629767, 16.2203918820307, 16.0164567626291, 15.927689902608, 
    16.0343659541599, 16.2534746817701, 16.4790639845745, 16.3647849039423, 
    15.8772594140698, 15.3842419799632, 15.3495434206044, 15.2596662863533, 
    14.4671905675399, 13.7003228172479, 13.6063113389169, 13.7194409171556, 
    13.1640564097315, 12.8451357845701, 12.6218641064046, 12.3998659496399, 
    12.5741118845189, 12.2733889097674, 11.8600388996777, 11.9976549071754, 
    12.3479268061016, 12.2799148593646, 11.8061959548285, 11.4095461863417, 
    11.0761324986525, 11.1272560011061, 11.2135674481589, 11.0734023226178, 
    11.0905845264905, 10.7623465940239, 10.9199587129867, 10.5041629526432, 
    10.4560549150593, 10.524374765281, 10.583037265942, 10.5179402293148, 
    10.3196905737662, 10.2211125883589, 10.1295708618833, 9.97885713851631, 
    9.76723516715058, 9.62089277113365, 9.82517553869975, 9.56994536302467, 
    9.52761579280329, 9.54172980373307, 9.48766540538324, 9.47125869430659, 
    15.9613607971049, 15.9706709490602, 15.8878435959784, 15.7911347479971, 
    15.9032494668314, 16.1675732676556, 16.3573163957752, 16.1244498500605, 
    15.7690757862166, 15.6892633595289, 15.6952742769087, 14.6446745428555, 
    13.3916017189703, 13.5203670504568, 13.5184988232885, 13.0908188088625, 
    12.7994100225633, 12.5810933861615, 12.6316545306421, 12.7826877348197, 
    12.5038629658613, 12.0582761021887, 11.7336161927381, 11.7465851520307, 
    12.0471253601804, 11.8684858155635, 11.475432733824, 11.26686824799, 
    11.2274528566192, 11.1855572432104, 11.0132274860627, 10.8022900851119, 
    10.7048678923519, 10.5951932714674, 10.5768507089576, 10.1894360320893, 
    10.3438478057551, 10.1842859249663, 10.0484825633455, 9.85825036963935, 
    9.83586188985253, 9.74281006499271, 9.55792489429517, 9.44564862012365, 
    9.36775534153666, 9.20039995079635, 8.8585132730361, 16.1539146402506, 
    16.3527151258779, 16.1872476199933, 16.00395972769, 15.8921930731193, 
    15.9037591167497, 16.1297327176817, 16.2673192672669, 16.0899668235647, 
    15.9542775157351, 15.3425482461932, 14.0277591232294, 13.1824397830089, 
    13.263786430963, 13.34363757897, 13.1470227943452, 12.9390518150067, 
    12.7341734575706, 12.7814721285606, 12.8800249502787, 12.5542664648894, 
    12.1425437277097, 11.7698100410952, 11.800691476329, 12.0410120715475, 
    11.7981822247082, 11.4706715907027, 11.5176810506531, 11.3755108785156, 
    10.9849605872868, 10.7951488803801, 10.6843140481753, 10.4359370638537, 
    9.8063527404827, 9.67873737027077, 9.75291301383588, 9.50440209298553, 
    9.25694013572357, 9.19322992078024, 8.76515073294782, 8.46758771981115, 
    8.35749139331784, 16.4267124522081, 16.3153200641896, 16.2883811710048, 
    16.2805970442435, 16.1248556328549, 16.0418729647479, 16.2420126954609, 
    16.3635174876074, 16.3400264661852, 15.8154089116163, 14.7250069517969, 
    13.5775327393213, 13.0651786656349, 13.0703648019761, 13.0431490178017, 
    13.1268003061611, 13.0204604153611, 12.9950052461642, 12.8714296842572, 
    12.6936326133942, 12.4918106110485, 12.1328131654186, 11.5924758225757, 
    11.6333091661222, 11.8021496562087, 11.8515049796992, 11.8454825588967, 
    11.7632792562096, 9.61430952181943, 9.33319174468243, 8.98697531779376, 
    8.25081637535274, 16.4679209634108, 16.2702594313268, 16.1689364859538, 
    16.1847258224493, 16.0848054789095, 15.9329191944069, 16.0942779130216, 
    15.8057036500095, 15.271078330942, 14.6487415502256, 14.2873540720363, 
    13.4127225908675, 13.1629061997223, 13.1680884873542, 12.9088787704282, 
    12.8744884789779, 12.9989843731583, 12.97914744271, 12.7419114960986, 
    12.4793906377062, 12.499184444166, 12.0696245554473, 11.7258792010378, 
    11.6523257149134, 11.4685844205253, 16.4530049950393, 16.1675228080952, 
    15.9866077669525, 15.8712044152071, 15.6041681058237, 15.3406480369671, 
    14.6641728453412, 13.9150878061747, 13.5085208702132, 13.6669487858747, 
    13.8506790759685, 13.3749421338527, 13.3574143478191, 13.2513844990026, 
    12.9833293656989, 12.7328324926957, 12.8741096694419, 12.9018738753194, 
    12.5933859155373, 12.4421461900026, 12.4448283285342, 12.1428238247855, 
    11.8147163495409, 11.8364946327874, 16.3794533963629, 16.1019457016285, 
    15.9493771624097, 15.4721928572983, 15.1204713446552, 14.7848456240907, 
    13.9012319700748, 13.3104680532297, 13.4069645355488, 13.5535794097968, 
    13.5366698995293, 13.2838045213518, 13.4304718143138, 13.2038219581513, 
    12.8352458572489, 12.6851032704873, 12.8070568881281, 12.5397892687496, 
    12.2167720291063, 12.1986607834161, 12.3979974917601, 12.1318960531285, 
    16.1815096768713, 16.0328171178739, 16.0384810997717, 15.1671865632494, 
    14.7023864123715, 14.3737257946487, 13.6696265213194, 13.2941243555355, 
    13.4581855871944, 13.5077389247327, 13.383832496344, 13.3692612866025, 
    13.148785910915, 13.0387043586163, 12.7819154165577, 12.6148814154876, 
    12.568186377805, 12.1176840726799, 12.0781378266383, 12.2241941760565, 
    12.1396497579465, 11.9189142889895, 15.9110201999802, 16.053095402702, 
    16.1683868218368, 15.627499334663, 14.7555902425648, 14.0434700820242, 
    13.5571449065459, 13.3218376856742, 13.4710064531285, 13.479886646897, 
    13.2905653890925, 13.0671608244993, 13.0827930947195, 12.8877138251484, 
    12.7068921260375, 12.6235672172183, 12.6565603188862, 12.1488567286269, 
    12.0850032091214, 12.1026143775967, 15.8940766509, 16.0625764310118, 
    16.0668991849133, 16.0967493318646, 15.3200048220498, 14.2076022461133, 
    13.4866641806137, 13.413133181069, 13.5075658784996, 13.5295497579957, 
    13.4813004000539, 13.2312812337439, 13.0643986458959, 12.8793890653428, 
    12.6848717819618, 12.6453700302789, 12.6128004711151, 12.39434287499, 
    12.4542608340335, 15.8453934742671, 15.9204275606256, 15.8194028255652, 
    15.8677811000906, 15.6039249321512, 14.4651145912515, 13.5638929170585, 
    13.6450604358996, 13.7104945795841, 13.7660291680082, 13.7429810274646, 
    13.4920562247435, 13.3268673342315, 13.1800516927819, 12.9166802319093, 
    12.6711986946131, 12.6527614933002, 15.4979979007076, 15.4594054798035, 
    15.5309789968229, 15.6961033945838, 16.0335678857195, 15.0885266385303, 
    13.9941877816387, 13.9235113151349, 14.1690296241839, 14.2256909837026, 
    14.0298487747548, 13.8766444475096, 13.6732058428012, 13.4429946267294, 
    13.2957075407187, 12.918242322289, 15.4024405306156, 15.339613788924, 
    15.4032511521105, 15.4974189646575, 15.980985335374, 15.4917205804088, 
    14.4849201469923, 14.242208858257, 14.5294361414449, 14.2868139205181, 
    14.0555625178299, 13.9185185499825, 13.2654098936906, 13.0852535010316, 
    13.0492614759158, 15.4660230543657, 15.5757899860936, 15.516913994844, 
    15.3725662319956, 15.8670103953443, 15.5704775013414, 14.7412647311254, 
    14.5554133816057, 14.4941062342211, 13.7977148206428, 13.6882732654371, 
    13.510617852493, 13.2022066091896, 13.012851617162, 15.8430844698062, 
    15.9699359504236, 15.6351153939313, 15.2864757634796, 15.7063819943123, 
    15.6082301455632, 14.9190931194913, 14.7805187503105, 14.1886514576158, 
    13.5096311099946, 13.3029802731349, 13.2236583583768, 16.0453343812429, 
    16.1604535132066, 15.6314714032731, 15.2047791169296, 15.4965114807538, 
    15.6157580454681, 14.9798190772216, 14.6528988755158, 13.9877423916154, 
    13.5416740924837, 13.3828587499907, 13.3856968277813, 16.0748166371427, 
    16.0030270022034, 15.463804933301, 15.2315473104189, 15.2488662238947, 
    15.3152669854475, 14.7624742602246, 14.3283116789128, 13.9619689315327, 
    13.5224275153695, 13.4988583228666, 13.5704520655965, 16.1963082074558, 
    15.7719962030696, 15.4024356410963, 15.5466563148506, 15.2236669537251, 
    14.792458201199, 14.5415828902196, 14.1923966559067, 14.1517335310029, 
    13.8413505755326, 13.5563922493618, 16.1411201898127, 15.5253569705719, 
    15.401342260936, 15.6710453116296, 15.4118159055664, 14.6379708284275, 
    14.3854964292816, 14.2756266269506, 14.3209117903392, 14.0207474047721, 
    13.6105107076626, 15.681846619912, 15.2523324758372, 15.3936010663005, 
    15.2510297325078, 14.9253875964453, 14.5816981351332, 14.2684303458067, 
    14.1434772777564, 14.0680139521165, 13.7836759323592, 13.5128425535823, 
    15.1888874356576, 15.0212090072762, 14.8937262420137, 14.7247469508163, 
    14.6534184457273, 14.5198392014269, 14.3271063754292, 14.0785839344894, 
    14.0629185292784, 13.9319607135005, 15.2857931986359, 15.182647216601, 
    15.1192257047361, 14.8617406376699, 14.5593432134379, 14.5425771056438, 
    14.4549263742102, 14.3259732503281, 14.2012982008974, 15.6610145547105, 
    15.4060501958714, 15.3643828817965, 15.1037487799041, 14.6977975988449, 
    14.3375320248121, 14.2884641303968, 14.4308415264418, 14.3263284883853, 
    16.0217398893713, 15.6738558802456, 15.4997261254889, 15.3776831083407, 
    15.0228063650608, 14.5259758897015, 14.108427449233, 14.1555001268177, 
    15.9120296012236, 15.651326056417, 15.3832917814109, 15.1408634178136, 
    15.0282980581986, 15.7580074873842, 15.4175774251711, 14.8209331833149, 
    14.7764022231345, 11.0459841734491, 10.7076628358506, 10.7141592390182, 
    10.7723059786126, 10.9776256870242, 11.0904761769335, 10.7048953991086, 
    9.78748340559323, 7.65751928421421, 6.76625560899773, 8.55356608029929, 
    7.09116153649079, 6.64897401779203, 8.97971031862114, 7.25615039669867, 
    6.62319130007796, 10.0961535158784, 7.98739536697413, 6.85028030835674, 
    6.51681598805875, 10.7133466745783, 10.7205168155948, 10.7697097596984, 
    10.9394560863547, 11.1641917167978, 10.8120807003867, 11.2347817984174, 
    14.2377032482042, 14.2755557001339, 14.2903273451039, 14.3217649942396, 
    14.3698033220677, 14.2513196974295, 13.8039936937349, 33.2864275689248, 
    33.2855133035496, 33.2848605013345, 33.2835647556008, 33.277207100172, 
    33.268272123986, 33.2549923718528, 14.2254019234868, 14.3056559791272, 
    14.3526303146085, 14.3887127051948, 14.3610032028539, 14.1473543128256, 
    13.5321127941588, 12.208258504056, 11.18584692061, 33.2658993207596, 
    33.2649289978701, 33.2641881179336, 33.2626392621178, 33.2606660702438, 
    33.2617122908558, 33.2673290213542, 33.2774488792579, 33.4065846733657, 
    17.4940237447818, 17.3082313065499, 17.1357573982407, 16.8956639551141, 
    17.166269037614, 16.9200098723995, 16.668026613412, 16.3204215312297, 
    16.2482985354732, 16.2821842369384, 16.2693608168309, 16.2001103904527, 
    16.1010776846324, 15.7092990111831, 14.7589976588341, 14.6865703288808, 
    14.5538654816157, 14.5341038037486, 14.037256101707, 13.4748014400316, 
    12.9730447195392, 13.3636379013785, 13.1716420767543, 12.9985591344996, 
    12.9405182910085, 13.0458714931799, 13.3604361622301, 13.2440901866965, 
    13.0061407816432, 12.434896949674, 12.7096689107808, 13.0977814029436, 
    12.6747883052295, 11.406143641844, 11.1303718945708, 11.0625693032701, 
    10.7909964870795, 10.8071982793825, 10.9402594567088, 11.0148977006467, 
    10.718880180573, 10.6283117110601, 10.4418942089774, 10.3105932581876, 
    10.1988065598801, 9.94044378579039, 9.93750569425623, 9.71052259486606, 
    9.59179616963373, 9.49025662502172, 9.1463273648331, 17.4657707862277, 
    17.3746722983196, 17.1473012619192, 17.1385043559371, 16.9980319449229, 
    17.0104030721074, 16.6983777325159, 16.2957782331128, 16.1336461207491, 
    16.3329545477491, 16.1211629451789, 16.1209342986075, 16.0800977720057, 
    15.7432571188652, 14.8029843067991, 14.647394399596, 14.4669296435412, 
    14.5781325115958, 14.4920725176373, 13.7295630986199, 13.1760184754165, 
    13.385995126529, 13.4389153376344, 13.0971050650792, 13.0285236110151, 
    13.283171289235, 13.4942413957451, 12.764944303075, 12.357241612943, 
    12.4006528666343, 12.5041850103387, 12.4629512395241, 11.8257434540391, 
    11.1256032877321, 11.0403699897865, 11.0320829073544, 10.8036024752937, 
    10.7705672094561, 10.9896870492255, 10.9507109801432, 10.7291454166935, 
    10.626329205186, 10.4248119303652, 10.1347257570694, 9.95140919751491, 
    9.96286707190987, 9.87363948851514, 9.72031421041698, 9.54936811632527, 
    9.41748590827225, 9.19187614872339, 17.3048817957646, 17.3127867741792, 
    17.1775839259726, 16.8101517862855, 16.5533461636789, 16.6125010021914, 
    16.5245586034667, 16.1937091749471, 16.0342485880013, 16.2641567670517, 
    16.0416231174047, 16.1776688056061, 15.9757840730158, 15.5861407060302, 
    14.8869909159228, 14.8149324933222, 14.7764007549532, 14.836685193364, 
    14.3375983927366, 13.8484769844738, 13.4883388548675, 13.3970075767277, 
    13.4643860696842, 13.3412811558371, 13.4134730615102, 13.4617021386096, 
    13.0430082357394, 12.2603045511497, 12.041052118764, 12.1141609721812, 
    12.0748358377492, 11.8209860701556, 11.3856893881317, 11.3004834848433, 
    11.0326545515325, 10.9552560906688, 10.7868538187229, 10.7590178421734, 
    11.0984703095706, 10.5866218532505, 10.295073716876, 10.3730620071782, 
    10.1696394420691, 9.72662237223484, 9.5723942900886, 9.83644719240189, 
    9.74896355695564, 9.75920252558592, 9.50488269721675, 9.26043394961534, 
    9.09796908228406, 17.2546896988696, 17.1302411789328, 16.9316841106649, 
    16.4822573651984, 16.3364535018478, 16.1794036688337, 16.1732183315982, 
    16.083158450128, 16.0693600130231, 16.1669355203839, 15.8726294655479, 
    16.0659493411229, 15.9063132576803, 15.4709015873665, 15.0732248793592, 
    14.9628546709614, 14.9431933674459, 14.4174455359256, 13.908269120374, 
    13.86796694758, 13.5904537580274, 13.4155349364975, 13.4584293131053, 
    13.5501806130731, 13.4687429140912, 13.3794322578749, 12.8228333256419, 
    12.0343570051821, 11.7624305444824, 11.6671931830657, 11.8097357936912, 
    11.5792982345119, 11.3981116436772, 11.2959363253739, 11.1046059452305, 
    10.925195080207, 10.8223331933456, 11.031192541443, 11.2385285481024, 
    10.3199283441472, 10.0725131022526, 10.2292317901672, 9.76329230275622, 
    9.21672537626942, 9.27444755041809, 9.32384321963105, 9.42029765473705, 
    9.40201254611006, 9.51133686030039, 9.02585294809042, 8.871303749005, 
    17.3644660130517, 17.1803335479513, 16.8303936529653, 16.5753806986534, 
    16.512415894703, 16.0996018558841, 16.0992165800432, 16.0183688947147, 
    15.924116005606, 15.7640965238709, 15.7456712745818, 16.0004083512787, 
    15.8737668153039, 15.4803608520618, 15.3429234235019, 15.0598693430472, 
    14.7587086783415, 13.5640764894809, 13.0405111399126, 13.1063027714218, 
    13.0558497060993, 13.1260510995989, 13.2090836258762, 13.5049949636455, 
    13.5692385140178, 13.2260565254604, 12.6884915316802, 11.6473050580687, 
    11.1820843366292, 11.2735313408862, 11.7151293219394, 11.626142841967, 
    11.2364655277289, 11.1176990764299, 10.9453369001792, 10.8437364293489, 
    11.0169301718818, 11.178376415845, 11.2702008977248, 10.2280818954962, 
    9.89621100790703, 9.91319484680761, 9.55778252465463, 9.21074162109023, 
    9.41849479992283, 9.29106361391808, 9.39069049503401, 9.41982253689183, 
    9.30356951276235, 8.81509281855824, 8.80071347591644, 17.4518130952085, 
    17.3432979541893, 16.986409921118, 16.8011356568218, 16.7667459270767, 
    16.1209044269016, 15.9172630482088, 15.8900920774844, 15.7459058407629, 
    15.5243845118224, 15.6772428531149, 15.7990761461217, 15.9058913014611, 
    15.6670035046582, 15.5313040221239, 15.265701077607, 14.6361101856454, 
    13.1967211636155, 12.664381738911, 12.781512507386, 12.9678806150424, 
    13.2517538633018, 13.2705042512506, 13.499593584011, 13.5584594538783, 
    13.11583208789, 12.5482459340397, 11.4308892012675, 11.1322420384249, 
    11.0337844935763, 11.3331192467537, 11.3967143459277, 10.9114147314063, 
    10.645723436463, 10.466038672811, 10.4399264414847, 10.6565513683398, 
    10.8438122109081, 11.1527823558936, 10.2453241748855, 9.87408732944989, 
    9.7007653553033, 9.49645280985696, 9.40132758990622, 9.58173831697806, 
    9.36682735314007, 9.35381171355861, 9.41921653937455, 9.18197600849663, 
    8.90464802196317, 8.70561945661348, 17.4558043604532, 17.377523764821, 
    17.0330693064121, 16.7549010193693, 16.7443530738744, 16.1008102496544, 
    15.9070575562723, 15.8384587105003, 15.5716049088994, 15.48065302544, 
    15.5188725219568, 15.6259210632244, 15.7038597077288, 15.4443813699183, 
    14.964861499803, 14.6651913165246, 14.1335927034744, 12.876566321194, 
    12.5984138689531, 12.6830611823082, 12.8894977353779, 13.1668479692404, 
    13.26268118032, 13.4498675772483, 13.4029858508331, 12.8188093061067, 
    12.0458594367142, 10.9823387509496, 11.2856706664559, 11.038552062971, 
    11.1334022550756, 11.0367867006963, 10.7589745518143, 10.4617630701104, 
    10.3857378210145, 10.5241274537062, 10.6289597038916, 10.6824045850439, 
    11.000164211682, 10.3828210491337, 10.1115670091633, 9.69167317663934, 
    9.49846812194178, 9.41940831714993, 9.63757970414679, 9.49244794409258, 
    9.25379404400176, 9.36756902535445, 9.20377517901775, 9.16963406543799, 
    8.95640023743502, 17.3634028690521, 17.3658246358887, 16.9787236940101, 
    17.0223814240003, 16.6976282426287, 16.2088431696177, 15.8685730675951, 
    15.8131554579118, 15.5537417985138, 15.3580517107704, 15.2329099329521, 
    15.3309192737962, 15.4627382892172, 15.1482046055186, 14.3695105883639, 
    13.7065754422805, 13.3708867859067, 12.6100485886776, 12.5396572264486, 
    12.7906617491001, 13.092796783476, 13.3204340905715, 13.3372116744598, 
    13.4661844129225, 13.0454419280075, 12.3101387405436, 11.5942711758469, 
    11.1947789561988, 11.3879757313267, 11.3208603726135, 11.3400711276434, 
    11.009918105024, 10.8182042411329, 10.3923629638011, 10.3677609209766, 
    10.4813573625864, 10.6196390133803, 10.8102759355055, 10.974064634991, 
    10.6022176529917, 10.4154363269062, 10.0755038403002, 9.66235032661858, 
    9.5113296348739, 9.67222541555976, 9.70500941594864, 9.35722129312334, 
    9.310394244787, 9.30072661188744, 9.10061153373308, 9.06158994818827, 
    17.3986667158327, 17.2908289350552, 17.1945801821965, 17.0462474851446, 
    16.7651288995155, 16.2548085588512, 16.0347539104344, 15.962899768923, 
    15.5444569597475, 14.9672180335633, 14.4804887916743, 14.3919400430312, 
    14.7504465872957, 15.0111559819478, 14.5505990924729, 13.8787638830298, 
    13.1332996098984, 12.6228558281956, 12.5277089718735, 12.8381827590429, 
    13.2582224218438, 13.4458336104685, 13.5034594385301, 13.5649585965064, 
    12.8445094592745, 11.9588078681198, 11.3584996727344, 11.2273122628383, 
    11.4127222167005, 11.3571609365915, 11.3952147168142, 11.1428797211722, 
    11.082152150374, 10.6482669009438, 10.4985327923225, 10.4541519512692, 
    10.5251611764857, 10.7123358432806, 11.0239993909291, 10.8513397767802, 
    10.5956487918495, 9.99779643077852, 9.74809577961225, 9.70748408362822, 
    9.72371725813177, 9.74464400683458, 9.4960092988615, 9.28629450743502, 
    9.26877893791128, 9.05862299307649, 9.12895492094108, 17.1420214298678, 
    17.2829900371906, 17.3087393246723, 17.2486728296354, 17.0011440794858, 
    16.4782139667217, 16.0565730718764, 15.7687474901461, 15.4212534518553, 
    14.5807619897156, 13.8096406550558, 13.6404300760746, 13.8716674546364, 
    14.2181521434489, 14.3674636069559, 13.7456926388614, 12.9287146238982, 
    12.620934648626, 12.5210622869133, 12.8499681193663, 13.2387602566045, 
    13.4836584587051, 13.5595465775973, 13.5045659776322, 12.7193368753595, 
    11.7494657358489, 11.2365835100839, 11.1299466526023, 11.5476039885015, 
    11.540013679942, 11.2621025335698, 11.2691705217837, 11.2300755898304, 
    10.9293051825339, 10.7844155885982, 10.5008113215952, 10.5431831549001, 
    10.6128501846099, 10.4887141899244, 10.6711547929571, 10.3824276101149, 
    10.1349476977509, 10.0004203476571, 9.95475420676805, 9.89843382818683, 
    9.76033474057124, 9.56952644954938, 9.27128670180274, 9.29671606243007, 
    9.0984879401001, 9.0621219646975, 17.026414787745, 17.0410072594216, 
    17.123250299049, 17.1944246010983, 17.0050213602565, 16.7925408455985, 
    16.2744799474981, 15.9539221575813, 15.404352222701, 14.636434176864, 
    13.9510111647121, 13.6960598950177, 13.6212521413131, 13.5605167236332, 
    13.5670930388006, 13.1684119125577, 12.6966849147026, 12.568884001954, 
    12.463890457536, 12.7792525366367, 13.0366853053108, 12.9925942123783, 
    13.086440955705, 13.0501652971849, 12.6470969888465, 11.7796597940572, 
    11.2176664034573, 11.2040089693408, 11.6615236950559, 11.5344242123472, 
    11.0684578944318, 10.9216119233417, 10.8681707127408, 10.8110298080792, 
    10.5707032004115, 10.2668924331704, 10.6060902678271, 10.6956870376481, 
    10.5095831686083, 10.3965259769262, 10.0898213996937, 10.0242859980402, 
    9.83104946059812, 9.63972565176543, 9.68473574371013, 9.42762805962057, 
    9.51028728213071, 9.1967661341122, 9.29594379563266, 9.18335996074945, 
    9.09926290283315, 16.8911927586206, 17.0988317297303, 17.0789336912173, 
    17.0632522044129, 17.2043013366118, 16.9672407869703, 16.5293117873497, 
    16.0399864164282, 15.3163422275315, 14.6598839744083, 14.2051846246886, 
    13.9271739097657, 13.856822227301, 13.7947440909241, 13.4572011022478, 
    12.8834030020328, 12.5327484147049, 12.6102812404149, 12.33514108536, 
    12.5438071935333, 12.8000175284128, 12.8477500525026, 12.784750011728, 
    12.6851418555971, 12.4656478912784, 11.8784757289153, 11.4661364324798, 
    11.3992943819087, 11.6385723344185, 11.474088734018, 11.0869292830773, 
    10.950935093992, 10.5739524216991, 10.4815440166915, 10.2983751341193, 
    10.3029685718137, 10.6047114568918, 10.681618471565, 10.4633699314478, 
    10.2312243646991, 10.100452619114, 9.95168143647944, 9.60130767513428, 
    9.46294770857986, 9.50266736540261, 9.34067306780644, 9.34585607246028, 
    9.16570215237378, 9.35665311350072, 9.2430798447568, 9.18295174198015, 
    16.7478575928025, 16.9125514969124, 16.8454550226438, 16.920938479608, 
    17.187635941952, 17.1069785825889, 16.5045555474336, 15.8667101119503, 
    14.982016882702, 14.3774059655026, 14.1820924077989, 13.9890415193057, 
    13.8508559185097, 13.8198188722944, 13.651383279872, 13.070922631033, 
    12.7097794126774, 12.7260120373225, 12.1859026578364, 12.0525107177775, 
    12.2944914791243, 12.5980345106945, 12.7003666561695, 12.4477824788023, 
    12.1341276667191, 11.8959225250324, 11.4010344619298, 11.4677289280653, 
    11.6102828084425, 11.2493159618153, 11.162242689593, 11.0991280176733, 
    11.1078264023173, 10.6422725635214, 10.6884076182864, 10.7455761888188, 
    10.7487416290988, 10.7260999023554, 10.5305712733222, 10.2440166465773, 
    10.1684920340877, 9.93461318611378, 9.78247667018594, 9.63314024804234, 
    9.60198344727681, 9.52752129082654, 9.58485572012975, 9.39937578560605, 
    9.51503013470043, 9.33007383167465, 9.22701808631436, 16.5154106068662, 
    16.6379813961738, 16.5471927375874, 16.686804532889, 17.02844819543, 
    16.7236153324003, 16.2398004452548, 15.5386735039274, 14.6870519650136, 
    14.2524229622653, 14.1378846887115, 14.1502370032534, 13.8936593509847, 
    13.7899074261539, 13.697456326168, 13.3130158211085, 12.9459998715399, 
    12.874129653888, 12.364738326745, 11.8393928949451, 11.8838632509081, 
    12.3306885063086, 12.885194858132, 12.4676977931176, 12.0951177181163, 
    11.793528570804, 11.698039359724, 11.4718604284803, 11.3820692624808, 
    11.1007940467573, 11.157045647902, 11.3207424943171, 11.2229495836489, 
    11.1391717266093, 11.177740609666, 10.9219663294554, 10.548636505616, 
    10.0858324776237, 9.94382707224849, 9.85101921454667, 9.7130283112852, 
    9.52175965401383, 9.47787306234127, 9.58236175434472, 9.54777971259491, 
    9.38634690850831, 9.22713278597333, 16.1907279426467, 16.0750342960575, 
    16.0053138234291, 16.2323364491046, 16.6024732381152, 16.7429284176083, 
    16.2563179674391, 15.4345867045455, 14.8311126167371, 14.8140130075914, 
    14.5558510654711, 14.2493952917654, 13.751569008146, 13.6633486528532, 
    13.8460174978274, 13.3334079322246, 12.9746584848946, 12.8380621605328, 
    12.3212882972325, 12.1048069076998, 12.0086321216371, 12.0265233866804, 
    12.54249856017, 12.321858596473, 11.9750052183009, 11.6917613907128, 
    11.7666636494106, 11.2147982003942, 11.2873043838266, 11.1662030562212, 
    11.1489313165746, 11.2642672277276, 11.0084762453421, 11.1217695767487, 
    11.004933174521, 10.7726406437135, 10.5257480107713, 10.0035809379084, 
    9.84207807833556, 9.7412913048095, 9.62029366813034, 9.49914492676056, 
    9.44459209921339, 9.4824293756751, 9.40764822860733, 9.35018140310813, 
    16.0805720750925, 15.8896661378517, 15.8244877401913, 15.9278795952628, 
    16.1716323356829, 16.4275241882262, 16.3400788746259, 15.7225282798062, 
    15.2362504459751, 15.2790886227607, 15.2691005154754, 14.4799081628987, 
    13.6092747353903, 13.5297813259674, 13.6257629502589, 13.0900886017948, 
    12.790421135707, 12.5829167969061, 12.3272915370963, 12.529742196893, 
    12.2817422350129, 11.8699137145955, 11.9346683738014, 12.2643123521046, 
    12.2696995686826, 11.8278261551259, 11.5411012989483, 11.1275683043961, 
    11.1316502797306, 11.1689440755194, 11.0713680816331, 10.8821241234668, 
    10.6306250452951, 9.88316702218715, 9.65420825351324, 9.86363385594004, 
    9.70799020293993, 9.47539315353272, 9.45520019835609, 9.39733902325257, 
    9.41226935079088, 15.877314466654, 15.9221807480133, 15.795915248626, 
    15.7404253496358, 15.8508268479731, 16.0788122525993, 16.2947794242788, 
    16.0163981729828, 15.6593831518147, 15.5814369390481, 15.6811088866068, 
    14.6791324210954, 13.3052545566767, 13.4433310239819, 13.3968385985618, 
    12.9434909897411, 12.6694603326407, 12.492891227097, 12.5255152059268, 
    12.7022026965323, 12.5192067440828, 12.0599201054285, 11.733987527954, 
    11.6730401484105, 11.9834940148467, 11.8921757649757, 11.5001669154191, 
    11.3052040067234, 11.2623304534689, 10.989991516549, 10.8404341912316, 
    10.7252711024541, 10.3770129714557, 9.93748085492685, 9.88569813787231, 
    9.78495578880963, 9.62509870076623, 9.46450663261448, 9.43273658431982, 
    9.32692830718512, 9.06336650316979, 16.0547785428618, 16.2782576723531, 
    16.1148709955367, 15.958958155844, 15.8748905981923, 15.8468096897337, 
    16.0485481641078, 16.1616317802892, 15.9725913178235, 15.8769889277699, 
    15.4545634275685, 14.093857931076, 13.0801652070498, 13.2067155608333, 
    13.2486606737727, 13.0097893463621, 12.8338484933589, 12.6418996071754, 
    12.6941321489539, 12.751864207339, 12.5497718592206, 12.1098946773285, 
    11.7161682008317, 11.7401047590262, 11.9692305714876, 11.8391951169104, 
    11.4726327315597, 11.539857589011, 11.4296777158266, 11.0403347951695, 
    10.8973968468366, 10.7252711024541, 9.7139261442914, 9.77591667162582, 
    9.59572584889449, 9.36890592189502, 9.28801707524479, 8.99387069370305, 
    8.69645890179875, 8.50788630481148, 16.3235747199289, 16.2214843013256, 
    16.1884517050051, 16.2043813664919, 16.10503192121, 15.9779495729415, 
    16.1726429168276, 16.2905022781728, 16.2841358760318, 15.8225392670982, 
    14.8282361011482, 13.5829149445539, 12.9630960198964, 12.9888119171427, 
    12.9697277108515, 13.0696396435898, 12.9676281671824, 12.9036495481419, 
    12.8047728771439, 12.5990959510216, 12.439656473585, 12.1083544664779, 
    11.596170789528, 11.5839300943337, 11.7607988246903, 11.8234678820315, 
    11.7947401847765, 11.7061531672498, 9.69470208852504, 9.49671953576043, 
    9.03661528223816, 8.3806347310664, 16.3810035492306, 16.1951768960611, 
    16.0595931639682, 16.0717307352278, 16.0386826512529, 15.9011912168883, 
    16.0137252882225, 15.6485259671631, 15.1386452944528, 14.6478388873338, 
    14.3071476268119, 13.3562722391377, 13.0682676709623, 13.1169309521404, 
    12.8606606402579, 12.7917189999147, 12.8967371523089, 12.8859027558452, 
    12.6455654471233, 12.3774474883727, 12.3874373558692, 12.0547689114613, 
    11.7116099311126, 11.6260686175713, 11.4224231929284, 16.3642244026003, 
    16.0846252600773, 15.874131310123, 15.745677048959, 15.5311589480609, 
    15.2680150562692, 14.5898197316648, 13.8131183128985, 13.4508296667288, 
    13.6513439593644, 13.8125561157962, 13.2717233188454, 13.2828495878733, 
    13.2029641269393, 12.9427830824379, 12.6438752105247, 12.7692647892889, 
    12.8095072944657, 12.5298876394732, 12.3487187444145, 12.3319184930163, 
    12.0986451231287, 11.7615356186717, 11.7953603557967, 16.282192758269, 
    15.9951918466423, 15.8155278113506, 15.3456346910399, 15.070248977604, 
    14.7018571728755, 13.8269000341886, 13.2305336241135, 13.3875434209108, 
    13.4791604225582, 13.4968709591662, 13.2157010514121, 13.3549926838203, 
    13.0973467389921, 12.7411725103378, 12.5952656594027, 12.7366668052195, 
    12.4209991321635, 12.0977748517529, 12.0912961596033, 12.3498202356973, 
    12.0642228228442, 16.1121103370762, 15.9366745817177, 15.9036293911264, 
    15.0004966548482, 14.6623262425794, 14.3744370774363, 13.5896452899778, 
    13.1913393202358, 13.394539806571, 13.3947043883758, 13.3006961521287, 
    13.2860413859825, 13.0776070075026, 12.9430952329784, 12.7082861011475, 
    12.5439645158698, 12.4678987289387, 12.0489272053138, 12.0303163291856, 
    12.1913660852669, 12.1452415529514, 11.930279173746, 15.8709739895333, 
    15.9607256368563, 16.0709181375962, 15.4448482533042, 14.5804494914803, 
    14.0361704197065, 13.5060984817172, 13.2535567887214, 13.4094760105105, 
    13.3789984437501, 13.1852801145624, 13.0348974259827, 12.9905712277084, 
    12.7874990663825, 12.6404177915418, 12.5641979006703, 12.5691259441902, 
    12.0866715562481, 12.0875896568801, 12.0856435181004, 15.8220961543125, 
    15.977104990027, 15.9785426502151, 15.9735640273603, 15.1307216690853, 
    14.0834344505454, 13.4482920736764, 13.3032492403473, 13.4484939085835, 
    13.5018551418862, 13.4126170681336, 13.1416474279478, 12.998411301244, 
    12.824543056807, 12.6384419568459, 12.595843279436, 12.5690741827221, 
    12.339779031772, 12.460894123532, 15.7375219585886, 15.7796025198279, 
    15.6965463814568, 15.7393637027661, 15.4274608933078, 14.2317574567103, 
    13.4238277529172, 13.505033146431, 13.6285040835947, 13.7617783617146, 
    13.7299911971419, 13.4444026690253, 13.3221643302098, 13.161473742442, 
    12.9506991151806, 12.6787982855131, 12.6324427344091, 15.3703446189442, 
    15.3446067801207, 15.4048171857302, 15.5767878479764, 15.850082920127, 
    14.7743906293386, 13.7471850266133, 13.7750540545491, 14.0328683737613, 
    14.1736212611601, 14.0299259418944, 13.837487644526, 13.6294575685782, 
    13.4026686489343, 13.2633054771915, 13.0031798873048, 15.2537485701064, 
    15.2969517970665, 15.311594954613, 15.4145459916085, 15.9388727840005, 
    15.2934753919964, 14.300902417052, 14.1532938717352, 14.4015610577479, 
    14.2218462731503, 13.9676597922407, 13.8424172688011, 13.2202377346266, 
    13.0238667768678, 12.9869181046561, 15.3580041005388, 15.5750023196745, 
    15.3965841799741, 15.2662895587509, 15.7572507615036, 15.4893565140279, 
    14.6507904961605, 14.4692625861413, 14.3857348016506, 13.719862337098, 
    13.6156233049401, 13.4621178056128, 13.1564046036226, 12.9897875761222, 
    15.7121583893142, 15.9219806538605, 15.5144458061023, 15.2010720163883, 
    15.5654647574072, 15.4737246747142, 14.7813349243044, 14.6325627549341, 
    14.0757823532521, 13.4395236470399, 13.2427306294731, 13.2185357700586, 
    15.9211252683283, 16.0292989068187, 15.5278360172024, 15.1540274845577, 
    15.3718255645363, 15.4361442923762, 14.8154726690659, 14.5429192222107, 
    13.9011472813473, 13.5087613244194, 13.380925446828, 13.3869307439064, 
    15.9316341838952, 15.8557429258516, 15.3456900927837, 15.1642630017446, 
    15.1205288869279, 15.2280311248082, 14.6311451967955, 14.2265481265998, 
    13.9166191170381, 13.5544235502593, 13.4801079600318, 13.5744790449298, 
    16.0411571134396, 15.6508974178713, 15.2810564584134, 15.4268785275583, 
    15.0285252091839, 14.7166001571209, 14.4419909633489, 14.106093455423, 
    14.1545992330112, 13.9049000706737, 13.5595487145579, 16.0069723226417, 
    15.4053739243189, 15.2922486528924, 15.4758608011294, 15.1578719751131, 
    14.495278390772, 14.2929390217937, 14.1616743035446, 14.2178815752679, 
    14.0287632562168, 13.6281262588572, 15.6825128630406, 15.1450199549673, 
    15.2703359662479, 15.008782637061, 14.7224769928151, 14.4215671680762, 
    14.1665073911919, 14.0419477732502, 13.9958454672104, 13.7691844515567, 
    13.5054982946314, 15.0721612198838, 14.9068832357479, 14.7807680713527, 
    14.6252097640809, 14.521386645097, 14.3925479492736, 14.2201412034823, 
    14.0815402065713, 13.9965910644537, 13.8739584528394, 15.0996790896686, 
    15.0565081561029, 15.0057669640072, 14.7873282635919, 14.5000974125816, 
    14.4205401177925, 14.3700893111773, 14.330574806795, 14.1577124508528, 
    15.5182449275844, 15.3109959945986, 15.2702804199904, 15.070038223949, 
    14.6341134251645, 14.2460013863936, 14.2497538625728, 14.352859237059, 
    14.2724538529967, 15.9378323383812, 15.6149696413973, 15.4108473483777, 
    15.2764414825984, 14.9400561595381, 14.4505024714655, 14.0735253944336, 
    14.1042250928642, 15.8085881954164, 15.517573198488, 15.325789429658, 
    15.1121922966859, 15.0180525946492, 15.6531024022444, 15.3777775998144, 
    14.8757961032165, 14.7949418328932, 14.3485354894691, 14.4862647825377, 
    14.5546623750108, 14.5863110071676, 14.3249450732292, 12.5653905874609, 
    11.0103213726053, 10.1349855507011, 9.32467097339369, 33.235474527434, 
    33.2332371906284, 33.2316140478617, 33.2313644674359, 33.2407752161715, 
    33.3148420322788, 33.4474479068949, 33.6068541019636, 33.8302155137561, 
    14.4370819175748, 14.518904777999, 14.5707029876738, 14.6493696887267, 
    14.5828190481536, 13.9179524602897, 11.7644855301414, 9.77498769733859, 
    8.64826891901789, 8.18319477571202, 7.89646482100186, 7.5656518276592, 
    7.23320176910747, 6.9648676198367, 6.67677150089755, 33.07963438161, 
    33.0773722305867, 33.0753788625576, 33.0689202545501, 33.0650024223323, 
    33.1043538218449, 33.3095965141596, 33.5954155692134, 33.8429838894356, 
    33.9808623114346, 34.0789606945779, 34.1672477387797, 34.226389180014, 
    34.2617427337786, 34.3109858335825, 0.184203799470898, 0.173662187291327, 
    0.174224256333103, 0.163856572613367, 0.160590569072566, 
    0.162760815870172, 0.154002989057993, 0.171954122638704, 
    0.152250575986985, 0.153618712816304, 0.189291155116613, 
    0.15139538908108, 0.163178751566738, 0.206914579583692, 
    0.140241778028618, 0.167090499189134, 0.164961267498105, 
    0.21526977107483, 0.157981047886401, 0.192117498092487, 
    0.147711466814618, 0.137654189835804, 0.214561370589432, 
    0.162334036807407, 0.208897769132409, 0.125305194451449, 
    0.161232044371871, 0.199420726052982, 0.136501226865834, 
    0.153581488038537, 0.20709761302072, 0.120050906009109, 
    0.159032164029936, 0.181795584096072, 0.114167378133493, 
    0.170349277738538, 0.187898740804831, 0.128309685647487, 
    0.13054551569294, 0.170136078750779, 0.161892217077149, 
    0.112563135693176, 0.162395880150529, 0.169316030820722, 
    0.138008721713799, 0.112633971411455, 0.162610175077377, 
    0.170167786635093, 0.125876387779054, 0.14207361453284, 
    0.160280124213201, 0.132773351194746, 0.145826472001813, 
    0.114850334675997, 0.16123722477851, 0.167690744687302, 
    0.137095381027189, 0.133856450220112, 0.155871112866621, 
    0.153976384254017, 0.151276565702346, 0.126551916430245, 
    0.172867681757206, 0.158824797761953, 0.108270883452907, 
    0.14334849647616, 0.140961576224902, 0.153388194105863, 
    0.183224410347533, 0.156609866159279, 0.134044525966385, 
    0.183718030563748, 0.156847393439858, 0.130365249211556, 
    0.147718211384947, 0.148846671836653, 0.15919389598164, 
    0.191660048263635, 0.16705187561661, 0.094814131586417, 
    0.136900330255417, 0.181090222698905, 0.169073537198843, 
    0.173763950267046, 0.155920345578059, 0.149675841248235, 
    0.168852922265529, 0.188054930422527, 0.172545950572998, 
    0.105934833916568, 0.141466535993899, 0.180222992106607, 
    0.178154470620406, 0.192456364438741, 0.167025806618033, 
    0.0701654118547208, 0.147409929257721, 0.172747029142004, 
    0.189934935215053, 0.168428782941726, 0.144447647421183, 
    0.149165922185195, 0.184870473890056, 0.175551717902095, 
    0.187693882167174, 0.181901129062382, 0.085380718753551, 
    0.150587265205101, 0.178977941866407, 0.197588873725335, 
    0.159709036788432, 0.168083591569032, 0.162355295581342, 
    0.184743374610776, 0.0492052871788941, 0.171425442249257, 
    0.184080337264919, 0.183539867022057, 0.113232300395898, 
    0.159987866971726, 0.192157714046322, 0.207883398076369, 
    0.153951657596351, 0.169076403415523, 0.176781619111967, 
    0.170240563818959, 0.0686929132011141, 0.171082730396602, 
    0.18918220115303, 0.16942815507202, 0.134729304810103, 0.169433070713887, 
    0.190333495653812, 0.062788348651389, 0.214042783358129, 
    0.150413039159616, 0.166346443384452, 0.182858504890894, 
    0.141828607312823, 0.0930079713324195, 0.176523691881166, 
    0.203894341296907, 0.153178092461547, 0.148113549994369, 
    0.175884106085321, 0.172678367741739, 0.081277684158717, 
    0.211447714590441, 0.152186715558094, 0.169062852687806, 
    0.166212413451234, 0.117557329568071, 0.11576803854397, 
    0.180328183857691, 0.0867985954500166, 0.221002790293794, 
    0.140508209879244, 0.152808011652687, 0.172776476827793, 
    0.147333295804188, 0.0983670344794508, 0.207612279368809, 
    0.160727376453536, 0.181700549009587, 0.142782282978725, 
    0.098268322323063, 0.13245978671271, 0.178746206515127, 
    0.102833347461035, 0.227727040494856, 0.136199707686054, 
    0.152067471744646, 0.152504508792809, 0.12848337122123, 
    0.102962970230734, 0.202221303036305, 0.17185774757071, 
    0.0881788243127305, 0.207001971438387, 0.124150831445538, 
    0.0820105014494701, 0.133779069912417, 0.165209033240582, 
    0.103908124902225, 0.219798901187976, 0.139172009935033, 
    0.157781297800814, 0.129491117656844, 0.113928614395465, 
    0.0967086162816831, 0.196448354777909, 0.180045892922411, 
    0.106095887368854, 0.227557357926427, 0.120600689752906, 
    0.0604585017379191, 0.12685243136549, 0.143712835931535, 
    0.093771858382547, 0.212605096472551, 0.15056161837313, 
    0.0710739000979882, 0.178211514979074, 0.112377432401278, 
    0.0980453669300772, 0.0811599721941958, 0.183124815406715, 
    0.180205720386477, 0.100914683349076, 0.227506260680247, 
    0.122988098795628, 0.0396304306654884, 0.128160453134097, 
    0.122424158476894, 0.08245045020098, 0.209374974891419, 
    0.161564273365299, 0.0949013405513899, 0.199703532616915, 
    0.107467058293797, 0.0730769003111377, 0.0656100732371118, 
    0.16598214074675, 0.173209967131829, 0.0882693389146503, 
    0.225907479407993, 0.129902550170347, 0.0584498573250304, 
    0.0404520905559489, 0.142995914056486, 0.105279668585562, 
    0.0661840043582417, 0.204783005949881, 0.167853844275192, 
    0.0959598375370642, 0.207762545857575, 0.104236627664591, 
    0.0540929852675392, 0.0631753438925348, 0.140572617096318, 
    0.162898286998628, 0.0799646301302322, 0.226533411770335, 
    0.139692583627334, 0.0879319734950438, 0.0614985611407883, 
    0.161073348569669, 0.0941068270974627, 0.0496136333950727, 
    0.188554273555273, 0.162195308865666, 0.0826398656079574, 
    0.210434035060203, 0.104900346103016, 0.0750477928166668, 
    0.0622351949258755, 0.0709762909507116, 0.108155940441748, 
    0.147532999456357, 0.0664051165264663, 0.222877815809627, 
    0.141545976331303, 0.0783244304685816, 0.0776922541890645, 
    0.171838990805927, 0.0844844374493383, 0.0480576559565172, 
    0.157578200216535, 0.15548372768778, 0.0696650813819374, 
    0.212619923535714, 0.106696896676141, 0.090624808052101, 
    0.0908129203161157, 0.0795326482731597, 0.0701016113632821, 
    0.122028678993701, 0.0489655617072832, 0.204493920168573, 
    0.131234933848051, 0.0474064209125417, 0.0841334749817962, 
    0.175712183561856, 0.0783370091256592, 0.0952100049179471, 
    0.0594186479190687, 0.116435615018828, 0.149267132022465, 
    0.0623964135654093, 0.209554723099659, 0.0984042426499264, 
    0.0647061312567357, 0.106192245962015, 0.0839775697874698, 
    0.0300972437454015, 0.10025725020495, 0.0505379780682169, 
    0.172369143616794, 0.1227001449768, 0.0251890143919349, 
    0.0906321784429376, 0.176278219082327, 0.0727626881554133, 
    0.0953630191035223, 0.065423056508795, 0.0640178228928102, 
    0.136136579510214, 0.0559137455211707, 0.197118420974908, 
    0.0784138651379723, 0.025301073837855, 0.10310923470375, 
    0.0866918865585642, 0.0067952742235103, 0.111557108153763, 
    0.100681162411048, 0.0653893963109197, 0.129096176941355, 
    0.127280374853837, 0.0361485942994901, 0.0981290032566209, 
    0.173677502426294, 0.0555251445071114, 0.0654943696753873, 
    0.0603074327780536, 0.00555535359539547, 0.122536180514764, 
    0.0601695805418458, 0.171179046120232, 0.0627931996077947, 
    0.00273018320844577, 0.0999459306810189, 0.0930154262667232, 
    -0.000775849769963194, 0.106193352152964, 0.118460041838218, 
    0.0672963300521874, 0.0723444473956687, 0.134964552998289, 
    0.0519039049559349, 0.0895208643873618, 0.168479473422907, 
    0.0287320018365426, 0.0291352733837721, 0.058202207219256, 
    -0.0312821159068278, 0.122166432767891, 0.118524954075709, 
    0.0713543530970024, 0.134668806501593, 0.0704701891582627, 
    0.0192991398535236, 0.103651211285061, 0.0993549879899811, 
    -0.0109449750958491, 0.081260818682711, 0.111971083327801, 
    0.0564761874100563, 0.00471891175641978, 0.135282299487579, 
    0.0445151640938816, 0.0609225429660635, 0.151127006480058, 
    0.0113172319580301, 0.00349728598282595, 0.0654226894101395, 
    -0.0384829705248061, 0.11602131474605, 0.115098798905067, 
    0.0693926380933297, 0.0884734672212462, 0.0987143618025825, 
    0.028656388120004, 0.0940631529717826, 0.1072372203954, 
    -0.0226536199490249, 0.0514073322979836, 0.0752933557418273, 
    0.0539623095061125, -0.0471465398472396, 0.107828880592317, 
    0.133663069216502, 0.0322035645971437, 0.0257908160866148, 
    0.121763165889788, 0.0186609041407531, 0.00904920758908828, 
    0.0711310319201198, -0.0356756980044864, 0.0961720911518984, 
    0.0811249293465514, 0.060721698823757, 0.0274761888928793, 
    0.12163047476813, 0.000842649717443964, 0.0718885264010735, 
    0.0985947084751946, -0.0235725546770262, 0.0231030493481476, 
    0.0427885972963028, 0.0543402600517418, -0.0624956991839961, 
    0.104658882924888, 0.103960222157466, 0.0305548200684797, 
    -0.00888885999569662, 0.0905994808545628, 0.0554479325621393, 
    -0.00628334167927946, 0.0805285294622752, -0.0306501195797449, 
    0.0782213902987135, 0.02501725536279, 0.0632034764906557, 
    -0.0304079277269226, 0.0760856190858634, 0.124478627376268, 
    -0.0281416980106741, 0.0483526823832104, 0.0627181357260565, 
    -0.0153681119890863, 0.00583664879409923, 0.0290746766790397, 
    0.0436524724241223, -0.0529571799769206, 0.088468757487844, 
    0.0264528895180584, 0.0443393378299371, -0.0443951398469488, 
    0.0476877547958277, 0.0927791918648231, -0.0584446735027855, 
    0.0691985281080677, -0.0209408555547429, 0.0614093108328183, 
    -0.0121608452125717, 0.0504528758268992, -0.0546894987344679, 
    0.0821493885784772, 0.0762322745644928, -0.032023512235413, 
    0.0191339891208229, 0.0456316097949948, 0.00981338784806939, 
    -0.0335096668039049, 0.0388181176758792, 0.0360573390521549, 
    -0.0357611760429436, 0.0797985284111445, -0.0512076851818795, 
    0.0587045467431496, -0.065397797834014, -0.00652364985250025, 
    0.0467985409903757, 0.104473656652776, -0.096425574316968, 
    0.025657288245344, -0.00861624977661908, 0.0263651707809889, 
    -0.0253334331418119, 0.00907516427490504, -0.0462014722039374, 
    0.0769716529342288, -0.0252636932943163, -0.0105809187882303, 
    -0.0131366193486878, 0.0364596401363852, 0.0435132462862001, 
    -0.0852457729872494, 0.0535325660636735, 0.0172260972391629, 
    -0.0219741102447478, 0.0751880365374899, -0.0887149207317333, 
    0.0358325054099699, -0.060661892964601, -0.0357365039597183, 
    0.0639635825401007, 0.0538388036968101, -0.100679008977755, 
    0.00971677114864714, 0.00711300575789169, -0.0368915096740946, 
    -0.0227787543258262, -0.0260824761308896, -0.0275901948967136, 
    0.0732826418062881, -0.10797098049063, 0.0159968870309606, 
    -0.0324977084813076, -0.0017680384824872, 0.0369664517693711, 
    0.0536593578872155, -0.102799840512257, 0.0642817692690386, 
    -0.0206989497970053, -0.0116364485917509, 0.0512489195128294, 
    -0.093823944744379, -0.0306263251301896, -0.0461345158657277, 
    -0.028399683935835, 0.0687225536007033, -0.0429632853962546, 
    -0.0800685201055541, 0.00546670302293578, 0.0208280263946933, 
    -0.0921134291204467, -0.0182647063859552, -0.0533865608745198, 
    -0.0167577698400293, 0.0767130152361945, -0.135966216765202, 
    0.0158528426351324, -0.0295187125146448, -0.0289682262037642, 
    0.0537221052365714, 0.0270361134491543, -0.0991433699663469, 
    0.075754715582134, -0.0363986867187027, -0.00816403170708948, 
    -0.00848367791430951, -0.0908813449660715, -0.0864142288489805, 
    -0.0347913796938372, -0.0119123226010469, 0.0669122522733542, 
    -0.115523667342715, -0.0439738667819787, -0.0332275611103391, 
    0.0265238413498884, 0.0130047834025492, -0.0981456176093215, 
    -0.00923435453317378, -0.0830481609594752, -0.0159053238108745, 
    0.0651954578169013, -0.139584172560807, -0.0199261689885201, 
    -0.0200597484851122, -0.0227598441701602, 0.0635853365235066, 
    -0.0160168456431301, -0.088297469860356, 0.0908818421653022, 
    -0.0403683787011137, -0.0206081165300514, -0.0821250165508239, 
    -0.0907328577572787, -0.0973175659163792, -0.0311806706920297, 
    -0.0031572929838182, 0.0641519694590333, -0.141170730381964, 
    -0.012077317149942, -0.062644605875767, 0.0420730092964171, 
    -0.00413301590269735, -0.0681080926255182, 0.0170621132265461, 
    -0.089940231079077, -0.0280463923553461, 0.019842805975024, 
    -0.141786601370123, -0.0529352055001579, -0.0156145943301919, 
    -0.00401904947526637, 0.0707146709957637, -0.0574662555813958, 
    -0.0573145941090735, 0.0972530928952681, -0.0737099068381773, 
    0.0173224026700538, -0.0471743835906405, -0.119658528509091, 
    -0.0825287566664923, -0.0839297505127588, -0.0379657225893244, 
    -0.00877146307871521, 0.0519697700251028, -0.152049524275272, 
    -0.00288877212779126, -0.0516964199906661, 0.0507105267675806, 
    -0.0270788675447195, -0.0375730755141025, 0.0526068177844902, 
    -0.0825292796112256, -0.0573069661360262, -0.0528259580598505, 
    -0.138087944908541, -0.043485420231312, -0.0229049936276168, 
    0.00644758677731948, 0.0714686014632349, -0.0922692515615851, 
    -0.0139235015305815, 0.0870573599701271, -0.107485675520697, 
    0.0387452131766838, -0.0653319927645104, -0.0849595311560138, 
    -0.0534819631876178, -0.0685016686885655, -0.0633437733158561, 
    -0.0305283099405368, 0.029833863813296, -0.164082682745397, 
    -0.00388972059210519, -0.0251914311588449, 0.0634408125737219, 
    -0.05010022504598, -0.00960903632595892, 0.0748794855344169, 
    -0.0974709041504569, 0.0249038941987145, -0.0951694792583196, 
    -0.110737216239211, -0.120873934055974, -0.00905379883161311, 
    -0.0416558011844297, -0.00885293614805156, 0.0592057218565989, 
    -0.120921338646168, 0.0178863801865555, 0.0589589682176603, 
    -0.0956135232514952, 0.0543423224137649, -0.0739254263400234, 
    -0.0319522275525007, -0.017202967005706, -0.0562982645850146, 
    -0.0917947276158349, -0.0691634264823602, -0.0120762277610429, 
    -0.161120450476865, 0.0183419443687077, -0.0136253192969409, 
    0.0753041099040483, -0.0744080980794634, 0.0229734374439729, 
    0.0730726843163108, -0.124698287395194, 0.0553273955092788, 
    -0.113380206110456, -0.0905682258028829, -0.0903362236396513, 
    0.0106846860470649, -0.0752086907784754, -0.0424359477564207, 
    0.0463725476787508, -0.139350658424188, 0.0328827258060875, 
    0.0280500433411192, -0.0610472432123779, 0.0634778582302919, 
    -0.077179099367053, 0.00563163308145658, 0.0115169315853672, 
    -0.0611386977880935, 0.0263596408231415, -0.0872186281775368, 
    -0.112632057530824, -0.0671982223231803, -0.131398185412739, 
    0.0579447038847588, -0.0331641621130096, 0.0724270649074469, 
    -0.102567926827653, 0.0517709154857092, 0.0515324999804156, 
    -0.121395528242473, 0.0697418514207045, -0.106607873929354, 
    -0.0285518981861563, -0.0558158558405589, 0.0109141105194156, 
    -0.0988384243409572, -0.0756940515395511, 0.0366405548348554, 
    -0.140066898483936, 0.0566447080378116, 0.00237916273222745, 
    -0.046156678423381, 0.0714344955168246, -0.0821748098407308, 
    0.0298222580658081, 0.0185140724857029, -0.0904493949334611, 
    0.0576432951475667, -0.061800339767689, -0.129390436975861, 
    -0.0601693609448898, -0.0945519819908146, 0.0764138130833886, 
    -0.0704013319624568, 0.0615945985699218, -0.120590938290081, 
    0.0692516850539735, 0.0222057805738307, -0.0921308176693301, 
    0.0670019938196372, -0.0960981272820943, 0.0106630223063458, 
    -0.0277337618668634, -0.00700845245551183, 0.016570314071974, 
    -0.0941029304081838, -0.100003156490844, 0.0139260345816423, 
    -0.114623990845124, 0.0916165643505669, -0.0217867568908636, 
    -0.0647537400893606, 0.0716616376352864, -0.101721132658711, 
    0.0454926549571329, 0.00950480350820035, -0.128312231389747, 
    0.0662820875489221, -0.0467691309195726, -0.114854837290851, 
    0.00209463887673366, -0.0695983711549058, 0.0664061209288214, 
    -0.0963238751230801, 0.0575708292513872, -0.121139281396082, 
    0.0831494041479255, -0.00328529452250946, -0.0794491378180537, 
    0.0627428227792121, -0.0987451253972083, 0.0235881704109243, 
    -0.0258898257552623, -0.0503973495925319, 0.041840917397141, 
    -0.073967224112921, -0.111685821337356, 0.00388584441999817, 
    -0.0830665411336611, 0.105796802125088, -0.0554379808806026, 
    -0.099376433838146, 0.0633401972202776, -0.121629495133962, 
    0.0547154644495554, -0.013100773966936, -0.140510934187557, 
    0.0641955314550247, -0.0343366764894766, -0.101321824809143, 
    0.0321370886316232, -0.0549364686056685, 0.0373707463434982, 
    0.00899240011588635, -0.0981242971287411, 0.0535066188913864, 
    -0.100231910375376, 0.0961055747919152, -0.0210494556511873, 
    -0.0979425575035012, 0.0572876712915687, -0.116213546325311, 
    0.0287336705033529, -0.0317368511451552, -0.113482610888445, 
    0.0493815376476787, -0.0532688542215058, -0.101151527813382, 
    0.0257642679291243, -0.0715952777421038, 0.0902524454885004, 
    -0.0761419654555244, -0.117518126197126, 0.0605765499608669, 
    -0.122614698213455, 0.0617589230682637, -0.0196677424409418, 
    -0.134807223738301, 0.0612534609699923, -0.106582541154529, 
    0.0263682229801723, -0.0545116938252011, -0.0119670386155228, 
    0.0210324344002463, -0.0999773428537326, 0.0355853274422738, 
    -0.0716990315206009, 0.0987338559375959, -0.0467074267374717, 
    -0.125058197291823, 0.0493663696498207, -0.128030160363272, 
    0.0345606318595247, -0.0401747134361807, -0.151773501469663, 
    0.0513525433654783, -0.0395344169378861, -0.0986908842242778, 
    0.0191123484272005, -0.0780114473885804, 0.0563164828336237, 
    0.0125226081207994, -0.0763149464362729, -0.106390121539842, 
    0.057458516068081, -0.0919051886995873, 0.065556796023707, 
    -0.0314490104719658, -0.143008400262967, 0.0518242201154118, 
    -0.116896571135865, 0.0145042995921747, -0.0556138433131153, 
    -0.0802602040729942, 0.0279440944521899, -0.0940017442312544, 
    0.0249543839121857, -0.0737844376436862, 0.0851209716851889, 
    -0.0622889960425531, -0.128983471352243, 0.0453439133198611, 
    -0.122846484106921, 0.0362364638560414, -0.0387243486907361, 
    -0.146189480524734, 0.0486398402286686, -0.105402801904715, 
    -0.0144258755566234, -0.0745393109528798, 0.0118754252185149, 
    0.0196993126069349, -0.0715748460813559, -0.095338036529041, 
    0.0425727876387108, -0.0759287320246869, 0.0635608159957966, 
    -0.0504760475686421, -0.143266144929426, 0.0389274145864491, 
    -0.121453697485413, 0.00533404060543072, -0.0540693940074245, 
    -0.131982545323907, 0.0254498040683127, -0.0896312307024445, 
    -0.00877237807073237, -0.0809918898329468, 0.0586540036368048, 
    0.0181725446119013, -0.0675971402142466, -0.10792707319457, 
    0.0380383988322161, -0.0986955240305047, 0.0285179588761979, 
    -0.040221559780687, -0.141350207445247, 0.0359868023494775, 
    -0.100909587100124, -0.0492196376055396, -0.0698150497739603, 
    -0.0412106026427256, 0.0268562966379871, -0.0485347400372419, 
    -0.0832743681419109, 0.0190808173851916, -0.0750126377142107, 
    0.0555110756348929, -0.063816681329824, -0.124835364325109, 
    0.0311959400038175, -0.121486349537205, -0.0165042595656183, 
    -0.0448135272520196, -0.138160744732229, 0.0128403741582704, 
    -0.0908151912797684, -0.061868462776399, -0.0791442876200261, 
    0.0251433508970165, 0.0248524764097781, -0.0739567061121787, 
    -0.0926686280503004, 0.0284305696444748, -0.0788349158448491, 
    0.0153387601717186, -0.0546105613598606, -0.13426607171346, 
    0.0207763582025833, -0.0982826459780162, -0.080496077737522, 
    -0.0694972127393464, -0.0876810654368098, 0.0223231411277673, 
    -0.0727399603499895, -0.0277947496951587, -0.0756833949201961, 
    0.041052050385927, 0.0291664666066692, -0.0724905101309894, 
    -0.101247231199151, 0.0254150269199767, -0.0979287867181328, 
    -0.058819117562948, -0.0442884925681039, -0.127871064351194, 
    -0.00394109063080159, -0.0916405551986433, -0.11223188733241, 
    -0.0755925098851227, -0.0047406812228776, 0.0360037943127994, 
    -0.0798905473321642, 0.00695649601614232, -0.0738206820689741, 
    0.00521708095424712, -0.118082769604813, 0.0113525967225221, 
    -0.089607061723868, -0.121718919824751, -0.0693138929830532, 
    -0.110754803877268, 0.00582283982412153, -0.0733362570422552, 
    -0.0884769797697492, -0.079221622165444, 0.018134389216393, 
    0.0428491876072131, -0.0818276587571671, -0.0922827232491537, 
    0.0203070772553392, -0.0764800560946216, -0.101104113136206, 
    -0.06340697194452, -0.120447599707085, -0.0173943454368754, 
    -0.0744031675878528, -0.145793301848548, -0.0286633190261068, 
    0.0288768873944031, -0.0592926133615877, -0.0396682318015084, 
    0.000831411781797971, 0.0336233672203545, -0.0986775880885602, 
    0.00800503390441768, -0.0721536930232176, -0.185713706506675, 
    -0.0820905081052652, -0.109534804611736, -0.0117945347876345, 
    -0.0782715757297764, -0.140000151101827, -0.0804857805299504, 
    -0.00738800309330959, 0.0483281487396001, -0.0730630834765355, 
    -0.00160108446579437, -0.068811041272705, -0.120399385175877, 
    -0.108569123605063, -0.0240025829830891, -0.0645676842848144, 
    -0.169750821093407, -0.053987723097003, 0.00885088441379709, 
    -0.0665843050255878, -0.0850530915838672, -0.00513834825593147, 
    0.0547557787400508, -0.0852110629396982, 0.00501300764833764, 
    -0.0625314217527688, -0.240909818330259, -0.100795265879382, 
    -0.103978515679948, -0.0235669367960154, -0.0591402275508243, 
    -0.158984870385006, -0.0309523932513482, 0.0320627692989955, 
    -0.0468224555702594, -0.0462835134953149, -0.112593697136982, 
    0.0342656899614687, -0.092036993434255, -0.0254222475390964, 
    -0.0534069790399331, -0.21700513736295, -0.071850809554913, 
    -0.00925460421010234, -0.0766244499253985, -0.112376568296741, 
    -0.0194506308679804, 0.0481967004948596, -0.0614566050184401, 
    -0.022716648089078, -0.250688102471763, -0.0968291677283393, 
    -0.0327182456151272, -0.039925527213802, -0.157846147276555, 
    -0.0509082146569228, 0.00741771063366725, -0.0427235978781133, 
    -0.0786793194307225, -0.0912047209560415, 0.0614292266498716, 
    -0.0726089410029178, -0.0317265146526091, -0.262070149013523, 
    -0.072700993630481, -0.0241775770483822, -0.0562569133049363, 
    -0.11804985420016, -0.0386878293274549, 0.0240773197060854, 
    -0.0366861183041326, -0.0691092566688488, -0.222234050845125, 
    0.0182885026755572, -0.0836633070519715, -0.0414297750656762, 
    -0.183823869385943, -0.0643197499225614, -0.00941924479575522, 
    -0.0570136216600023, -0.0923775741264913, -0.0782678624004196, 
    0.04849841732182, -0.0514472706919129, -0.0576276958571066, 
    -0.263002094357013, -0.0744148478466012, -0.0419891536404849, 
    -0.114556616622473, -0.056822025151999, -0.00156819329799373, 
    -0.0327034866694048, -0.0941555344906596, -0.183026504787625, 
    0.0452150534952572, -0.068788786954436, -0.0487324687845865, 
    -0.222437123110418, -0.0689338353372484, -0.0265498811328161, 
    -0.0504029482171636, -0.103209032129933, -0.0809411345294359, 
    0.0155521391397225, -0.0382555107956358, -0.0864763921940838, 
    -0.233345139302708, 0.00473376817407742, -0.0818177010855004, 
    -0.0615108919606971, -0.1200547529399, -0.0633627276849959, 
    -0.0160035366786353, -0.0418900925993683, -0.100307264693535, 
    -0.155246567021504, 0.0298771472773422, -0.0571830451148588, 
    -0.0605557997009286, -0.225617435389114, -0.0718034115453472, 
    -0.0583362739427952, -0.111887382454076, -0.0874437768957581, 
    -0.011149477420797, -0.0393143165972609, -0.0978587642336468, 
    -0.197246077269951, 0.0183603073842388, -0.080965020443421, 
    -0.0680048950301635, -0.139848457243484, -0.0618523730594057, 
    -0.0317214330407303, -0.109655294774159, -0.143692739067701, 
    -0.0034923983923745, -0.0482455018840443, -0.0732904373074592, 
    -0.204094020492329, -0.0323403180303077, -0.076180060751034, 
    -0.0992389711839998, -0.106889227254484, -0.0831435035703615, 
    -0.025092327147725, -0.115830640744787, -0.169679914468107, 
    0.000814043415287718, -0.0801322282859391, -0.06514508152516, 
    -0.14810031027996, -0.0577430015105962, -0.0663865714326584, 
    -0.121635952151321, -0.142554374320272, -0.0228929553751127, 
    -0.0480257074786502, -0.0842212828106146, -0.181978491631911, 
    -0.0359364204061233, -0.0830351281343312, -0.119311080912215, 
    -0.104302770193779, -0.0776636476981192, -0.0384752430732838, 
    -0.146038555720142, -0.159149934030916, -0.0207857232684117, 
    -0.0651337724891664, -0.144830232663852, -0.0457435935163243, 
    -0.0702114101454053, -0.113322646676041, -0.118043944724157, 
    -0.137679283560455, -0.0299118398773687, -0.114427589934728, 
    -0.163889157722871, -0.0422198715292113, -0.105522478265338, 
    -0.11256127134368, -0.0713139068427514, -0.0705180290420854, 
    -0.167653118184374, -0.158823125173369, -0.0240876588831544, 
    -0.0762815382156035, -0.146466693256214, -0.049858571588871, 
    -0.0822242363667829, -0.14189779575031, -0.10484741639339, 
    -0.119461606947633, -0.0388609454415019, -0.158333812035759, 
    -0.160009666723165, -0.0272493739610903, -0.0830829513964145, 
    -0.127652317078022, -0.0438254808594536, -0.065971276360114, 
    -0.113760200744137, -0.172645960857923, -0.152760162355408, 
    -0.0238794527707222, -0.111065960335709, -0.146816349305058, 
    -0.0516381041266065, -0.130885740093913, -0.102725654303724, 
    -0.103227437131621, -0.058018130332693, -0.189646397450595, 
    -0.154990864462805, -0.0101753116937106, -0.078188896645641, 
    -0.140578862789944, -0.0470704283380568, -0.138214616208713, 
    -0.147552648800658, -0.133329314312377, -0.0290478297393912, 
    -0.154510894456275, -0.150783889626092, -0.0317543126602122, 
    -0.103103336573069, -0.122702388749842, -0.0409949280848642, 
    -0.0761605466947052, -0.0869813529194837, -0.202169722009902, 
    -0.152707472181113, -0.00436928376303103, -0.0971418563347992, 
    -0.142920158716826, -0.0511778818133702, -0.131730435572141, 
    -0.116977632343048, -0.0943717186187552, -0.0393924016633262, 
    -0.189391828678688, -0.140984748471197, -0.0116461195902404, 
    -0.0873039021376547, -0.145276898961786, -0.0379278782768024, 
    -0.100867346178206, -0.177887904331127, -0.117225062289972, 
    -0.00378864339007082, -0.121540644155522, -0.135349237744956, 
    -0.0447963430222736, -0.109022750137963, -0.124937230091434, 
    -0.0528002561790067, -0.0665342801844544, -0.0623106194351945, 
    -0.213457815467474, -0.124204122202403, -0.00116788013461638, 
    -0.0898801158980123, -0.148092996843968, -0.0425599658563102, 
    -0.0966119632243325, -0.135933459269074, -0.0691331585279739, 
    -0.0100496576253488, -0.150487485103986, -0.124111258398014, 
    -0.0293347159522745, -0.0912861358366794, -0.155773144421932, 
    -0.0488645523680635, -0.0769290158405365, -0.202170014842543, 
    -0.0788628905598539, 0.00301395418833189, -0.100087130013855, 
    -0.131710494500459, -0.053125832153616, -0.0873272469739566, 
    -0.134812224107905, -0.0675369029490125, -0.0304814282745562, 
    -0.188846063663083, -0.107317305836236, -0.0106565050022847, 
    -0.0858433601245675, -0.166303696769175, -0.0422981593572408, 
    -0.0733630817403853, -0.16162123480762, -0.00414772877851534, 
    -0.120580719100232, -0.119873835981437, -0.0496486186400486, 
    -0.0824990980077878, -0.161355538893252, -0.0593093197139655, 
    -0.0503582310022727, -0.20717014845941, -0.0743916850196131, 
    -0.000574555931349909, -0.0879690256603527, -0.148527950020058, 
    -0.0446162955812361, -0.0692889672383146, -0.156740255972773, 
    -0.0692976904392181, -0.0210764358656204, -0.156646672928133, 
    -0.104220504979308, -0.0291218196699272, -0.0843639901117338, 
    -0.171223420070589, -0.0421414416103593, -0.0455872714163181, 
    -0.192461023165392, -0.0438327140819194, -0.00387104509057642, 
    -0.0976408002551659, -0.132990507198884, -0.0433526591784469, 
    -0.0755495271219862, -0.172094373209996, -0.0599685990565685, 
    -0.0373760618617313, -0.184643537024813, -0.0803130999311522, 
    -0.015523662350618, -0.0933794579930082, -0.152645327987172, 
    -0.0341624370500205, -0.0329896531094418, -0.187609638697191, 
    -0.0850574619411161, -0.0145117091227391, -0.120022398029619, 
    -0.107894880341294, -0.0290599559593173, -0.0901762588966588, 
    -0.177838321847181, -0.0392875716159412, -0.0341761319584694, 
    -0.186950946680223, -0.054464013945065, -0.0147642337354556, 
    -0.0973259976389711, -0.130730332666634, -0.0350236202841205, 
    -0.0386079175247009, -0.175734312446425, -0.0864590367376897, 
    -0.0245108575714895, -0.142493762302752, -0.0220191813679335, 
    -0.10970143354428, -0.153574954745573, -0.0333656719942409, 
    -0.0229210297423413, -0.181050357104554, -0.113167350265502, 
    -0.0176704760649394, -0.101170141859324, -0.102820574585799, 
    -0.0374023868765431, -0.0659295856982114, -0.162385243793116, 
    -0.0552237059422921, -0.0276230454423536, -0.150654815748403, 
    -0.0245056447221779, -0.120658176455951, -0.128265782647526, 
    -0.0404100475858416, -0.0325810844989242, -0.163638341587886, 
    -0.12811497100919, -0.0205196490196923, -0.103416004778138, 
    -0.0377667797190979, -0.102583948813391, -0.128044990981025, 
    -0.0333560583835093, -0.032994291586574, -0.14898050552418, 
    -0.141295810330893, -0.02744343520178, -0.123693616002781, 
    -0.0890739522139528, -0.0508563967021742, -0.061410221313085, 
    -0.14060350495761, -0.107813427051593, -0.0324106304742548, 
    -0.109485528708798, -0.043207223834606, -0.129114192918037, 
    -0.091020977580501, -0.044180644244019, -0.0603681538933241, 
    -0.141547408673872, -0.152621676040537, -0.029079753664867, 
    -0.116134754112062, -0.0489997520186545, -0.0970041409368702, 
    -0.106018706452163, -0.075012581886117, -0.0615171029079487, 
    -0.11385442087696, -0.0538322708591475, -0.133596212318999, 
    -0.053294639256838, -0.0644481884839746, -0.094473262302992, 
    -0.12662554930735, -0.137056381502807, -0.0397609127233976, 
    -0.11480786649599, -0.049192802666884, -0.125217327467468, 
    -0.0702127574848815, -0.0719685445293975, -0.105532038278076, 
    -0.122744442800082, -0.0576945622269374, -0.131115062730071, 
    -0.0147807268570782, -0.0678666369816351, -0.121331942402815, 
    -0.104061037295196, -0.105318524030095, -0.0640150676254498, 
    -0.1225746833825, -0.0594831706989, -0.13287918741207, -0.04737470121864, 
    -0.0874017368530655, -0.142546532125857, -0.12940016659289, 
    -0.0588857992595335, -0.128970025032511, -0.0612003433291023, 
    -0.137420478599403, -0.0724515402226027, -0.103344272485216, 
    -0.100424326181848, -0.131119136040273, -0.064418244380088, 
    -0.136489380002163, -0.0108042927996322, -0.0882411183817182, 
    -0.164694526364041, -0.118509026464329, -0.0630030489142508, 
    -0.131095868220939, -0.0621735645969828, -0.142357898694851, 
    -0.0555890915347576, -0.117501044109486, -0.133647618825048, 
    -0.141570139359228, -0.0667988548564104, -0.130668085241777, 
    -0.0757853591713728, -0.172480797401531, -0.0944294377052398, 
    -0.0755259006921628, -0.142425142107165, -0.0662432332775092, 
    -0.142217517309758, -0.0146604903104821, -0.112462502894024, 
    -0.158592530419055, -0.131687257239197, -0.0674305325818074, 
    -0.126940012846544, -0.0709880582903394, -0.168215864417187, 
    -0.0733822609955427, -0.0936795933625382, -0.152503324740511, 
    -0.0725463990845068, -0.129728263973984, -0.0929567934951734, 
    -0.174315438950934, -0.109065761591596, -0.0680567964607725, 
    -0.143797728189277, -0.074334033030807, -0.152453016916674, 
    -0.0203010688985004, -0.122228238925716, -0.150133997854439, 
    -0.0768890504873992, -0.123924353864374, -0.0849580963964596, 
    -0.173235897678908, -0.08095368937986, -0.0756228026936446, 
    -0.157139523503083, -0.0815348309118098, -0.122872942730412, 
    -0.151771743655868, -0.128340897574786, -0.0725721257298116, 
    -0.147712347180682, -0.0940851512079345, -0.156364200299458, 
    -0.0299325013117996, -0.103689951216206, -0.154359580085947, 
    -0.0907810917332375, -0.113956715083562, -0.162232211262475, 
    -0.0966101169842766, -0.0803494286428693, -0.163684817399111, 
    -0.0924666672762129, -0.121974628977548, 0.00655307997527613, 
    -0.135061824012785, -0.131166874099207, -0.0931064654462107, 
    -0.140691187286529, -0.150381401956915, -0.0569702258552868, 
    -0.113149861833926, -0.157989236397991, -0.0970953908064361, 
    -0.110847886330635, -0.148456199671204, -0.0988971218288006, 
    -0.116183489458095, -0.168059052337665, -0.12690803689895, 
    -0.00888032132692628, -0.137124127593981, -0.13252656278342, 
    -0.117909004493484, -0.134822774181958, -0.143078241984586, 
    -0.0627403627792902, -0.15160718848078, -0.17035227541399, 
    -0.126364546864627, -0.146702698822224, -0.0972931444553376, 
    -0.156025238374041, -0.167685261903303, -0.132993913807509, 
    -0.00957929543386232, -0.173482663600657, -0.147350626245082, 
    -0.145753356850318, -0.156904314574924, -0.0630014153325932, 
    -0.180949701405943, -0.175726453379347, -0.142450549961157, 
    -0.185358954507481, -0.114615634555208, -0.167970379371614, 
    -0.171526617361112, -0.0117150656184447, -0.184846127602329, 
    -0.156859148209489, -0.160770205010928, -0.200923957408659, 
    -0.0756600303375617, -0.173759511721809, -0.188282553624685, 
    -0.190550564283689, -0.128623543245029, -0.170055186925047, 
    -0.213073121609967, -0.0192290877742008, -0.150133825286839, 
    -0.193266842959912, -0.204576913486495, -0.0852858746202378, 
    -0.170925243503312, -0.217040487898327, -0.115576631979502, 
    -0.17914092944421, -0.214784252699751, -0.0283201471095463, 
    -0.142832799278532, -0.213248190722766, -0.0779365609672175, 
    -0.169703054731334, -0.211685101248258, 0.00565245467091932, 
    -0.099701722981906, -0.196683505486143, -0.0408652133028302, 
    -0.139051800769778, -0.206135766742852, -0.0593836279784703, 
    -0.174289885170483, 0.00312645498340617, -0.0976085763747788, 
    -0.200169510623461, -0.024535636856033, -0.147625259633211, 
    -0.0475411688674998, -0.177273993086656, 0.0132801214011825, 
    -0.105409647524033, 0.000392883750071251, -0.149835928366134, 
    -0.0511372992579538, -0.098551454355191, 0.00110847202564375, 
    -0.0421208128691714, 0.0235125097359769, 0.00810930949414044 ;

 NLmodel_value = 17.8503597407106, 17.8193642555481, 17.8543400413646, 
    17.4276819634862, 17.4017312411222, 17.0055186663776, 16.8892228363505, 
    16.6550101112547, 16.6727579687687, 16.5127129703001, 16.4957469743843, 
    16.4537188496371, 16.0928224214996, 15.9077490036503, 15.3178399173616, 
    15.2137826643969, 14.7701069954081, 14.5745962210981, 14.4684744128471, 
    13.9372858504207, 13.4398422633629, 13.3560566764397, 13.4007382080576, 
    13.5740392396616, 13.5901561049451, 13.6777261953069, 13.7064379246056, 
    13.2831157816019, 12.66909161519, 12.2993236199165, 12.1580834600032, 
    12.1781024214249, 11.9925469119524, 11.5290434357383, 11.0823708117183, 
    10.9363632779115, 10.6903465702308, 10.763236423528, 10.7851981650146, 
    10.9627094607907, 10.7891409942332, 10.7328685556861, 10.7938249687936, 
    10.6982203903337, 10.5967222738595, 10.4229846920914, 10.1750171970436, 
    9.92133732834223, 9.67830749824837, 9.54344660336579, 9.35664587404753, 
    17.78623832546, 17.7542546281895, 17.8284117826359, 17.6804281095445, 
    17.1113177468432, 17.0682179915573, 16.789584044299, 16.7091896199551, 
    16.6031397352502, 16.5572064051071, 16.4304960434169, 16.3363568186587, 
    16.1722555624937, 15.9411377614162, 15.4738826211477, 15.1698276964978, 
    14.6033417164072, 14.5915017268275, 14.7821085099822, 14.2280506909117, 
    13.7984915149185, 13.6932245125357, 13.946256525847, 13.9834173049776, 
    13.9726612643943, 13.9217191078455, 13.7032176262609, 12.8876930077719, 
    12.5389923923367, 12.5590619866189, 12.1338222201189, 11.928158074274, 
    11.7842199087432, 11.7151279580624, 11.3225137628758, 11.1416426249549, 
    10.9443387635713, 10.9977561310098, 11.2346143682124, 11.1673853953265, 
    10.8887797463883, 10.8232329526459, 10.8775817464059, 10.7636254334987, 
    10.6080513272022, 10.44991602153, 10.0759207585652, 9.86757995150442, 
    9.69778483329099, 9.69736128557445, 9.58795311049037, 17.7080164152781, 
    17.5459508565642, 17.5668505754436, 17.3568238646189, 16.993599190857, 
    16.6614463355263, 16.4266132028243, 16.5924946027847, 16.5075523302679, 
    16.5833523211421, 16.433039171903, 16.462523860856, 16.2986786218724, 
    15.9805039261469, 15.7045440840628, 15.3257465769989, 15.0194939680982, 
    15.2201047245685, 14.7203070699576, 14.3865633790296, 14.1335669238706, 
    14.0349299179905, 14.1595293758327, 14.0553664616844, 14.0106261668248, 
    13.660721138173, 13.1139429087822, 12.5684669667236, 12.5340080179973, 
    12.4966148476501, 12.0642511765317, 11.8634986560973, 11.9261317315055, 
    11.9534859004051, 11.4696899395643, 11.3794351811205, 11.1838199373005, 
    11.2661592931694, 11.4724127522811, 11.1340693893616, 10.8172119033441, 
    10.8654085976016, 10.7780453116189, 10.5435979134583, 10.4378751816582, 
    10.3390367098304, 9.92481050839457, 9.78928939189919, 9.67324692197197, 
    9.78819644075969, 9.7032533188978, 17.8461510318323, 17.5343389485913, 
    17.391900005185, 17.2187760494824, 16.9105230137567, 16.5937322233199, 
    16.2983296924417, 16.4733498267078, 16.4379170898389, 16.5637914036273, 
    16.4234482825667, 16.3737237494425, 16.2321931711053, 15.9545601437475, 
    15.7443251592032, 15.3315057781708, 15.2585678372505, 15.1487893728037, 
    14.6840549538672, 14.107702882671, 14.2470942283893, 14.2392729754185, 
    14.1583199587297, 14.0023382965554, 13.836510235937, 13.3273345051136, 
    13.0056812379618, 12.493365325114, 12.4115607488801, 11.9908589504001, 
    11.718919669789, 11.4916286073327, 11.46954268037, 11.8026530860085, 
    11.5074841919094, 11.423618309285, 11.2378107840847, 11.4405021606469, 
    11.4600381038421, 10.9848151739476, 10.8618902439017, 10.9472884208258, 
    10.5860775087212, 10.2581545995435, 10.0832596146775, 9.82609806483965, 
    9.60243887791832, 9.62511897156371, 9.78870616229214, 9.80202340314271, 
    9.62920200692774, 17.9114208216967, 17.6782909176303, 17.2819200235319, 
    17.0361011029422, 16.8401982558295, 16.6256609016455, 16.3928487297027, 
    16.429057957143, 16.4396316887959, 16.4410157977847, 16.3116814011706, 
    16.3154908797639, 16.1301474062748, 15.9032492026344, 15.7914478667821, 
    15.5161681005243, 15.4714853574944, 14.3436033523869, 13.5890320443316, 
    13.3813886795018, 13.5774328392176, 13.7809658629896, 13.8221944155036, 
    13.9080776310354, 13.7608374072008, 13.3152036814697, 12.7703387715772, 
    12.2130844245627, 11.8679657371617, 11.4944883763177, 11.3862164159023, 
    11.3655040301587, 11.1909186477714, 11.357487912583, 11.290370325348, 
    11.2412240411407, 11.0901478168104, 11.1657685825167, 11.2439797223129, 
    10.9508953866386, 10.6821345135173, 10.5361541846568, 10.1979617565869, 
    9.98469845054406, 9.94912658048825, 9.63359428768864, 9.54554151378842, 
    9.69284495312533, 9.73707794004013, 9.62566304552345, 9.6065363666667, 
    17.797045741543, 17.5951670329857, 17.2159235712024, 16.8572640515532, 
    16.8706739953938, 16.5758007195156, 16.2674504394232, 16.2978436111923, 
    16.2134073219153, 16.1158448702509, 16.2172316233392, 16.1244094663006, 
    15.9605121158289, 15.7846872968632, 15.783323953581, 15.4739851095658, 
    14.8126386051737, 13.7889875244002, 13.1937404255727, 13.2217428836456, 
    13.3727134950009, 13.7559516894654, 13.6977888799019, 13.7708039835795, 
    13.647172284707, 12.9828219389465, 12.4403286897764, 11.7026035015917, 
    11.3965099916137, 11.3373605934843, 11.253836544449, 11.4136556016609, 
    10.9414107139635, 10.8977786713088, 10.8580433282122, 10.7766130462687, 
    10.6480210806282, 10.7447617663704, 11.0400372186833, 10.8595498586308, 
    10.587487051165, 10.2946618709497, 9.92703322252793, 9.88709924734134, 
    10.0130232745904, 9.65947491991373, 9.5659912191405, 9.72735571591937, 
    9.65978215725963, 9.61124162661307, 9.48152741293185, 17.7903232441273, 
    17.5059628094998, 17.2756332133434, 16.9354487041527, 16.9988238135944, 
    16.6761143214815, 16.3985929137516, 16.2509065060954, 15.9574836824959, 
    15.9079343346214, 16.0373041359091, 15.984588044998, 15.7303781295054, 
    15.5549528982856, 15.3856367905075, 14.863539347573, 14.1954944245346, 
    13.3982840582215, 13.0333757424945, 13.135405104057, 13.280373523453, 
    13.6817669489062, 13.5657409266276, 13.6283029374253, 13.5211093418819, 
    12.7031407911791, 11.9538500311589, 11.1668963317514, 11.3660747993183, 
    11.1694255204883, 11.2762225179785, 11.4480447717485, 11.022241278616, 
    10.7136225262325, 10.5665269068912, 10.6246277141703, 10.6384986386983, 
    10.6068809087994, 10.8218032351998, 10.8575287551301, 10.7359645544998, 
    10.3548214020536, 10.0400161007419, 10.0074729598754, 10.1287088428085, 
    9.81497778426771, 9.53496105415486, 9.6270719614086, 9.46145163876458, 
    9.65875191625077, 9.77588919192158, 17.7116484888206, 17.6771581412361, 
    17.3219487612094, 17.2458210098791, 16.8841691768387, 16.7311373413773, 
    16.2067780639548, 16.0320201606828, 15.7229061818235, 15.8191558824344, 
    15.9403938698801, 15.7907106354923, 15.5849476571426, 15.51744831106, 
    15.3555811799818, 14.3591731273597, 13.6298862379952, 13.0942546718574, 
    13.135897042716, 13.2913605436677, 13.3550850812397, 13.5158415560855, 
    13.4603397125454, 13.6483454779775, 13.3576180240404, 12.3671338573822, 
    11.5262314296308, 11.149038498773, 11.270028436982, 11.1538692037399, 
    11.1610868001642, 11.3136176231398, 10.997107227453, 10.4412537516448, 
    10.3207541044676, 10.4530282069205, 10.5850103321791, 10.7749443503919, 
    10.7529196591543, 10.9141635725894, 11.0630319279201, 10.7358828226753, 
    10.3775048149202, 10.2792947671977, 10.1614023363786, 10.0487473064073, 
    9.68540022642446, 9.47801981528641, 9.20270429644025, 9.58041416590621, 
    9.80873145928602, 17.9080898204861, 17.6454998627146, 17.5249058991049, 
    17.118589548664, 16.8184958598448, 16.3770794377714, 16.290813346571, 
    16.1311650450167, 15.8698764369826, 15.841727170307, 15.6870929364536, 
    15.311851787269, 15.1929059928634, 15.4495177230598, 15.4267407535255, 
    14.3068501853335, 13.2610305874218, 12.8418368052907, 13.2123605646537, 
    13.4693830219465, 13.5174045583249, 13.5328721626988, 13.5190571567445, 
    13.673353507381, 13.1760508775773, 12.1662902070976, 11.312544141626, 
    11.225978315485, 11.2512123125036, 11.2048973877085, 11.1214244663425, 
    11.1707714042929, 11.1213681443938, 10.5247530852681, 10.4002153573233, 
    10.3812621420302, 10.4476437332141, 10.685563738944, 10.7567869714186, 
    10.9891603466028, 11.0751349682024, 10.7494453204837, 10.4180738535929, 
    10.3875133875124, 10.180612626077, 10.0728859929323, 9.79571605433243, 
    9.37627775342143, 9.03257583798311, 9.66158937236226, 10.0158746865946, 
    17.7563407819754, 17.823948729732, 17.5590959508169, 17.2966125556548, 
    16.945571172266, 16.5050088965958, 16.3595992624997, 16.0183693449192, 
    15.8750720681533, 15.6804028606444, 15.1376454749464, 14.7416876635494, 
    14.6684153748176, 14.8503903609522, 14.8847638890016, 14.0460550870161, 
    13.114223655634, 12.8636310668878, 13.159873413823, 13.4313016634326, 
    13.5460340739175, 13.5154563940814, 13.4067658389308, 13.3970929486191, 
    12.9433781172502, 11.9663787055569, 11.1221732819767, 11.0771468669312, 
    11.3269188554769, 11.3424745475679, 11.0970218932588, 11.1539111990626, 
    11.2365195124116, 10.8791313828917, 10.8273322891031, 10.4769946986881, 
    10.4228448182146, 10.5849062452841, 10.6804586056438, 10.8943508751507, 
    10.7350561988025, 10.664607728498, 10.4692492958592, 10.4092293864193, 
    10.2170782175553, 10.1258178405792, 10.1901198004029, 9.30233580155356, 
    9.26421934072703, 9.76760375494866, 10.0828333548087, 17.7355123840051, 
    17.5322651184604, 17.34812332948, 17.2587816969053, 17.0189893074044, 
    16.9214332320516, 16.5644626751232, 16.2832686851433, 15.828265832998, 
    15.4379156673791, 14.920071082634, 14.7084576016467, 14.582091207906, 
    14.504245534083, 14.3499282922431, 13.7547667234048, 13.1312033733708, 
    12.8845071167934, 12.8509735205054, 13.0987421634762, 13.3572685249993, 
    13.4288962284866, 13.2153350419556, 13.0469625758771, 12.6976983010362, 
    11.9374671552427, 11.1568405266778, 11.1763495783772, 11.575978388336, 
    11.5927444791899, 11.1537160247772, 11.1902138069968, 11.1918433102042, 
    11.152347416116, 10.8878740444983, 10.5426020499504, 10.60358143234, 
    10.6301914917396, 10.8699722497262, 10.7941983192988, 10.4434557414901, 
    10.3878755445601, 10.3496408130222, 10.3645167513706, 10.2656698262247, 
    10.2537846005654, 9.96422821164403, 9.44053968696611, 9.54582513524189, 
    10.0388207185579, 10.1098968691155, 17.5534637179742, 17.5720247016578, 
    17.3773974662243, 17.3877192594114, 17.4027944294186, 17.1426580134969, 
    16.7576930235133, 16.0756925097525, 15.6946002371996, 15.1390278996086, 
    14.7336186124016, 14.69369131712, 14.5482230077851, 14.375931709985, 
    14.1112976514592, 13.4563838370312, 13.0183707434256, 12.7370291744505, 
    12.6355427370276, 12.8035182552294, 13.088113861897, 13.2955764614229, 
    13.1543954788681, 12.9465463903389, 12.6195918570733, 12.2291333245926, 
    11.4544836473002, 11.5348842888414, 11.8879853642633, 11.7625775568193, 
    11.3112167734787, 11.2670102645842, 11.0973931242812, 11.0538146050551, 
    10.917043389964, 10.8203145209576, 10.7948121819124, 10.7071939163725, 
    10.8282976153433, 10.6957312367559, 10.4139380090624, 10.4067263231837, 
    10.4142132595161, 10.4706662823644, 10.4369791425827, 10.3179700719152, 
    9.95600420303565, 9.60936410336476, 10.0670261818676, 10.2305627544226, 
    9.93509572001105, 17.2602429900533, 17.2992574364694, 17.3297518516937, 
    17.4041081591447, 17.4629824023473, 17.4346289262132, 16.6643626003591, 
    16.1254425629397, 15.7088122736745, 14.9951404075846, 14.7437648774536, 
    14.7396598570465, 14.5154233120378, 14.3729744957398, 14.0723978386983, 
    13.4365586479088, 13.0588215996159, 12.8200268926104, 12.7582685781153, 
    12.7425165037307, 12.7935297989952, 12.9453167078606, 13.0725937166165, 
    12.9069238001435, 12.7590567389862, 12.6040681852433, 12.066878156773, 
    12.0456561907661, 12.1811599743021, 11.8295930918669, 11.2917392080792, 
    11.1267851107226, 11.2348059938921, 10.8799042951729, 10.9052579217912, 
    10.8515872064073, 10.7914006824592, 10.6951870271619, 10.8039851961355, 
    10.7188691184311, 10.5853987397391, 10.5304989627346, 10.5715488352416, 
    10.3946444033724, 10.1984609978325, 10.0020841926533, 9.67494343861929, 
    9.69192302625737, 9.9744064340022, 10.0291047027022, 9.69827748726292, 
    17.0137861010058, 17.0614838242115, 17.2424023785023, 17.3753893771627, 
    17.4701983809902, 16.9860497475905, 16.603924767574, 16.1259864709554, 
    15.8228759528799, 15.1010153601815, 14.8451630375806, 14.8580950710534, 
    14.4826676904147, 14.3770136240345, 14.2447972565198, 13.5968123317832, 
    13.1801376735048, 13.0657076609979, 13.0575463015353, 12.7646132005225, 
    12.5880631584292, 12.6114329272978, 12.8660441229554, 12.779503349864, 
    13.0175338499897, 12.990390548944, 12.8360613404142, 11.8743136883675, 
    12.0426298021266, 11.6866636479333, 11.0692722144663, 10.9098049106379, 
    10.8386095911798, 10.8947761481514, 10.7878358906213, 10.4331832614179, 
    10.3112177757178, 10.2833440769909, 10.5162955343901, 10.4439274622892, 
    10.4249378347026, 10.3468755190291, 10.4932928152347, 10.3373717535785, 
    9.98248608945606, 9.53009815630354, 9.27970136283088, 9.57446462780615, 
    9.75007095546634, 9.56834265493055, 9.3069648155516, 16.8540755122753, 
    16.8402933485286, 16.890310607788, 17.0997078904986, 17.2318852887721, 
    17.0841217465833, 16.6184042142029, 16.1571449071788, 15.9382913007831, 
    15.124485838237, 14.8468621794355, 14.755317260417, 14.3953274096318, 
    14.414831925724, 14.5316827321508, 13.9218085401945, 13.4764263158099, 
    13.2416699765966, 13.2276144204812, 13.2248966769448, 12.7165811688806, 
    12.425784314075, 12.6538944814797, 12.8075848844337, 13.0820632707401, 
    13.2154036299875, 12.4801578235493, 11.4137400075858, 11.70422651454, 
    11.5051668755041, 10.8877030780985, 10.6181611336443, 10.5891058489659, 
    10.9062574398776, 10.5837923230519, 10.2465223905273, 10.0657850199759, 
    10.0957586422331, 10.2326002281877, 10.3604219199003, 10.2240744444944, 
    10.1123219069697, 10.1934404055316, 10.0549763685381, 9.5976163256735, 
    9.48440009586515, 9.59421863264887, 9.72092002497149, 9.53772952963689, 
    16.9463179022023, 16.8045647886872, 16.7997335216421, 16.9550359261299, 
    17.0773889308806, 16.8876185342791, 16.5586090193461, 16.2523358601204, 
    15.9308715747076, 15.219668285516, 14.9731744328391, 14.5779767075927, 
    14.4482819923558, 14.5271537282271, 14.5770784550628, 14.0557061738388, 
    13.7298149980279, 13.3847460455364, 13.3428954749992, 13.4094818958987, 
    12.8325269928819, 12.3454462131082, 12.2255852826584, 12.582567079873, 
    13.1008001753526, 13.175490425539, 11.9629131682727, 11.3918907656351, 
    11.594322816236, 11.5318040276947, 10.9642977423235, 10.7278465727336, 
    10.7911317743496, 11.0748464698794, 10.3237510056295, 10.2564202645582, 
    10.2855801419864, 10.3478564899112, 10.4973804614521, 10.322582781443, 
    10.1207018371708, 10.0129974249794, 9.95107640262139, 9.90614071005152, 
    9.77678769402571, 9.92038238128179, 9.76180641113999, 9.78588848359974, 
    9.84656206524829, 9.78847616612594, 9.5280568313334, 16.8472336451186, 
    16.7323476425046, 16.6909747311006, 16.7388624527658, 16.7815095608952, 
    16.6294810067451, 16.6032357967721, 16.350397402086, 15.9820623725349, 
    15.4157034212739, 15.4000958269495, 14.7712657122508, 14.2269487244384, 
    14.3663454932586, 14.4301004149868, 14.1014857745137, 13.8693768389672, 
    13.7121332526363, 13.6986857814676, 13.4566258062363, 13.0644118614625, 
    12.5898119302568, 12.2963932413936, 12.2873856018955, 12.7603185448516, 
    12.95024400176, 11.9000265896419, 11.5804254372678, 11.7977346333943, 
    11.6376169721825, 11.2649282244812, 11.1605958139164, 11.1734478762443, 
    10.9559156713714, 10.4724860059345, 10.5780027521729, 10.163847181461, 
    10.2400795903422, 10.1521414091514, 9.89633151727504, 9.63761998248983, 
    9.50787904632719, 9.67788952633258, 9.66283483727796, 9.36229594625858, 
    9.55040934043489, 9.54258734250874, 9.08752449625896, 16.9828817086667, 
    16.9115026887631, 16.761048571013, 16.6443950305829, 16.5125161726459, 
    16.1435844092578, 16.0393215626031, 16.3226645519385, 16.1698456975052, 
    15.8920820658494, 15.3411851134931, 14.5655888776751, 14.0409586203473, 
    14.0817189621432, 14.1576443013293, 14.0804635859387, 13.9666292893193, 
    13.8660263588878, 13.5543877388871, 13.3208411804632, 13.0978008801453, 
    12.5836299157792, 12.5637411473849, 12.4471809440416, 12.6005529268457, 
    12.5091432112421, 11.7183431066921, 11.6491541607325, 11.8423365625346, 
    11.2084889094456, 11.2413523728137, 11.2469639574457, 10.981470610058, 
    10.3928107855475, 9.40920067896097, 9.75035752041243, 9.5233283788144, 
    9.21599162683033, 9.39664974155399, 9.47366531731928, 8.68207565296107, 
    8.68101714202387, 8.83781885365114, 8.65515999772241, 17.1888641769733, 
    16.9147553609055, 16.7565140854085, 16.5296261354602, 16.3714607617799, 
    16.1105886203982, 16.0546592060723, 16.2377026375454, 16.3175244483307, 
    15.9862490278234, 15.1437701655626, 14.4409599150166, 13.9674528166859, 
    13.8792569553922, 13.8557656820634, 13.8543651119763, 13.8319056808011, 
    13.7125114892447, 13.2262263037526, 13.1339125914847, 13.0091925425684, 
    12.7639093658562, 12.7933017971174, 12.3876099988514, 12.2193470683339, 
    12.0930347020097, 11.716048594166, 11.4389070064906, 8.95545679200173, 
    9.00899702864757, 9.11334224087559, 8.41735145067434, 17.0871614538069, 
    16.8126615687677, 16.6318806390489, 16.4393529056449, 16.3877336319002, 
    16.2020349084592, 16.2190940927515, 16.1568922853358, 15.8558686149142, 
    15.2500105068019, 14.7623658229522, 14.210171207953, 13.9992157204083, 
    14.0410557690349, 13.7045055415254, 13.4294495542572, 13.7390331495572, 
    13.5868893839735, 13.1506090749026, 12.7961348357363, 12.8099341980561, 
    12.6902586238669, 12.536346661825, 12.1782109039611, 11.8871959935944, 
    16.8832255860532, 16.608358855346, 16.5909755257153, 16.4850459420683, 
    16.3880157275521, 16.1737698208118, 15.6372611190867, 15.2053571421236, 
    14.8488073481345, 14.5878471928113, 14.4801383244186, 14.1877588359812, 
    14.2824227930689, 14.3536454852081, 13.9839692589876, 13.309601782832, 
    13.4083701851358, 13.4790207957432, 12.94871532772, 12.7400239880376, 
    12.8507080458189, 12.726811931617, 12.5738625805873, 12.1678654067575, 
    16.8228389098811, 16.5686700461872, 16.6023951951156, 16.3655899132781, 
    16.1322389178623, 15.8315859649247, 15.0555297228812, 14.575698509849, 
    14.3999422787073, 14.297327178897, 14.2844653290748, 14.1558683385227, 
    14.4645389946751, 14.4048925847578, 13.8122090177499, 13.2968204726347, 
    13.4260480477391, 13.4019559624357, 13.273984881852, 13.2603789719238, 
    12.8972183890506, 12.4287094325118, 16.7226865223797, 16.5789696415406, 
    16.6625142155656, 16.0673054174012, 15.8459227631039, 15.3566401322808, 
    14.5969555691546, 14.2772791690164, 14.2942348736448, 14.2246124692158, 
    14.2718675091762, 14.423095286285, 14.3533486991976, 14.1324822796605, 
    13.682000074374, 13.2598340479148, 13.5002259552031, 13.4362744035677, 
    13.2833546868082, 13.0840402828123, 12.8520319687785, 11.9903360716012, 
    16.5501205519504, 16.7240657741488, 16.6390749502858, 16.2203574565103, 
    15.6767148444558, 15.0041671902219, 14.3611974346362, 14.3597527165787, 
    14.4025984495965, 14.3789828686038, 14.372418839695, 14.2783189914636, 
    14.0155316842423, 13.8477492867427, 13.5186147330836, 13.3597481466569, 
    13.4352651969227, 13.1664786422886, 13.0749367594535, 12.8283551883685, 
    16.572038035371, 16.8563720736901, 16.6919436036918, 16.5474131544918, 
    15.9307553120803, 15.2310754661731, 14.6925185457551, 14.5784932271113, 
    14.5275674282103, 14.6344996550505, 14.5432229273957, 14.0243912050785, 
    14.0525737330386, 13.8660241042004, 13.5175354470529, 13.5710304917609, 
    13.4586195678204, 13.240166563745, 13.1265900372375, 16.5172450219906, 
    16.7815628772928, 16.8094910263523, 16.6625096801874, 16.3239641534878, 
    15.653413003731, 15.1864738076245, 14.8140351192561, 14.4254666379979, 
    14.5613749777705, 14.6445262079677, 14.0476370915043, 14.0736725169841, 
    14.0520944496922, 13.7853919711467, 13.5134240328168, 13.443473485265, 
    16.3768327059503, 16.5289376991216, 16.6133651704598, 16.7137820943478, 
    16.9850348735992, 16.4647908945418, 15.8888843328891, 15.0854944139157, 
    14.6047419629701, 14.5417985705729, 14.3256155194621, 14.0903889761779, 
    13.9638199203521, 14.0025747553593, 13.8701945837817, 13.499578585126, 
    16.4049799726103, 16.4385667616755, 16.2808773990585, 16.4635472178462, 
    16.857889511711, 16.721051906749, 16.4388787734755, 15.5867333276357, 
    15.0182089392435, 14.7345098722043, 14.2394545338224, 13.770630735458, 
    13.2922410359133, 13.4469017004959, 13.2210332340716, 16.5391948905696, 
    16.4671025036648, 16.1293451919646, 16.3677040426478, 16.7625919473232, 
    16.6331429135577, 16.4221238155561, 16.0070168654833, 15.4445238708145, 
    14.6212097186539, 13.9487883758227, 13.6285509717434, 13.2351488453162, 
    13.171701434321, 16.7205135071067, 16.5308759817331, 16.081245353571, 
    16.2270786566928, 16.5994782904008, 16.3557484082825, 15.9326018128927, 
    15.9800990555957, 15.3355440060985, 14.4564351767573, 13.919486027593, 
    13.5751064915092, 16.7437366683897, 16.5870673745623, 16.0957944833803, 
    16.073797329405, 16.2099911011722, 16.1865692930266, 15.3451621825532, 
    15.1302938807657, 14.9738300098207, 14.4094115492405, 14.0174115101033, 
    13.9296209430966, 16.6483318404397, 16.5138439515645, 16.0927880772776, 
    15.9653350143179, 15.7884316284524, 15.8994965161988, 15.1941623489535, 
    14.709372063182, 14.8471454352425, 14.1698320930069, 14.0073201292893, 
    13.7892649450444, 16.5621814234444, 16.2939084801695, 15.9409363827527, 
    16.0528352258446, 15.849501709951, 15.6699424079917, 15.3914778386405, 
    14.6549572012055, 14.5774835951189, 14.2041027093458, 14.1251074877391, 
    16.472451929818, 15.949583592439, 15.8678256948725, 15.8840748970989, 
    16.1127657176094, 15.8403765264337, 15.1809282194032, 14.700700845447, 
    14.4761126755916, 14.5460955433228, 14.3795615863479, 16.1778353752983, 
    15.9478977343335, 16.0308279677709, 16.0389248940055, 15.9993642852059, 
    15.6537501661525, 14.8742774932456, 14.8814490135509, 14.6065123392349, 
    14.6276384864567, 14.3747771276027, 16.002950408664, 16.0743790962773, 
    16.133900384502, 16.009296726208, 15.8375131172456, 15.3138110342287, 
    14.9347814965013, 15.1436953037366, 14.8128847232925, 14.5755424153618, 
    15.9493551480765, 15.9115721515649, 16.0424534735098, 16.0761469195518, 
    15.8846920974942, 15.4811051518593, 15.295901652117, 15.5907870746962, 
    15.2340108554743, 16.3481193822365, 16.0151020225034, 15.9977522381192, 
    16.097638440826, 16.0175371222089, 15.7314441929951, 15.4389208285004, 
    15.4980363613501, 15.6540221407543, 16.6944323546645, 16.4945263286039, 
    16.3564190237691, 16.1145290705168, 15.9073971483159, 15.6825300887709, 
    14.9379465606369, 14.2458517865576, 16.6820939377778, 16.7565308332594, 
    16.484145430968, 15.788194936651, 15.317515030127, 16.5426385879913, 
    16.4728910553864, 15.7436571866165, 15.1545350128701, 13.7006228156734, 
    13.715547090697, 13.7612604972007, 13.6330971469287, 10.1265062875853, 
    8.63733547707405, 7.98375815541605, 7.37269986156393, 5.93225557816058, 
    5.19221186312679, 4.56840855304761, 3.96675628749563, 3.42135431721151, 
    3.00437072649328, 2.65198670562551, 2.34948081332731, 2.1393886121908, 
    12.4239525618394, 6.74107942973307, 32.5343868696338, 32.5344244237141, 
    32.5296424967253, 32.5195893502946, 32.8952139376065, 33.5120557042474, 
    33.8698178585661, 34.0222982941287, 34.0970810437007, 34.1948237362654, 
    34.2980477209731, 34.3876538494436, 34.4554869336033, 34.4973957550662, 
    34.5336739329331, 34.5643828712591, 34.5845760070264, 32.5855975566913, 
    34.0588134954031, 12.6607657589389, 12.7086477705858, 12.8295314119109, 
    12.7905311142195, 11.4880408528067, 8.97103350924196, 7.88363591696834, 
    7.35797510501927, 6.95287644028138, 6.3472629602577, 5.39725613082596, 
    4.83029537716885, 4.34837589308301, 3.85326182710722, 3.35806918810827, 
    2.96694214797873, 2.65803168939965, 2.39040975809725, 2.12986126270448, 
    2.00441497461993, 32.4898385949903, 32.4903840895078, 32.494548581556, 
    32.5063876614614, 32.6127292638401, 33.069366792685, 33.6106856452714, 
    33.8618074027999, 33.9546534267837, 33.996159461373, 34.0639572957593, 
    34.1404199641841, 34.251608957752, 34.3659567344986, 34.4530566604771, 
    34.5003687688578, 34.5330097384353, 34.5600746408929, 34.5825908260572, 
    34.5933907051992, 17.7922159928112, 17.7866386499822, 17.8076456147411, 
    17.3791571113, 17.3512749800077, 16.9634097656074, 16.8806434779327, 
    16.6563011553336, 16.6429340308202, 16.4894155207383, 16.4601686184148, 
    16.4564167528663, 16.0754875002294, 15.8732367884389, 15.2780570398155, 
    15.168276762167, 14.7301549140542, 14.529508365959, 14.4186514933546, 
    13.8988344182334, 13.4135088542745, 13.3173835610253, 13.2256655967656, 
    13.4253456068517, 13.6400272585074, 13.6939182621891, 13.6220626950491, 
    13.1289928126393, 12.5949727399291, 12.2317503312608, 12.0820524925694, 
    12.1399103584386, 11.9354896080545, 11.4122008901657, 11.0149202689319, 
    10.8570140018306, 10.583147568907, 10.6990994289464, 10.7928227925911, 
    10.914070521055, 10.7221352732674, 10.6767007816669, 10.6860658691524, 
    10.5677263123084, 10.4676933038803, 10.2584310443917, 9.94098026193457, 
    9.72442153938329, 9.475019209658, 9.32289163886024, 9.12571396622014, 
    17.7240737474109, 17.7280262768921, 17.8070268732075, 17.605684778736, 
    17.1061631195789, 17.1024647420636, 16.7414233468228, 16.7197747070072, 
    16.564863262983, 16.5467555718974, 16.3934224717312, 16.3429671625142, 
    16.1266229145278, 15.9387920210216, 15.4215938954543, 15.1282944757628, 
    14.5769298392657, 14.5825448565444, 14.7379706482434, 14.1627242038394, 
    13.6373676017949, 13.6654820830088, 13.8049007340689, 13.890133025107, 
    13.966529952082, 13.8147688279819, 13.6123053444321, 12.8040785596442, 
    12.4612045026287, 12.3913380448176, 11.9815095535981, 11.9009300019428, 
    11.7654453046945, 11.6347268884841, 11.2211029524861, 11.0121565107587, 
    10.8099304326889, 10.9108497429079, 11.2030313773487, 11.1171473276379, 
    10.8493618607138, 10.7221589938458, 10.720855749875, 10.5717567226892, 
    10.4117235875909, 10.2361316864282, 9.85151548581658, 9.6774719214625, 
    9.51999063273185, 9.48721010848723, 9.38203409220742, 17.6601214724611, 
    17.4991203442403, 17.5299310782637, 17.3530070918565, 17.0151709500742, 
    16.6830802330875, 16.4026061670502, 16.5760384675633, 16.4642151054005, 
    16.5435994451547, 16.3931155309027, 16.4210718834055, 16.2658281826453, 
    15.9713269997812, 15.6457413409457, 15.2856076024406, 14.9612554668767, 
    15.2113570621735, 14.7294798871184, 14.3474284239013, 14.012259390166, 
    13.990990830621, 14.084558568059, 14.0184836598188, 13.899282944499, 
    13.4384904054512, 12.9715003394568, 12.5271090759058, 12.4846914545209, 
    12.3014641990466, 11.9298144409155, 11.8515235315204, 11.8565032826009, 
    11.8775570481657, 11.3868245745812, 11.2672310023047, 11.0746472964315, 
    11.1428384668726, 11.3896509221393, 11.0577196307852, 10.7333412745529, 
    10.7285257785557, 10.597775332924, 10.3293622561876, 10.2127921720271, 
    10.0798441385273, 9.7122790492039, 9.62041374222652, 9.52863519615287, 
    9.70149089742669, 9.57982291932688, 17.7949581532638, 17.4864368571631, 
    17.3610501359095, 17.1756301451218, 16.8496509339677, 16.6608465579921, 
    16.3417134277731, 16.4550765593251, 16.4096464550561, 16.5311738566737, 
    16.3607956589114, 16.309948714746, 16.2236743714341, 15.9524998390801, 
    15.7035074183188, 15.2942951014457, 15.1955514617635, 15.073983501214, 
    14.5120275301272, 14.070112677763, 14.1741864503913, 14.1853360425312, 
    14.1122132295958, 13.9515786917211, 13.7272696403662, 13.1790814020994, 
    12.8594822039915, 12.4120389678872, 12.2074628794793, 11.7475037635951, 
    11.6615150205419, 11.5080138886651, 11.4058995429531, 11.7233012692211, 
    11.4364133364724, 11.3341173097575, 11.1495871600676, 11.325240412028, 
    11.3813174707356, 10.8862825593584, 10.7601194484314, 10.7769140685858, 
    10.3940780669011, 10.0121730808458, 9.85960144700836, 9.60216320738772, 
    9.44308782701937, 9.48848468395324, 9.62419901561178, 9.64816729321852, 
    9.46792430493793, 17.8503929253127, 17.6216961296213, 17.2314398508971, 
    16.9893696935972, 16.7741113324697, 16.6323808246217, 16.4166951041527, 
    16.4212901483133, 16.3902783436352, 16.346753650734, 16.2450458738536, 
    16.2470885089262, 16.1112604689543, 15.8836473854724, 15.7560135987329, 
    15.4484848427544, 15.3674079835996, 14.233718729184, 13.4539742945747, 
    13.2963370603161, 13.5263062363145, 13.7227444374044, 13.7757403366575, 
    13.8678547173556, 13.6711019077913, 13.1617883339947, 12.7129680347125, 
    12.1173384786294, 11.6426628949535, 11.3332604283883, 11.3960069382355, 
    11.2914665562786, 11.1687795874354, 11.3254547672321, 11.2248315328965, 
    11.1462125998902, 10.988743717046, 11.037972636455, 11.1718194121468, 
    10.8468765566289, 10.5309561160603, 10.4173167884685, 10.1188349385074, 
    9.82582620727767, 9.77394730571539, 9.46133642314001, 9.43095581456206, 
    9.60304465764725, 9.57039690519519, 9.54145765447547, 9.48890278585333, 
    17.7562214176451, 17.566707891393, 17.1729359045808, 16.8013001563691, 
    16.7957317249283, 16.5676372016485, 16.2711440601846, 16.2820207512645, 
    16.1824356677694, 16.0400888825489, 16.1486766823571, 16.015207372671, 
    15.9266667514737, 15.7591674845807, 15.7368240614956, 15.4711766667073, 
    14.8209357059251, 13.7217712232111, 13.1180612902632, 13.1582831689469, 
    13.3230403573805, 13.695259254695, 13.655189243617, 13.7489272517157, 
    13.540823829658, 12.857413183043, 12.3945070576655, 11.6386904055377, 
    11.2191803538889, 11.2062164665938, 11.1982613717617, 11.2654221740353, 
    10.9127432719989, 10.9204420424964, 10.853491542536, 10.6898072098132, 
    10.5766143811597, 10.6414260110061, 10.976957429061, 10.7731788242179, 
    10.4432001208271, 10.1651329067879, 9.86578363507191, 9.78363998969436, 
    9.86855795465447, 9.50837333496975, 9.45086170600934, 9.58366278587951, 
    9.4984372696504, 9.45248108106405, 9.34508025800086, 17.732857027667, 
    17.4738048136508, 17.2103185520391, 16.8509945634114, 16.9359905202211, 
    16.6718395593773, 16.4646745945458, 16.2594719509175, 15.9274152419373, 
    15.8826265545743, 15.9915328172495, 15.8970540211483, 15.6754115004972, 
    15.5335898400147, 15.3453882785891, 14.8804003274174, 14.1357751406246, 
    13.2993178940968, 13.0174680180248, 13.1786895693057, 13.2325028665806, 
    13.5536568533788, 13.5253509429898, 13.579743178039, 13.3529866749846, 
    12.5213962063967, 11.8894450961314, 11.0937166338412, 11.2069598367972, 
    11.0749990370754, 11.2071208085161, 11.3432235492928, 10.8590729625769, 
    10.6621797056134, 10.481372758566, 10.5076440896983, 10.5479217833225, 
    10.5514603369053, 10.7511530058119, 10.7814859839195, 10.5995546469798, 
    10.2300267271476, 9.89152161407281, 9.88012595552673, 9.96730216683083, 
    9.6976457433076, 9.41789789088151, 9.46894964700534, 9.34138373842506, 
    9.52388141693109, 9.54200331876241, 17.6790562995943, 17.5958853638475, 
    17.239382138511, 17.1578601879914, 16.8465171901374, 16.7654495757805, 
    16.2479588876801, 16.0561300211654, 15.7176949643053, 15.8259211834026, 
    15.8569623990253, 15.667677665295, 15.5071707810427, 15.425971452968, 
    15.1765622964796, 14.2913943006956, 13.6346406524658, 13.1103176920857, 
    13.1587953736404, 13.3807108862955, 13.4073871695077, 13.4372732809439, 
    13.4000082018009, 13.5406312380813, 13.1400734420367, 12.1807030437012, 
    11.4870389794486, 11.0568897539663, 11.1534274801825, 11.0846879104955, 
    11.0942602425663, 11.2810735268476, 10.8924522617288, 10.3721705737493, 
    10.2451691976248, 10.3646061080425, 10.4503625295462, 10.6873493229791, 
    10.6665961452738, 10.8182535935904, 10.9589254571933, 10.6200254422218, 
    10.2502137619297, 10.1231349667036, 10.0272967384139, 9.92846883289838, 
    9.56069128458489, 9.3190852681669, 9.21753707311922, 9.58715857080374, 
    9.65235418642811, 17.8392682909923, 17.6821750813739, 17.4969898031885, 
    17.1034973963521, 16.7803867002416, 16.4047219603611, 16.301042572808, 
    16.1698460708456, 15.8465912172695, 15.7859787585271, 15.5393407605318, 
    15.1730455467118, 15.1487772132386, 15.3921632181598, 15.3470422196493, 
    14.3206176847759, 13.369943729482, 12.9106950782131, 13.1015412664479, 
    13.3888965312514, 13.5147514852986, 13.4640741760923, 13.465707756572, 
    13.5894375012327, 12.9792136347987, 11.9677226282643, 11.2855471467353, 
    11.0406768314155, 11.1499022013011, 11.164720708231, 11.082987258451, 
    11.1276585476823, 11.0549747934142, 10.4798444420405, 10.2905709653872, 
    10.2679082432951, 10.326610932205, 10.5761373807063, 10.6678263916285, 
    10.8908832358308, 10.9981825635162, 10.6652298607404, 10.328502924047, 
    10.2587138903592, 10.0890648261323, 9.95327975717687, 9.69297610481676, 
    9.20993480312706, 9.06439646115612, 9.74060287325007, 9.92003541545988, 
    17.762298328357, 17.729746667354, 17.5130145461381, 17.2715527962215, 
    16.9411965407506, 16.4593306143115, 16.3185718390863, 16.0025296117998, 
    15.8658557444358, 15.5618779916885, 14.9931576770665, 14.6314425999142, 
    14.6532524329216, 14.8164683225499, 14.8962299288053, 14.0751926473887, 
    13.1182000904713, 12.8400504070963, 12.8934647477701, 13.1953431310709, 
    13.4583757806268, 13.4139386242729, 13.3709272263042, 13.4104399309323, 
    12.8260238339148, 11.8615045498826, 11.104528576467, 10.9584580466968, 
    11.2627572981601, 11.3502307240814, 11.0171354227258, 11.077660013155, 
    11.1830966655384, 10.7442334891551, 10.699618046336, 10.3902797551103, 
    10.3837004454085, 10.5350899776264, 10.6258202568946, 10.8048290311467, 
    10.7172896242264, 10.5488795046136, 10.3530274711354, 10.291267046403, 
    10.1280266087347, 9.98186548718007, 10.0302627901625, 9.14401760065508, 
    9.16677704604115, 9.70338420115101, 9.98466594790315, 17.7256408985636, 
    17.4757401782288, 17.2740343865791, 17.2083983512825, 16.9416212058625, 
    16.8495811916239, 16.5103208521589, 16.374487185164, 15.8509775162753, 
    15.4332475024999, 14.8831594872239, 14.6437604272906, 14.4916988387473, 
    14.376264228832, 14.3184565958825, 13.7247144442808, 12.9814160081861, 
    12.7971729090493, 12.6922942625753, 12.9595286131323, 13.2896958522177, 
    13.3258475929839, 13.1292434269819, 13.0413946247582, 12.6481487175762, 
    11.8473963830174, 11.1421386665472, 11.1869999825675, 11.5552734897699, 
    11.5443148994902, 11.0831487226252, 11.1117113629701, 11.1147557382104, 
    10.9577950713645, 10.7854147735633, 10.4403703801782, 10.6066090103886, 
    10.6040060782007, 10.7939987434161, 10.666938718407, 10.3252329080764, 
    10.2712409820315, 10.2495721972436, 10.236693647831, 10.1482416462049, 
    10.1130611469662, 9.77350818840097, 9.28702013605787, 9.51795744181874, 
    9.91230924338673, 9.94816287550275, 17.4530911316063, 17.5110399636682, 
    17.3582623095451, 17.3291486256141, 17.308631728836, 17.1021874942232, 
    16.7842967346249, 16.1315689726448, 15.7050682588315, 15.1952110520396, 
    14.7254103904639, 14.6427986458589, 14.4975537877232, 14.317405862163, 
    14.0936224345687, 13.4940117458121, 13.0000794889573, 12.7022906433425, 
    12.6322965417604, 12.7976090640915, 13.0508109948458, 13.1938946568796, 
    13.0612738140628, 12.8598050496019, 12.5258911147727, 11.9935622207688, 
    11.3655169539979, 11.5104529533792, 11.8265983409146, 11.6597839035375, 
    11.2496600951728, 11.148681900539, 11.0143831273737, 10.9542515076474, 
    10.8197829272464, 10.7507283486858, 10.7379085026784, 10.6589238514197, 
    10.7591007083378, 10.5557384285802, 10.368188645786, 10.3131504005985, 
    10.3344730854619, 10.3543359364676, 10.2960777002537, 10.1363709439627, 
    9.81045937128619, 9.4495669140739, 9.88038214423191, 10.0395455367394, 
    9.83666770571288, 17.1894907332069, 17.2281824934793, 17.2818828871457, 
    17.3441269917432, 17.385070424116, 17.3808445085002, 16.7193490447535, 
    16.17746617413, 15.6670892510582, 14.9724496654059, 14.6872629702006, 
    14.6880458133056, 14.4862547084029, 14.3466129385626, 14.0588376078266, 
    13.4408904159945, 13.0500939723856, 12.7847699331353, 12.733814421864, 
    12.6774551994373, 12.668274943162, 12.8169057015208, 13.0095421127817, 
    12.8220701262726, 12.6001831583128, 12.3065444340723, 11.9009433324683, 
    11.9667300648111, 12.0695412089517, 11.7305170285435, 11.1744558168433, 
    11.1012760172918, 11.1480305718575, 10.8340768359554, 10.8389558328678, 
    10.7491185708603, 10.6643122103548, 10.6356007374239, 10.7270545425704, 
    10.5955466846887, 10.4600102991917, 10.4793883372802, 10.4226322260679, 
    10.2201667384637, 10.0337592737138, 9.85847469911046, 9.48864443831823, 
    9.56829900636198, 9.76876924513661, 9.87313716885188, 9.5972933827083, 
    16.9675115759922, 17.0233447962311, 17.1813484540736, 17.3113157599805, 
    17.4378629470214, 16.9282124694488, 16.5826754848122, 16.1269516408882, 
    15.7633981337193, 15.0719459369535, 14.8024683902762, 14.8162923734982, 
    14.477068600038, 14.3416810286981, 14.1967016755587, 13.5499674123242, 
    13.1235082669621, 12.9571728358886, 12.9709821553285, 12.7011683516002, 
    12.5075101462417, 12.4776827285077, 12.8182067222609, 12.7577889328513, 
    12.893923532675, 12.7046402564953, 12.6760916655219, 11.8462830096809, 
    11.9643537848992, 11.5834261412051, 10.9515313755156, 10.8565879033651, 
    10.748163141849, 10.8092750862813, 10.7404982272838, 10.3232519410228, 
    10.1985363123387, 10.2190597593112, 10.4979907433247, 10.3879900984758, 
    10.3380586858337, 10.2581121215226, 10.3859049305578, 10.2644424224822, 
    9.88797150992235, 9.43137588394533, 9.14789367717826, 9.50540975868553, 
    9.59620194464017, 9.42031135591519, 9.17151350620672, 16.806904842758, 
    16.8008023323294, 16.8477064553175, 17.0595727732958, 17.1567429464243, 
    17.0479167250812, 16.5771577653115, 16.1365080338882, 15.9450826943559, 
    15.0992573911706, 14.8227499086178, 14.6980162556131, 14.3989864994215, 
    14.4128779885114, 14.498406417503, 13.8309530981135, 13.3512460699167, 
    13.1364361812641, 13.148978826013, 13.1413559972768, 12.6656206312957, 
    12.3437232067868, 12.606838945381, 12.8092205617416, 13.0496680787619, 
    13.0469225009671, 12.4173165990615, 11.3610442022215, 11.6984293878637, 
    11.4248579754241, 10.7716066142784, 10.577904146606, 10.5346924795574, 
    10.8266554381675, 10.5588796328356, 10.2787953342711, 10.0175072033997, 
    10.0528636172581, 10.1579304055497, 10.2846575754729, 10.1641161330509, 
    10.0583708596586, 10.069110570401, 9.92194358976673, 9.46886316395105, 
    9.33005986827716, 9.42928872136948, 9.60907755758914, 9.44666032671027, 
    16.8894576124005, 16.7442504033391, 16.777004118982, 16.9197027807509, 
    16.9806596860438, 16.8029535804731, 16.5312905926659, 16.220030924124, 
    15.9578156581482, 15.1763449076289, 14.9689436528363, 14.5461510439372, 
    14.4238504905827, 14.5556872226283, 14.5560328096353, 13.9195517727371, 
    13.5336751447062, 13.2838305452177, 13.2940728173362, 13.3414980419942, 
    12.7984670441823, 12.324382994846, 12.2497179582087, 12.6172985826818, 
    13.0196477521631, 13.1614408473418, 11.9635156914457, 11.4068360951153, 
    11.5453073216548, 11.4986106073223, 10.8950898241873, 10.7169967242397, 
    10.7831278798212, 11.0236945675447, 10.3820869451878, 10.2205677041145, 
    10.2357958749655, 10.2110230667949, 10.3205829521573, 10.3032609785845, 
    10.0675336776314, 9.93945126191988, 9.82407857054761, 9.78465010037315, 
    9.70923483445131, 9.72463750902998, 9.55992214381411, 9.63317749474339, 
    9.68152269224668, 9.62181249030419, 9.37629403958155, 16.7903991742801, 
    16.7149988533865, 16.6870005094028, 16.7123243651097, 16.6605376011521, 
    16.5157062254154, 16.5707596829568, 16.338997354219, 16.0441140905316, 
    15.4123027024222, 15.3326963865279, 14.7506497800692, 14.1404288498668, 
    14.299663890928, 14.3783534813793, 14.0060925234104, 13.7248410397055, 
    13.5869416544138, 13.5955351436001, 13.395855866594, 13.0365443542615, 
    12.544596463735, 12.2720250346845, 12.2652387924125, 12.681873691385, 
    12.9915164189691, 11.895150461746, 11.5067053694208, 11.7729921626931, 
    11.6595262917086, 11.2560982556252, 11.1486267039523, 11.1472490891386, 
    10.7768186299125, 10.3880728356641, 10.5937274865895, 10.1574045895582, 
    10.2006001545415, 10.223479479809, 9.87575558724442, 9.51722540274616, 
    9.372760549011, 9.48910438075761, 9.50686613705886, 9.09081988772954, 
    9.13931352823098, 9.28613991832716, 8.91162706344379, 16.9435492091307, 
    16.898202019701, 16.7546602208043, 16.618006364641, 16.4233420662841, 
    16.0568670014763, 15.9667348665891, 16.3297458375658, 16.1279817031007, 
    15.815316809531, 15.2876498206544, 14.4137422560289, 13.9377017823941, 
    13.979648669854, 14.0883736200539, 14.0232203108882, 13.9057194582816, 
    13.7805271074751, 13.5257803807702, 13.3143693269375, 13.1283389735768, 
    12.5732828939, 12.5213736039736, 12.4056109097047, 12.532696579491, 
    12.4993605668743, 11.6430154390727, 11.5312146056481, 11.7535848611384, 
    11.1998795435222, 11.2027390440098, 11.1908222694298, 10.9365202901827, 
    10.3495461333691, 9.61474396916552, 9.74223348585847, 9.54766014947524, 
    9.28393453779535, 9.25516776050695, 9.30610622826749, 8.63593119981002, 
    8.44046682508614, 8.65099652634553, 8.42529049175941, 17.1481175893894, 
    16.8679235073395, 16.7571700914176, 16.5430523754554, 16.3540186327367, 
    16.0984116970798, 16.0568539587654, 16.190621218722, 16.2495160906605, 
    15.9256559750718, 15.0850440815478, 14.2788590961607, 13.8475651967, 
    13.8151901610099, 13.7618997684579, 13.7966849279154, 13.9092829963668, 
    13.7315796528297, 13.23318918853, 13.0962305637224, 12.9686768653256, 
    12.7433307449879, 12.7225418070874, 12.3153369212066, 12.1086526805435, 
    12.1350027194151, 11.7919036451407, 11.3836021374541, 9.01734881925945, 
    9.07763307096418, 8.8943967500292, 8.15829580164465, 17.0162756009991, 
    16.7566848598531, 16.6299239356543, 16.4674221906312, 16.3776587095744, 
    16.1720853711837, 16.1664116371183, 16.0631533170466, 15.752031916468, 
    15.1727009882071, 14.7428592077143, 14.1377126711564, 13.9583186049827, 
    14.0538623809239, 13.716897202806, 13.3814321408227, 13.732395621973, 
    13.5482733868741, 13.1554725785494, 12.7469389032598, 12.7634669106629, 
    12.6590275779544, 12.5088276370901, 12.1167466364315, 11.8223945170908, 
    16.8375211669667, 16.5900142762952, 16.5702123919838, 16.4734464662492, 
    16.3213223816848, 16.0010947666557, 15.4508543934514, 15.0436064089527, 
    14.6959956601143, 14.4674358708817, 14.4187300447435, 14.1113840351564, 
    14.2460360734884, 14.3087446517971, 13.9968211245766, 13.2857528560218, 
    13.4157628319721, 13.407315418897, 13.0879433558904, 12.8710681739956, 
    12.8655086098849, 12.7117336014973, 12.5424909618794, 12.1514632869608, 
    16.8265007992396, 16.5866085501046, 16.5905685503608, 16.354400560179, 
    16.0711543591329, 15.6480431321846, 14.8876166864873, 14.4881509846223, 
    14.295855633799, 14.2626847286683, 14.2595602826864, 14.061033821143, 
    14.4138375669075, 14.3408316630765, 13.6764271406015, 13.2328245616653, 
    13.4112026771452, 13.5183067773293, 13.3684004492969, 13.2405108697094, 
    12.7888772593793, 12.4301555642913, 16.767291931114, 16.6155095807025, 
    16.6585401905941, 16.0844967501224, 15.849916420604, 15.3563556264719, 
    14.5806262521076, 14.2490073027535, 14.2748633282015, 14.227283576004, 
    14.2786029863181, 14.3507709529156, 14.260284010167, 14.088924547906, 
    13.6262386308006, 13.2769104706791, 13.4902884058475, 13.303292918478, 
    13.0385635879437, 13.0582968816481, 12.7600309123953, 11.9213300962229, 
    16.6080842138612, 16.7975941925083, 16.691109436095, 16.2101564437184, 
    15.7438445957209, 15.0836681197607, 14.3657270865002, 14.3546270467004, 
    14.395643284094, 14.3933253662055, 14.2919992199104, 14.1278157087682, 
    13.9598979688594, 13.7708564603418, 13.5507209940456, 13.3818011415208, 
    13.3031188629278, 13.0730343546931, 12.9172883634002, 12.8571982007542, 
    16.6442444434345, 16.9273204107718, 16.7527185555385, 16.6513249298166, 
    16.0487949835209, 15.2526735806854, 14.5344601387255, 14.5503788943933, 
    14.4984677249675, 14.5245491309021, 14.3239488770444, 13.8964040809677, 
    14.04899053527, 13.8521088762645, 13.5414909213983, 13.5702661712227, 
    13.3075729429229, 13.2100372384545, 13.0670719010907, 16.5949387378355, 
    16.8815566702605, 16.8988935202323, 16.7868082313276, 16.3631866943834, 
    15.6549555010937, 15.0846926627667, 14.9058996716609, 14.4934579814752, 
    14.4268736706397, 14.4753677030502, 13.9516014805961, 14.0356271744051, 
    14.0150914996395, 13.78441817481, 13.4092271820666, 13.3610035769576, 
    16.4112033636193, 16.5033246422212, 16.5974424852151, 16.7556576068197, 
    17.0025593348725, 16.3962430423776, 15.8495457373094, 15.2635628054325, 
    14.7356708833965, 14.4816501432629, 14.2853136680423, 14.0669366985594, 
    13.8153169543207, 13.8521331335728, 13.6880436633541, 13.5236346461584, 
    16.3784329273269, 16.3286925325342, 16.2160611923723, 16.5161503901994, 
    16.9145492096023, 16.7015434503626, 16.3294109523312, 15.7380085465874, 
    15.1591047838009, 14.7437173340258, 14.2447095511076, 13.7679052955767, 
    13.238380995196, 13.3302561092702, 13.1394576582043, 16.4815239419431, 
    16.3383633932014, 16.0950890642974, 16.3771624956439, 16.7216534168198, 
    16.7310539290177, 16.4479794781606, 15.9938460154559, 15.4626651407131, 
    14.6113784734002, 13.9236725844783, 13.6754367720994, 13.2217066908928, 
    13.0257393769751, 16.6534698927139, 16.4824750610391, 16.079950242518, 
    16.1769566632947, 16.4116925625452, 16.3216455229125, 15.9468714740226, 
    15.8536675500995, 15.2569635186588, 14.4125387223212, 13.8763377882681, 
    13.7023927567103, 16.6575473260022, 16.5721394336872, 16.1527263441163, 
    16.0117933129977, 16.0778034762423, 15.9650505632642, 15.2637828678498, 
    15.0432464689058, 14.99270531, 14.4435294760241, 13.9885018212325, 
    13.8381998652551, 16.5816520786719, 16.5118351065594, 16.1329519630096, 
    15.9304322267722, 15.751059048188, 15.7018409828385, 14.9869944173361, 
    14.6768985348554, 14.7012895146025, 14.1432968198906, 13.9773516051845, 
    13.7054519391805, 16.5360438254864, 16.3785397241938, 15.9969456242669, 
    16.0303136926479, 15.8495840117367, 15.6257076012643, 15.2040143143408, 
    14.6101515649187, 14.5115722895441, 14.1867806136313, 14.0674956582904, 
    16.4573193141582, 16.0392841623874, 15.9304517247142, 15.8909765668782, 
    16.1826494925707, 15.8180248997346, 15.1256852772127, 14.7165821021107, 
    14.4952834493819, 14.5258833347634, 14.3525935716917, 16.1867934826174, 
    16.009429053446, 16.101170090541, 16.1915347925992, 16.0858357903579, 
    15.5994192021119, 14.8191167528697, 14.8673716776678, 14.6486576467081, 
    14.5446733737803, 14.3505917607762, 15.9815284033073, 16.0979228207016, 
    16.1699657992341, 16.1036889405257, 15.8681973057073, 15.2678766401067, 
    14.9606113492894, 15.1745748147871, 14.8091685353066, 14.565947524675, 
    15.9118247586609, 15.9335923009642, 16.0907001428372, 16.1172929154977, 
    15.8683327323559, 15.4562894950867, 15.3485776066496, 15.6059446737079, 
    15.2431828528857, 16.331050948442, 16.0244153133195, 16.0543566486741, 
    16.1140188506751, 15.9732029906355, 15.6379676129308, 15.4047684450694, 
    15.5556818234391, 15.8288105608416, 16.6739091564084, 16.5196202431446, 
    16.3620061691642, 16.0921332185363, 15.7690582319, 15.5133945203921, 
    15.0127675410944, 14.2743976809896, 16.6557538623894, 16.7403387347425, 
    16.4360922488567, 15.7424601219352, 15.234563483756, 16.4559992638103, 
    16.3512561720436, 15.6957950433081, 15.1473380538183, 13.9314239003044, 
    13.9772717828893, 14.0525021269893, 13.8887059035234, 13.3899626395848, 
    12.470138956786, 10.6835183489039, 9.41393661693309, 8.96365022038104, 
    8.53536303700088, 7.90515534592795, 7.235459173857, 6.71475948447939, 
    6.2693228686202, 5.90224366647207, 5.49634410603202, 5.27184303638464, 
    5.08520529479343, 4.80509617452574, 4.5114714040698, 4.34841122736352, 
    4.20036028853035, 4.07025738513598, 32.9879621079745, 32.9917654703942, 
    33.00661468271, 33.0228758110023, 33.0487616814404, 33.1509410844952, 
    33.4317615419256, 33.6824001125732, 33.8956016707641, 34.0173192401012, 
    34.0748923606437, 34.1149753274659, 34.1442686676377, 34.2110696721405, 
    34.2464143215164, 34.3043592010291, 34.3396598694583, 34.353280729434, 
    34.3784131718746, 34.4104711405873, 34.4216495958861, 34.4299067856121, 
    34.4379829404317, 12.2894951932145, 12.2974340886813, 12.2594531772786, 
    12.1772476390268, 12.0232541865317, 11.2098928238206, 8.97732825476131, 
    7.88256562459444, 7.60772868814629, 6.97239558831644, 6.1470836231413, 
    5.27054302360717, 4.71433366850667, 4.29066888851302, 3.83925937804262, 
    3.43128593522438, 3.09611844071284, 2.81011683272489, 2.56134138955988, 
    2.33726958776347, 2.17316163821943, 2.03409513479534, 1.93882934833345, 
    32.6017822479058, 32.593070762605, 32.5735066953329, 32.561532423086, 
    32.5540811702726, 32.5722314640953, 32.8744887095852, 33.4106634333765, 
    33.7084131609023, 33.9326896425578, 34.0121677827589, 34.0317002536811, 
    34.1057159008559, 34.1777043582802, 34.2733707752952, 34.3665810988481, 
    34.4283165836742, 34.47175096358, 34.5069257906995, 34.5382918233012, 
    34.5612382612836, 34.5800965428949, 34.5924868906942, 8.10105603008503, 
    7.49381828942148, 6.52432346185931, 9.93082110123008, 9.94530114150129, 
    10.0695777065435, 10.3855530617107, 10.358717578892, 9.60283693203118, 
    8.47366797045026, 8.20257949629574, 7.74164956867014, 7.11002835651068, 
    6.19446471524929, 5.95850741402643, 5.80439040861563, 17.7298976556585, 
    17.7450376313607, 17.7342974071271, 17.2609229946714, 17.2814574292731, 
    16.915374326026, 16.8309445180792, 16.633473637732, 16.5917313823001, 
    16.4665141853151, 16.4589484802956, 16.4316064816343, 16.0679428037977, 
    15.8140260707041, 15.204797536084, 15.13569156895, 14.6973104426085, 
    14.5249053968178, 14.3394223726352, 13.9029802617663, 13.5119789673959, 
    13.3031522393443, 13.1190925239674, 13.2789395337287, 13.6506748267934, 
    13.7398011847849, 13.6018104108255, 13.0742797889604, 12.5864154389389, 
    12.1659454923659, 12.0914841859133, 12.1739042115227, 11.873205763272, 
    11.3148837191224, 10.9824984337096, 10.8080957232274, 10.5000494958261, 
    10.6318783005841, 10.7833852917404, 10.8695605362333, 10.6819874804726, 
    10.6373893404728, 10.6208592419199, 10.4944747255318, 10.4128964725304, 
    10.2080895615181, 9.85121399515498, 9.65672053605814, 9.42561193679781, 
    9.25272571150525, 9.06917529367305, 17.6507850323835, 17.6905456481143, 
    17.7526082355275, 17.5069148412651, 17.0859371169861, 17.0745505272319, 
    16.7080988602586, 16.6885583965033, 16.5105104153375, 16.5392543266253, 
    16.3550814302087, 16.3260694080016, 16.0654892371594, 15.8813300067178, 
    15.3452457882467, 15.08551009489, 14.5429567648375, 14.5797136924519, 
    14.7287664470925, 14.1811529747062, 13.6256697097123, 13.6201581627141, 
    13.6770199949632, 13.816077397981, 13.9582493629167, 13.7345820795642, 
    13.6175528862884, 12.787937500943, 12.3683021345591, 12.2100569140499, 
    11.9026604689591, 11.9085777457076, 11.7311624768824, 11.5231275118861, 
    11.1172100101814, 10.9103271892505, 10.6873182297984, 10.8138382546171, 
    11.1499110357193, 11.1164695911416, 10.8797404616857, 10.693108267206, 
    10.6193062490305, 10.475217901136, 10.2991249174629, 10.1228320367444, 
    9.75167531848291, 9.61024368449707, 9.4644834806659, 9.38846862786576, 
    9.20657400483435, 17.5919250797271, 17.4518774671936, 17.4801620708077, 
    17.3312551866912, 16.9877896145985, 16.6878660307789, 16.4014222779895, 
    16.5495760114868, 16.4271416117326, 16.5113388926583, 16.3517989802954, 
    16.3871932398234, 16.1936160936658, 15.940993166286, 15.5730691682188, 
    15.271359138945, 14.8920968677399, 15.1906041183259, 14.7079741430556, 
    14.3945440394521, 14.0023440128263, 13.993296112397, 14.0190443882684, 
    13.9882010166799, 13.8800920083243, 13.3305891512811, 12.9818713940814, 
    12.5214359204987, 12.3807430353671, 12.1458478660024, 11.8780978845567, 
    11.8499945142839, 11.8130290694931, 11.7944323126558, 11.3112796547917, 
    11.1568033890094, 10.983075045538, 11.0344167592132, 11.2997856486501, 
    11.0196983564549, 10.6996916670424, 10.6468141700481, 10.5195328947216, 
    10.2159046294349, 10.0435428371751, 9.90643068295394, 9.61709080166908, 
    9.55421677774797, 9.48767021298571, 9.61967143085849, 9.48225946929763, 
    17.7209056078496, 17.4257201168245, 17.3229718284293, 17.140605766684, 
    16.7887943566188, 16.5621182562249, 16.3715177523853, 16.4257043312614, 
    16.3952880444339, 16.522985839878, 16.3152540458171, 16.2823593059695, 
    16.2102482880047, 15.9557487662487, 15.6708977220956, 15.315170750221, 
    15.1532306362984, 14.993841718308, 14.4116685172725, 14.0994415309864, 
    14.1306409552851, 14.205811671212, 14.1427220409356, 14.0306183881561, 
    13.6976581589569, 13.0930337964791, 12.7880030211951, 12.3387558299353, 
    12.0209652336024, 11.594778319909, 11.6596689224633, 11.5617838767485, 
    11.3751557659072, 11.6861268634048, 11.3949773965049, 11.2863570187409, 
    11.1141696345513, 11.263802589384, 11.3354135703731, 10.8383422757984, 
    10.6923278798464, 10.6484824585106, 10.2814686133331, 9.86064741427961, 
    9.6937818929073, 9.47282040054163, 9.36014493311948, 9.40516983966826, 
    9.51730680178261, 9.51665544339887, 9.35918613111984, 17.7798000316343, 
    17.554070235171, 17.188297739037, 16.9819146965005, 16.7474340280076, 
    16.5949847678298, 16.4190083687017, 16.4321977969361, 16.3699657906049, 
    16.2933779104497, 16.2183005743449, 16.2310437801796, 16.115571916492, 
    15.8902111406666, 15.7167964364924, 15.4331612025209, 15.2714400116085, 
    14.1548050378979, 13.3591360348009, 13.256824419392, 13.5081118211672, 
    13.6982618146324, 13.7736943119606, 13.8656961374161, 13.6264020693276, 
    13.0675548668475, 12.6421066052974, 12.0319085024124, 11.4985722601066, 
    11.2640199352407, 11.3548934603626, 11.296570300434, 11.1886651114577, 
    11.3424101791258, 11.2067943435275, 11.1064783790157, 10.9471506878459, 
    10.9791662790176, 11.1274591682104, 10.7887486363152, 10.4407214680279, 
    10.3620007895182, 10.0762772778701, 9.72502715319778, 9.66994674215439, 
    9.36977594481555, 9.390269741162, 9.54843413572157, 9.43205821180191, 
    9.45612785425076, 9.39891285592136, 17.7058923301795, 17.5354057210574, 
    17.1464951766726, 16.8300242241726, 16.7860965609314, 16.6045154826351, 
    16.3121555034201, 16.3182401547484, 16.2012334612657, 16.0252714309812, 
    16.1278777156431, 15.9738703509245, 15.9658094322669, 15.7782715745161, 
    15.7424587943842, 15.5215170647656, 14.8925419557786, 13.6743468244281, 
    13.0761526896552, 13.2006096716044, 13.2857272370539, 13.6418589981435, 
    13.634473130267, 13.7384000608786, 13.4451975367572, 12.8027194251178, 
    12.3877750836728, 11.6518981848147, 11.1323344564358, 11.1451831783662, 
    11.159039540986, 11.2038307478382, 10.9131482667836, 10.9444571017292, 
    10.8083735931805, 10.6298201103396, 10.5477668009512, 10.5866046163116, 
    10.9447729152705, 10.7224164943944, 10.3454001592492, 10.0835107001199, 
    9.85204719848373, 9.71835600391491, 9.77953068931278, 9.42568412387703, 
    9.37525403450063, 9.50129173350368, 9.35037574440734, 9.33992801995396, 
    9.28984329384083, 17.6653046863352, 17.4166936940544, 17.1614294636246, 
    16.8133917528209, 16.934700720948, 16.6961635677543, 16.5415587838153, 
    16.3095386569182, 15.9407834894735, 15.9120061523441, 15.991733506016, 
    15.8733045442629, 15.696398928193, 15.5699258440456, 15.3765349377864, 
    14.8828553888944, 14.1120894877449, 13.2460253126726, 13.030656057569, 
    13.2696794957411, 13.2774905641736, 13.4437517073075, 13.5104397032859, 
    13.5538240833359, 13.2274880413707, 12.4653105119632, 11.9040441000289, 
    11.0798368313016, 11.1585808391004, 11.0327239818538, 11.1631423862507, 
    11.2638928148132, 10.7970718394629, 10.6653464873427, 10.4675828727508, 
    10.4764983575523, 10.528584457664, 10.5326579594909, 10.7301508873035, 
    10.7413846654453, 10.5128769322245, 10.1370464323789, 9.81109998361216, 
    9.77845495401785, 9.88492226089194, 9.64009320877854, 9.34716730595696, 
    9.35995160115422, 9.23322156466826, 9.40605389563169, 9.33849551584814, 
    17.6430412093003, 17.5035209744624, 17.1763215428927, 17.1156693508771, 
    16.8676719273519, 16.8329856916132, 16.3363983570629, 16.1413769321887, 
    15.7648226887402, 15.877030299115, 15.7930733030322, 15.5986123231243, 
    15.5001700912351, 15.405521340661, 15.0729423636332, 14.2283035011204, 
    13.6131853440278, 13.0813158066138, 13.1213726414805, 13.3324970857769, 
    13.4534783771163, 13.3841012209637, 13.3540332496295, 13.4457227119532, 
    12.9484051601537, 12.0711855079192, 11.4613004590246, 10.954764764724, 
    11.0848327727795, 11.0646232393616, 11.059665899944, 11.2364286011382, 
    10.8372403248107, 10.4063204337286, 10.2389564470242, 10.3349112819115, 
    10.405274435376, 10.6389800052452, 10.6540900555617, 10.751870858962, 
    10.8959956110287, 10.5600971925712, 10.1620052754413, 10.0293123308655, 
    9.94952013209441, 9.86121136729935, 9.52240358229905, 9.24246521013122, 
    9.19500867298943, 9.55141846200236, 9.5611729112073, 17.7535732339772, 
    17.6597566329635, 17.4705247725167, 17.1259387593772, 16.8022360102604, 
    16.5261917787388, 16.3807909657824, 16.3136052476653, 15.8811708365725, 
    15.7709326564877, 15.4291857957896, 15.0942440138648, 15.1580250578342, 
    15.3897719391743, 15.295472468518, 14.3386332712354, 13.4715875043116, 
    12.9639066256996, 12.944229643216, 13.2411373025731, 13.4799340803062, 
    13.4102703514924, 13.4020653882391, 13.4899650800547, 12.8095531907634, 
    11.8464524031876, 11.2679847403172, 10.9232159877368, 11.099834811676, 
    11.162203005401, 11.0646053298486, 11.1329264022937, 11.0277052121996, 
    10.5114553550725, 10.259709756482, 10.2176022601204, 10.3310771042702, 
    10.5244777119086, 10.6448103390066, 10.8220082275846, 10.9488694376985, 
    10.6644690927923, 10.3048392993579, 10.1973028591192, 10.0443241875379, 
    9.88485031979079, 9.62897177502944, 9.12614586323947, 9.07432753954292, 
    9.67575404862328, 9.81273408398187, 17.7639776615665, 17.6206516558014, 
    17.5102957134137, 17.278693395729, 17.0001712608989, 16.4796138277773, 
    16.393732445414, 16.0906358617398, 15.9415765340805, 15.5031425826871, 
    14.8978113268739, 14.5870783318496, 14.6639506632386, 14.8511451018777, 
    15.00194135752, 14.1491830655595, 13.2577003726826, 12.8638100899422, 
    12.7754946787052, 13.0876397180784, 13.4072492718173, 13.3683112525841, 
    13.3684412585862, 13.4183718724488, 12.7614099939542, 11.7665496735521, 
    11.1628874866526, 10.9260542547377, 11.2471418025186, 11.3647133541599, 
    11.0010076887822, 11.0866626747989, 11.1623575580472, 10.6909138177387, 
    10.6326406390759, 10.3860904374963, 10.4450222128224, 10.5148099744085, 
    10.6073806111548, 10.7680942995713, 10.7089107162645, 10.5395948776011, 
    10.3367173869914, 10.252679983757, 10.1050808144305, 9.90862803242369, 
    9.92457371033909, 9.0316924655307, 9.06191606403106, 9.59785684072389, 
    9.88900025486444, 17.739302580331, 17.4122364045752, 17.202694933374, 
    17.1781214249781, 16.9275154049792, 16.8015455734509, 16.5127300619629, 
    16.5086502081155, 15.9483358994711, 15.4590369822088, 14.8778420379787, 
    14.6198537783804, 14.4482598038558, 14.3452688469398, 14.3765490511313, 
    13.7430070735257, 12.9933675331525, 12.8202570896962, 12.7047949509485, 
    12.9804318221785, 13.2750627756217, 13.2623595310492, 13.119450809205, 
    13.097990404462, 12.6564821986999, 11.8137144126735, 11.1373553010821, 
    11.1696687224762, 11.5211574067141, 11.51862568081, 11.0625746412712, 
    11.0765303630908, 11.0747108122426, 10.8434712736919, 10.7651818616262, 
    10.4283379464031, 10.6222760347446, 10.6124998943916, 10.752278192017, 
    10.600759249016, 10.3030961775088, 10.2481483336925, 10.2200947682006, 
    10.1743831477854, 10.0717485888896, 9.99321624029428, 9.67197709835639, 
    9.1239386964738, 9.42260544439338, 9.76832425522312, 9.85097002279281, 
    17.3119609381725, 17.4106604487639, 17.3144004099482, 17.2454793924188, 
    17.223401292816, 17.0485880579384, 16.8363302982085, 16.2925526774788, 
    15.7851105135382, 15.2945153100909, 14.7926039106121, 14.6535896050062, 
    14.521984866451, 14.337271377138, 14.0964645643325, 13.5422345644982, 
    12.9697919055333, 12.7267794434627, 12.7125635991354, 12.8558924785261, 
    13.0401081191017, 13.1430339078802, 13.0057600482232, 12.8469367414251, 
    12.5157117230011, 11.910785415183, 11.3075908123921, 11.474206380367, 
    11.8168483118824, 11.6378013100121, 11.2066959682852, 11.1114618807882, 
    11.0132627475351, 10.9443526549827, 10.8357462867327, 10.7535941294796, 
    10.7160398739456, 10.6553599978356, 10.7102275043247, 10.5015338040832, 
    10.3548465936654, 10.2635005640582, 10.2965598618033, 10.2920766869944, 
    10.2075312929421, 10.0209551352522, 9.6847153713591, 9.29729146722892, 
    9.73314843936794, 9.91795343889381, 9.73669553232637, 17.0719867502621, 
    17.1227830661488, 17.1958081100908, 17.2629675226087, 17.2970637065433, 
    17.3398571963287, 16.8155223423016, 16.2494856977406, 15.6623598212971, 
    15.0372325896811, 14.7147764039433, 14.6817313680533, 14.5290014918107, 
    14.4053777286548, 14.0885794730824, 13.5326176139797, 13.0923185989409, 
    12.8437107840192, 12.7485984474682, 12.6524602880081, 12.6276629070917, 
    12.796441562054, 12.9958249036565, 12.7888267784844, 12.5083864338456, 
    12.0956442192887, 11.7453703441097, 11.8996736890331, 12.0032759792646, 
    11.691435505625, 11.1490136980255, 11.1210461619164, 11.1056357518041, 
    10.8665219573685, 10.8012356708649, 10.6979819718357, 10.6417038812486, 
    10.5987714342225, 10.6778214287951, 10.535391405004, 10.4229880556118, 
    10.4501190354314, 10.3684190832353, 10.1419863560226, 9.96962505890763, 
    9.76469725768235, 9.37691359714353, 9.45099123196783, 9.66002384091812, 
    9.73687964264807, 9.56276584497969, 16.8744015306147, 16.9592155858188, 
    17.0908969222808, 17.2262104931544, 17.3911092285315, 16.90433244513, 
    16.6070107919392, 16.1410439351247, 15.6947311435076, 15.0768728915266, 
    14.791821490757, 14.7893924632608, 14.519395561416, 14.3650552117944, 
    14.2081537336776, 13.5877959326209, 13.172812175504, 12.9379240911681, 
    12.9306104902973, 12.7294543765674, 12.5120692563643, 12.4644375393735, 
    12.8302018546814, 12.7620367826897, 12.8119366541885, 12.4372395976621, 
    12.557924085903, 11.9023047442099, 11.9371512852846, 11.5957558704387, 
    10.9288991061601, 10.9602570082332, 10.7869864911178, 10.8081052710171, 
    10.7932999810819, 10.4197681496391, 10.1707122509892, 10.539333591709, 
    10.3808438708674, 10.3431104403098, 10.216162175707, 10.3587740428695, 
    10.2727248053334, 9.88062530744449, 9.40069897734198, 9.10717101566301, 
    9.3823798898379, 9.50024133188451, 9.36318625078106, 9.20303797812396, 
    16.7222931227551, 16.723212410006, 16.7852999182643, 16.9919863581564, 
    17.0759448367957, 16.9972942459155, 16.5540405871425, 16.1128309465936, 
    15.939082246072, 15.1105752001557, 14.8353311011202, 14.6631005499501, 
    14.399077258435, 14.4066255465559, 14.4757841692024, 13.7847196154948, 
    13.2880780730386, 13.1056415164479, 13.1209061197351, 13.15320039119, 
    12.722045939568, 12.3614009014969, 12.6406940963218, 12.8485634144158, 
    13.0299124273769, 12.8532947524247, 12.4494387162118, 11.365189298301, 
    11.7159448683099, 11.4415855970065, 10.7775952835533, 10.680921852954, 
    10.5482404250214, 10.7573867129568, 10.6380898012071, 10.4022145824813, 
    10.075864246937, 10.0968735049031, 10.1893128151758, 10.3400958392756, 
    10.2385275529797, 10.0053443108098, 10.1178000785481, 9.9274584517041, 
    9.48037530892371, 9.30890560410342, 9.31007529914018, 9.5095819434059, 
    9.42346796300848, 16.7962500092037, 16.6502681952604, 16.7367505157964, 
    16.8566050386983, 16.8730342714194, 16.7056768084253, 16.5086086959348, 
    16.1823746782489, 16.0008106264336, 15.2040764315012, 14.9831516000393, 
    14.5425620025803, 14.3771611488631, 14.5020650303396, 14.5106867299349, 
    13.8211589449014, 13.3967782283177, 13.2191198285103, 13.2911311488714, 
    13.3157110376888, 12.817149657122, 12.3701668428558, 12.2843633777788, 
    12.655204322385, 13.0032416531669, 13.1376547837245, 12.026342329381, 
    11.3998609007847, 11.5302505409232, 11.5120130753295, 10.9154052783479, 
    10.7540145401293, 10.7589900055819, 10.9610506129538, 10.5706991008963, 
    10.3256789277163, 10.2384298026556, 10.1705808442179, 10.2785690341178, 
    10.2637514649416, 10.0980853178396, 9.92327175902595, 9.8176649948473, 
    9.84684903646662, 9.7466680324747, 9.6585845935724, 9.50876481495253, 
    9.51817329169424, 9.65677501531846, 9.606260679359, 9.47762412152912, 
    16.6888689861578, 16.6584107105936, 16.6389921884976, 16.6619475328875, 
    16.5197717260432, 16.3975175854968, 16.5472207583188, 16.3119602948044, 
    16.1194065353932, 15.4645994752986, 15.2985732340155, 14.7260541163123, 
    14.0989696089108, 14.2492046837833, 14.3384797651886, 13.8836984142237, 
    13.5732949480654, 13.4817800961764, 13.5715109262582, 13.3991584329831, 
    13.0792968767775, 12.581249874611, 12.3229705700696, 12.3254382094964, 
    12.7028433514085, 13.0900768178819, 11.942813158486, 11.5077162259718, 
    11.7150154703396, 11.6743082247506, 11.3095740319448, 11.1689892567726, 
    11.1847336417793, 10.7846598162094, 10.5833960668177, 10.1382272486614, 
    10.1608036762216, 10.2501578712436, 9.91746470847698, 9.63766965015755, 
    9.4838420045481, 9.41367003922273, 9.42954097478458, 9.02243190931967, 
    9.01138817256543, 9.28997727134361, 9.0238201427124, 16.8367094081787, 
    16.8264464488478, 16.7298814709926, 16.5634619350361, 16.3322809088107, 
    15.9873588603528, 15.9152722074539, 16.3310500110351, 16.1409645398588, 
    15.7789250960849, 15.2493113590222, 14.3774565634711, 13.9042323073614, 
    13.9671236187938, 14.0605739361046, 13.967359371494, 13.853068970863, 
    13.7401792022258, 13.5593780377057, 13.3490571133304, 13.1518519295195, 
    12.6133446384894, 12.5391957139112, 12.420964713742, 12.5362217865609, 
    12.6204112004844, 11.7252470850082, 11.506217155372, 11.6941592334352, 
    11.256159532023, 11.2242630395934, 11.2042225840412, 10.3554245302006, 
    9.73533903287284, 9.67771827566801, 9.39062320530706, 9.15960770738828, 
    9.15467844664684, 8.6498045844547, 8.44632433512629, 8.62004278930976, 
    8.41109249042045, 17.0336774701559, 16.7633163443109, 16.7486581265837, 
    16.552622803012, 16.355211330356, 16.099861993764, 16.0775472344021, 
    16.1654672940514, 16.207508332265, 15.9054041737929, 15.0497012111809, 
    14.1936570600443, 13.8189917588527, 13.8165965582486, 13.7048939678813, 
    13.7742172287921, 13.9568778299248, 13.7841577148293, 13.2459681047052, 
    13.0535821812936, 12.9691566897704, 12.7631944341836, 12.7142104496653, 
    12.2435375184359, 12.0963836448508, 12.2377422004876, 11.8581435873322, 
    11.4292645588732, 8.99219720911922, 8.99858794771387, 8.75779556864861, 
    8.08608070118188, 16.900875007509, 16.6533126091995, 16.570614898088, 
    16.4648553632952, 16.3674958472046, 16.142357324163, 16.1236046110429, 
    16.0038583291167, 15.6905345843901, 15.1426966208964, 14.7449962459703, 
    14.1017732164124, 13.9698796551323, 14.1027177468, 13.7445557428601, 
    13.3654119227894, 13.7230114282204, 13.515620480584, 13.154197336485, 
    12.7725561375173, 12.7641940385394, 12.6354743279722, 12.5073366180497, 
    12.1412554990349, 11.8249378832217, 16.7687542054868, 16.5646808288836, 
    16.5214613116933, 16.3968939119674, 16.197573493712, 15.8560065316337, 
    15.3590844892828, 14.9301208402791, 14.5538678750734, 14.362288347129, 
    14.3931716453205, 14.0737663583991, 14.2180969424831, 14.2825983631003, 
    13.9917129229491, 13.2775823134605, 13.4118766694223, 13.4383324579742, 
    13.236787608257, 13.0253039744209, 12.9264857274078, 12.723488742273, 
    12.5086664164875, 12.1313995717955, 16.7736773576593, 16.5733815536891, 
    16.5325617222905, 16.267170110205, 15.9332569762201, 15.4092369494859, 
    14.7425979002993, 14.3830162630335, 14.2088381551194, 14.2007478866072, 
    14.2216871149128, 13.9843909777639, 14.3881981202682, 14.2798923734523, 
    13.604813999389, 13.2328984798181, 13.4057781255146, 13.5088275039883, 
    13.3197404405869, 13.1687769045294, 12.8317739972457, 12.4606885159803, 
    16.7313444488296, 16.6156569014532, 16.5997509549977, 16.0424689328798, 
    15.7627840888967, 15.225740192023, 14.4881211254648, 14.1992792064755, 
    14.248257119202, 14.2387004086988, 14.2761714444502, 14.3137908800669, 
    14.2264620931089, 14.0557375178174, 13.6153979037339, 13.3273017075586, 
    13.4605964567524, 13.3633235047189, 13.0605826866302, 12.9660691770725, 
    12.5824929751795, 11.8884386375379, 16.5921851571372, 16.7859245875932, 
    16.6686113651673, 16.1313376165766, 15.6784178486285, 15.0839094181887, 
    14.3533198486631, 14.317528520698, 14.3746705097328, 14.3727951113413, 
    14.2094829731723, 14.0576284671597, 13.9777328373987, 13.7511364962039, 
    13.5378330272055, 13.4155308973868, 13.2841938699403, 13.1432642995586, 
    12.9876796025548, 13.0799103420795, 16.6286189985179, 16.8918503526808, 
    16.7312889008338, 16.6127676245103, 16.0310157455298, 15.2561968093077, 
    14.4296304274073, 14.4469107794062, 14.444098020091, 14.4096226638974, 
    14.2292488925486, 13.8878790516944, 14.0439145576439, 13.7936257654234, 
    13.5804637336609, 13.5009397408989, 13.3397783877955, 13.2501493921521, 
    13.0744944487853, 16.5934184854759, 16.8220323696243, 16.8142870944001, 
    16.7682317449692, 16.3272303153569, 15.5522722530701, 14.8620877383682, 
    14.8583491921635, 14.5458202509327, 14.3405221632348, 14.3891821968488, 
    13.9388597831952, 13.9936681469663, 13.9919734713166, 13.7866668724691, 
    13.4732165056786, 13.3770607340026, 16.3938636982848, 16.3735624576478, 
    16.4120472576792, 16.6278807347487, 16.8713866085595, 16.200012645654, 
    15.6458383225232, 15.3232739986845, 14.9144582444357, 14.5602377686295, 
    14.2558898534106, 14.0461599202698, 13.765091680533, 13.7753403682623, 
    13.6279835441575, 13.5471225987277, 16.2870252730609, 16.1860081717316, 
    16.1025007314673, 16.4287434727367, 16.849551159736, 16.5299251930791, 
    16.180001214832, 15.8431677420841, 15.3389807775489, 14.8106034337235, 
    14.2230494100394, 13.7100331525704, 13.1837248535355, 13.2081903474137, 
    13.0886277650247, 16.3810320721585, 16.2308633606052, 16.0212627607807, 
    16.2604648791012, 16.5991146997378, 16.7189926232467, 16.4332477120839, 
    16.0382859090136, 15.537630837393, 14.6254153608361, 13.8707126714608, 
    13.6496539293927, 13.2050955788799, 12.9711010982947, 16.563216205125, 
    16.4415853644616, 16.0733155320805, 16.0522636916083, 16.2734152597628, 
    16.4113986778958, 16.1211658436529, 15.840676233156, 15.2369907182923, 
    14.3901717567154, 13.839637988359, 13.6795258807668, 16.5722099036445, 
    16.5349209653281, 16.1639598572271, 15.9103446342356, 15.9346293431135, 
    15.9035078997335, 15.3545140029915, 15.0657271724707, 14.9535462229777, 
    14.4969818357072, 14.0092200805143, 13.8201772028842, 16.5133965800447, 
    16.4513966309634, 16.0988391290709, 15.8603003841919, 15.6696291574036, 
    15.5357556891543, 14.8827062115254, 14.6698950604118, 14.6317174793075, 
    14.1956953253985, 14.0198100681107, 13.7444853325713, 16.4699758052279, 
    16.298090588564, 15.9730230145441, 15.934020470502, 15.787496451783, 
    15.5124990562265, 15.0330908294155, 14.5655472784131, 14.4752072672315, 
    14.1519749941288, 14.0531886740312, 16.4105688715629, 16.0395165338065, 
    15.9143312760292, 15.8660854894141, 16.1074159349959, 15.7320029270019, 
    15.0920184524297, 14.7040062237269, 14.5206008873781, 14.4431840435598, 
    14.2590665120337, 16.1898248884171, 15.993881661884, 16.0933276700036, 
    16.2058309808358, 16.0150978577138, 15.4903645983658, 14.8341862294588, 
    14.8622590136382, 14.6693631064508, 14.4982492921665, 14.4141196292317, 
    15.9421331977995, 16.095803514361, 16.1723630154676, 16.0703666153485, 
    15.7459998806134, 15.1884095069584, 15.0067370735934, 15.1379566389222, 
    14.8003465924156, 14.668648934744, 15.8521479438295, 15.9477638001672, 
    16.1030016297691, 16.0574604977157, 15.8011121631572, 15.4586550528668, 
    15.4380474381181, 15.6535697085813, 15.2743487490177, 16.2586612271451, 
    16.0184602362949, 16.0764604044309, 16.1046030794601, 15.8931469729226, 
    15.5987806606519, 15.4823959079932, 15.646301330583, 15.9232695057882, 
    16.6797984393609, 16.5418058134134, 16.3906523410586, 16.0469979780323, 
    15.5393161685255, 15.3891534595422, 15.3103476858768, 14.6789146374267, 
    16.6552019557444, 16.7045311777538, 16.528786167458, 15.7228090003924, 
    15.2407307027132, 16.423976871727, 16.3589512351464, 15.9507335863898, 
    15.2015649332994, 11.4977936219781, 10.8578788242334, 10.9036461580754, 
    11.1592863640127, 11.3092174991524, 11.4583742514404, 11.0541854997406, 
    10.0773717393039, 8.5104131022696, 7.54026427296393, 9.17328851815845, 
    8.06579065073576, 7.06831871243231, 9.44777038169996, 8.03917345975186, 
    6.84437163650041, 10.211641231758, 8.75140924037809, 7.40175498009556, 
    6.45474050725283, 11.0264177004692, 11.074453274149, 11.2689333407061, 
    11.5342388873466, 11.7076733307625, 10.9893742617517, 11.4812782167026, 
    14.7019848483224, 14.5325228954299, 14.3255615625171, 13.5060045530894, 
    12.6762033205653, 12.173425170589, 11.6966791376585, 33.1686793489075, 
    33.1576613443559, 33.1516966516225, 33.1381315108662, 33.1517491716455, 
    33.173314557462, 33.1838080432533, 15.0103007235372, 14.7287029121382, 
    14.2525943272631, 13.5668114834649, 13.0375728661524, 12.5440248207675, 
    11.6852212231139, 11.0536826272126, 10.3384627611212, 33.2052068648637, 
    33.1936418495889, 33.179502971793, 33.1690490281673, 33.175219861216, 
    33.1916822242255, 33.222209833503, 33.3295532297698, 33.630713953222, 
    17.7097507265736, 17.7398021159128, 17.6634827621919, 17.2183817389147, 
    17.216714407284, 16.8969469015738, 16.7926597822524, 16.6309681941824, 
    16.5617849484201, 16.4706414653913, 16.4744622424109, 16.4201663335419, 
    16.0933169946967, 15.7279081819626, 15.1285360005434, 15.1166867873794, 
    14.7069870486725, 14.5334110698588, 14.249610665578, 13.9293730867336, 
    13.5534093706105, 13.3862557959785, 13.1577042568037, 13.1453750722148, 
    13.5466538587984, 13.7701787269163, 13.6310881567458, 13.2139549824669, 
    12.6827277798832, 12.2326456667565, 12.2797284029859, 12.33027656001, 
    11.9597642124855, 11.3544042859991, 11.0691764892911, 10.881023732696, 
    10.4894185017982, 10.6676034703267, 10.8575290259478, 10.9434317802821, 
    10.7169882375299, 10.6831486832115, 10.667639804368, 10.5369617910405, 
    10.4347465497058, 10.2809626651701, 9.94286301076958, 9.73734296112276, 
    9.57974976116088, 9.41633410910533, 9.26254660686186, 17.6262743207678, 
    17.7013555562145, 17.6993655114219, 17.4224604483866, 17.0713493083846, 
    17.0396657387868, 16.6720590898872, 16.6547279452408, 16.4769682665084, 
    16.5651994140173, 16.328191278055, 16.3136201682654, 16.0440943435656, 
    15.7950381168494, 15.2970431620465, 15.0705574029111, 14.5608714498809, 
    14.5637356805207, 14.7499345713149, 14.1732763588582, 13.7461749512605, 
    13.6926743005449, 13.634256168254, 13.6422326656409, 13.9375421239553, 
    13.7968258302917, 13.7469005098064, 12.872808784504, 12.3715698716117, 
    12.2055642148544, 12.0327687844258, 12.0189608823945, 11.7309113363049, 
    11.472543211775, 11.0965322038131, 10.9447736307953, 10.653588151673, 
    10.8323049951335, 11.1719938644963, 11.1827977195481, 10.9497017858719, 
    10.7485110484389, 10.6587430481964, 10.5212955242237, 10.3075384010836, 
    10.1727304864077, 9.81789751786791, 9.71173705147674, 9.56892277965051, 
    9.48182987035387, 9.25946210544775, 17.5358272535418, 17.4522986771294, 
    17.4764364711703, 17.3111221706568, 16.9572643383978, 16.7494863074257, 
    16.4959448976616, 16.5126023109649, 16.4073215271187, 16.4916875755432, 
    16.3393737285596, 16.3715540941589, 16.1139299655021, 15.904788269551, 
    15.522773852547, 15.2614059844416, 14.8824516462583, 15.1611292730576, 
    14.7905099924363, 14.4086746582248, 13.9675838923466, 13.9369644173246, 
    13.9559675853798, 13.9425520255474, 13.9452119977987, 13.4208835179127, 
    13.1430521584226, 12.5920446155343, 12.3107830391449, 12.1103300660316, 
    11.9664690452053, 11.8975706853692, 11.8097754291053, 11.7787187685341, 
    11.29790170585, 11.122520330964, 10.946360453305, 11.0147659623112, 
    11.2997166131347, 11.0627652105678, 10.7598424529765, 10.6683898752576, 
    10.5592354671575, 10.2801507371108, 10.0411754964456, 9.91627033018185, 
    9.60833503621416, 9.59141496048528, 9.51383056268924, 9.61533510012202, 
    9.4235689540716, 17.6558295678935, 17.3953901709183, 17.3151553120308, 
    17.101126271356, 16.7446850509232, 16.514715639331, 16.3870637235113, 
    16.3774071129792, 16.379264599366, 16.5046800053124, 16.2768935680977, 
    16.2955070800313, 16.1868376301382, 15.9485175479525, 15.6364359792545, 
    15.3238593461622, 15.1064023072762, 14.9326157684933, 14.37312893689, 
    14.1885338219989, 14.1421613958388, 14.1774941751154, 14.1940416172406, 
    14.1391332185982, 13.765028302184, 13.1181489503401, 12.8982981612399, 
    12.3343834035411, 11.888561048356, 11.5586204280332, 11.7416284004094, 
    11.6588742054565, 11.3777823493618, 11.7161275479074, 11.4071236389645, 
    11.2795544148103, 11.1394030373597, 11.2490337030679, 11.3409895055617, 
    10.8745138406226, 10.6791769202409, 10.6269882334197, 10.3018157027902, 
    9.88083219502552, 9.67370112059357, 9.47583786405763, 9.39204681645855, 
    9.3802737117198, 9.50804171907304, 9.49467005996039, 9.37313893403071, 
    17.7025730027694, 17.4938860145448, 17.1633740808815, 16.9851485539666, 
    16.7395699826476, 16.564784034593, 16.3966194339668, 16.4189399895952, 
    16.3360457305613, 16.2467062710238, 16.2175077225949, 16.24952654527, 
    16.1296322940101, 15.9339001127245, 15.7017129287906, 15.4023487069204, 
    15.1652171515717, 14.1072252717839, 13.3274935595546, 13.2857733807144, 
    13.5649969796027, 13.6995083734346, 13.7836208243481, 13.9522836848406, 
    13.6979742069483, 13.1394641319511, 12.7247793415403, 12.0145891884752, 
    11.4725522593499, 11.2572276909567, 11.3751970720854, 11.3986505495132, 
    11.3183061612016, 11.4277944580533, 11.2826117422119, 11.1717195007293, 
    11.0178169514543, 11.0874984917915, 11.1643138608174, 10.7891561696343, 
    10.4438837959837, 10.4599896433079, 10.1209292144312, 9.72001039321294, 
    9.6661972405252, 9.37092814840595, 9.39027746326017, 9.50837636220084, 
    9.39231477743651, 9.41353462331925, 9.37873695264095, 17.6550138851716, 
    17.5152496653895, 17.1435880818428, 16.8923716695617, 16.7828084587209, 
    16.6125848472408, 16.2962071664727, 16.3169097134703, 16.1965214284401, 
    16.0142405872526, 16.1005319233216, 15.9614887080228, 16.0314317718305, 
    15.8241890807523, 15.7354902411181, 15.5808221465915, 14.9902508745502, 
    13.6753235380005, 13.0652498134316, 13.2257436313744, 13.2689652099283, 
    13.5809910163636, 13.6211715316963, 13.799628722764, 13.5072630764633, 
    12.9151731695219, 12.4807665983383, 11.7051890754507, 11.1064184324531, 
    11.1710853706724, 11.1505602705845, 11.2784882065868, 11.0434917684956, 
    11.088510981328, 10.8288911976429, 10.6502196992614, 10.5996994979323, 
    10.6615597147891, 10.9697872499044, 10.7197040578169, 10.2812119006043, 
    10.1470291630582, 9.94226204833367, 9.71067181321763, 9.75447050326873, 
    9.39121513239526, 9.35557947045449, 9.46090547013283, 9.3370024340389, 
    9.3504708790803, 9.40154883618234, 17.6062788858651, 17.361794238333, 
    17.1328201582947, 16.8046346960279, 16.9312235253781, 16.686664724191, 
    16.5303490829515, 16.297379381832, 15.9264193370836, 15.9358415824926, 
    15.9835079860982, 15.8565317075359, 15.7459004249166, 15.6335202783965, 
    15.4735771360713, 15.0061486499249, 14.2946931652638, 13.2403558460463, 
    13.0149340866194, 13.2434799910741, 13.312574267738, 13.3910921969281, 
    13.5411068638787, 13.6307306863226, 13.2566740186811, 12.5671936911351, 
    11.9908283141593, 11.1560281424026, 11.1259201122558, 11.0430119968788, 
    11.1546806780454, 11.2406775257917, 10.9161945468839, 10.7435930597942, 
    10.5878074212238, 10.5548722675876, 10.5011463279388, 10.5636353594482, 
    10.7724554066558, 10.7224238782463, 10.3977883924159, 10.0552947020456, 
    9.78301064994744, 9.72087749779106, 9.86792381861858, 9.60139774258037, 
    9.32858648308381, 9.33895830548757, 9.2324502761086, 9.38571801134301, 
    9.32289052642252, 17.6043275113336, 17.4315129955822, 17.1165122613439, 
    17.0781044431214, 16.875932423692, 16.8483303722004, 16.3544325150053, 
    16.1957615976489, 15.7967409821413, 15.8966045166123, 15.6999754646305, 
    15.533152243858, 15.5153517129741, 15.4116811014763, 15.0553250014989, 
    14.224052735523, 13.5970794249924, 13.0204055603205, 13.0030315477016, 
    13.210382672428, 13.4534526697969, 13.3960042045313, 13.3934365910372, 
    13.4583360195091, 12.9374199946253, 12.1478255533295, 11.4960859930902, 
    10.8913390411266, 11.0563706443342, 11.0228042879924, 11.0446681741484, 
    11.2304032230629, 10.8106891109179, 10.4857991329601, 10.3658814614822, 
    10.4172912572799, 10.4086943393695, 10.6210039537816, 10.6626897903847, 
    10.7255839695191, 10.8210872497668, 10.4929016151088, 10.0793853675574, 
    9.95828836758617, 9.94424193276671, 9.92217894712232, 9.53742914511865, 
    9.24240891510777, 9.22691729811142, 9.54568054632322, 9.42343766406105, 
    17.7023937313751, 17.6240042523748, 17.4715236928041, 17.16752568711, 
    16.8123510879512, 16.6352084073807, 16.4201929396495, 16.3980783687382, 
    15.8689701757111, 15.7276880843063, 15.2943579078574, 15.0086291615116, 
    15.165544111617, 15.3613631087753, 15.1811604384189, 14.3028795927999, 
    13.4643272863736, 12.9511637936387, 12.7989991708824, 13.1304972062483, 
    13.4449040773422, 13.3998269205156, 13.4314000629916, 13.4536257524332, 
    12.7751130086914, 11.8747608149675, 11.2622930299573, 10.9073779363711, 
    11.1279108182012, 11.1528599300352, 11.0544730593175, 11.1599898897316, 
    11.0343076163853, 10.5454022442312, 10.3243742051516, 10.2958617907827, 
    10.3755970781997, 10.4970969696748, 10.7228361064544, 10.7810636767382, 
    10.9426304196177, 10.6936926808168, 10.3188093787615, 10.185901919098, 
    10.0780208551553, 10.0043150156989, 9.63960446558013, 9.13712186669058, 
    9.09923328199745, 9.58129474051833, 9.64479444423134, 17.7631077458316, 
    17.5548150848337, 17.5260806217685, 17.2925927665077, 17.0339660990896, 
    16.5162014897119, 16.4376696478621, 16.1497322112235, 15.9817557754488, 
    15.4354903646108, 14.7892760659206, 14.5301187406617, 14.6532151373108, 
    14.8832743572239, 15.0710450813161, 14.2272529384705, 13.3412462967837, 
    12.8562082253664, 12.7099054867052, 13.0469135337517, 13.368634365221, 
    13.3539025423493, 13.4347480726321, 13.4347903632368, 12.7481865648522, 
    11.7446682058833, 11.1806577668531, 10.9510435640183, 11.2114122014591, 
    11.360403147652, 10.9875665209469, 11.0587968711757, 11.1807866908033, 
    10.6700210695459, 10.5541046600881, 10.4096795910809, 10.4590058711044, 
    10.5047368393628, 10.7206298366442, 10.7587937299932, 10.7742860212918, 
    10.5872170840404, 10.4049651248923, 10.297334117711, 10.1593787840563, 
    9.97610371259715, 9.85104448993683, 9.02912054384606, 9.08666686196185, 
    9.48425182409536, 9.80922636382659, 17.6570708869063, 17.4176547878141, 
    17.2161771229303, 17.2185216241679, 16.9629451562159, 16.7777357489101, 
    16.5079936829721, 16.5143391059719, 15.9855582166597, 15.4179662879223, 
    14.8179683061695, 14.5647751836333, 14.3954157665847, 14.344252139542, 
    14.4325693767614, 13.8021904635083, 13.0413299893832, 12.7584526039273, 
    12.7298886462404, 12.9796154361308, 13.2215179881146, 13.2248313676478, 
    13.1759689338018, 13.1810901505407, 12.7185262602587, 11.81500358606, 
    11.1677318317731, 11.15778221636, 11.5604448851172, 11.5099913732758, 
    11.0023187186371, 11.083195639459, 11.0510994283316, 10.7503341345317, 
    10.6683167707767, 10.3639773133047, 10.5973236342355, 10.6058651045168, 
    10.7287371896225, 10.5571842953499, 10.3211233251312, 10.2773266532891, 
    10.2216031718001, 10.1597839507255, 10.0956045894391, 9.91368366733541, 
    9.67910119670077, 8.98599407310795, 9.35564780048916, 9.67639737042009, 
    9.81280778777503, 17.2270248176146, 17.3692333397173, 17.3302518435258, 
    17.2086264664833, 17.1755361856588, 17.0228620825213, 16.8494402222685, 
    16.4165894030853, 15.8662021617032, 15.3654119330462, 14.829020102073, 
    14.6657798560185, 14.5415460581383, 14.3545232376368, 14.0999535189779, 
    13.5547214220725, 12.9225035664176, 12.7088649937063, 12.738004204267, 
    12.8345700879588, 12.9791357776892, 13.079042314174, 12.9605476372447, 
    12.8578327071169, 12.5580560557531, 11.9177505446699, 11.3047952283465, 
    11.4081911724965, 11.7311657569962, 11.5851442084321, 11.1200538343041, 
    11.0625221637224, 10.9822034288518, 10.9109796956871, 10.8065130500888, 
    10.6655322739022, 10.6619305375296, 10.6484669406525, 10.6966755807218, 
    10.5123587227305, 10.3031192080803, 10.1797477874472, 10.224788871855, 
    10.2275166719514, 10.1420939223411, 9.93260698450897, 9.6336451380022, 
    9.14696235235934, 9.6423128507956, 9.87461253843348, 9.74643938948395, 
    17.0088399031772, 17.0728748336525, 17.1567224473107, 17.2245807001481, 
    17.2378882079963, 17.3444799193718, 16.9193355203692, 16.3349978167095, 
    15.6942640512455, 15.1188996187743, 14.7660695666575, 14.7050494843373, 
    14.5711370144528, 14.4598986226054, 14.1381468237951, 13.5887660024397, 
    13.0814297346701, 12.8549342535881, 12.7301350474798, 12.6098716350882, 
    12.5713907575253, 12.7545265847603, 12.9706588942536, 12.7484158315637, 
    12.401512275104, 11.959695573164, 11.5725433664119, 11.7955264255862, 
    11.977877255467, 11.6471528650053, 11.0859100551482, 11.0593403687553, 
    11.0357046540481, 10.8464819794567, 10.7282787327922, 10.6437837465701, 
    10.5780896215909, 10.5436702557648, 10.6557535177356, 10.4882014645237, 
    10.4173686352334, 10.3947611621409, 10.3061524694624, 10.0526113760997, 
    9.91058319784741, 9.72607069646121, 9.39382433156328, 9.34174053359759, 
    9.6293388407412, 9.64240023489274, 9.57327150286731, 16.8108326812184, 
    16.9093121139716, 17.0311542828906, 17.164125014636, 17.3546687634539, 
    16.9366588712306, 16.6866066087087, 16.1745686091752, 15.6461329770867, 
    15.1023551236375, 14.8198235994041, 14.8176550095712, 14.5722449459649, 
    14.4225781264466, 14.2354557278251, 13.6626806929135, 13.2221317912704, 
    12.9556961332271, 12.9066930883605, 12.7342831456092, 12.5203420663598, 
    12.4493349664671, 12.8348441563556, 12.7320112030005, 12.695595501353, 
    12.2034093920353, 12.4186793041367, 11.890502681765, 11.8929468463022, 
    11.5592920908821, 10.8771164708575, 10.9868012515491, 10.7348151035473, 
    10.7388266313334, 10.7667478492325, 10.4623020855005, 10.0795594450055, 
    10.2789420016847, 10.3186227525845, 10.2406015716424, 9.89972274066075, 
    9.39350067705834, 9.07301933758222, 9.33588179905932, 9.56146920756605, 
    9.29547988171577, 9.28399559760725, 16.650006866518, 16.6579868802429, 
    16.7448282432917, 16.93563120903, 17.0351003014548, 16.9743134940211, 
    16.5732277471609, 16.1132037043384, 15.9132366615001, 15.1388118234643, 
    14.8819984292056, 14.6974090007833, 14.4255420917241, 14.4432735296473, 
    14.4965282935444, 13.8166683723787, 13.3085999709159, 13.0943031473044, 
    13.090239934969, 13.1634423847711, 12.7865985265944, 12.3834423274707, 
    12.6488219293037, 12.8454495461497, 12.9558879414688, 12.6067471465802, 
    12.4301365354771, 11.3472941505053, 11.6723314846066, 11.3893789153756, 
    10.7145423561948, 10.7157574939757, 10.5249635202737, 10.6312337810015, 
    10.6421800849781, 10.4374788436013, 10.0677493449479, 10.0130742978805, 
    10.1078619352333, 9.96305810518, 9.4515474622927, 9.25124672227668, 
    9.23103976902999, 9.48749965320391, 9.44371021395447, 9.28458235949869, 
    16.7118426699076, 16.5919782343871, 16.688697457245, 16.781291252959, 
    16.7894875794198, 16.6358516647511, 16.5089840289473, 16.1704206760532, 
    16.0403804509915, 15.2620890375698, 15.0307968303721, 14.5864079283305, 
    14.3724333987182, 14.5065470517222, 14.5276728920842, 13.8146666024285, 
    13.3363385411334, 13.1664519150133, 13.3039439905555, 13.3301382654044, 
    12.8657865476777, 12.409926313509, 12.2991577067283, 12.6665095111778, 
    12.9257905366465, 13.0424197970778, 12.1109525878687, 11.3658075613749, 
    11.4761180704032, 11.4337296121074, 10.8792298580434, 10.8521379234759, 
    10.5337993351453, 9.84376494052953, 9.77644344255796, 9.54766873779567, 
    9.4275387501126, 9.37217684577455, 9.4909348549127, 9.48799645959115, 
    9.55338222079802, 16.6116528751373, 16.620721478322, 16.5927303702831, 
    16.5513287836764, 16.3986630628715, 16.3140900926077, 16.5697569530761, 
    16.2984220531059, 16.1982387201691, 15.5433197804319, 15.3193456423452, 
    14.7186729736745, 14.1040898181518, 14.2717725053289, 14.3374751238938, 
    13.8178930766283, 13.4878526181125, 13.4332134273907, 13.5912478001602, 
    13.4524075667286, 13.1395661274166, 12.6298838645562, 12.3720400931554, 
    12.3409494244881, 12.6605406715297, 13.1059699818585, 11.9425092092307, 
    11.4530736319275, 11.5938323601977, 11.2792476419508, 11.1156513078101, 
    11.1134901230078, 10.0712896851101, 9.62749797114963, 9.52017663432942, 
    9.32491414147399, 9.38492406998736, 9.08112447630671, 8.90512244137895, 
    9.20410060972335, 9.22674074210911, 16.7391626619586, 16.750725364893, 
    16.6607657578604, 16.5032023905812, 16.2493984282722, 15.9250515380088, 
    15.944614023703, 16.3329321447117, 16.1807942244631, 15.7706877078225, 
    15.2421434076142, 14.3734480799257, 13.9214778259258, 13.9893764766224, 
    14.0627395849734, 13.939095490391, 13.8113059666227, 13.7378363579481, 
    13.6114359455089, 13.4136006551708, 13.2156983584821, 12.7044674441039, 
    12.5753966564285, 12.3975658360937, 12.5113260392663, 12.7228132241297, 
    11.8037735841375, 11.4183777143353, 11.5929969995497, 11.2488192750078, 
    11.2162076116677, 11.1134901230078, 9.64723075408535, 9.41568903272522, 
    9.14461383420702, 9.09362538210868, 8.77826056184328, 8.53458799151915, 
    8.63482090089082, 8.58372609246417, 16.9401015761728, 16.6723667593627, 
    16.6516416852176, 16.5329277335977, 16.331547291087, 16.0697913580969, 
    16.0620571375435, 16.1511435425161, 16.2200226420176, 15.910485825975, 
    15.0194295504214, 14.1643059527792, 13.8280725789598, 13.828436265632, 
    13.7230415390177, 13.841723441903, 13.9741390051263, 13.8485572619691, 
    13.3035034712587, 13.044016301917, 13.0170056254361, 12.8267846918825, 
    12.7209215739629, 12.226558810942, 12.0157003462362, 12.2903280662764, 
    11.9271009535539, 11.4546446388989, 8.91431894531683, 8.97541060803605, 
    8.67428604789451, 8.12589556955253, 16.8099744376938, 16.5789189200971, 
    16.4980257696988, 16.4187977722562, 16.3417837012985, 16.1136161307346, 
    16.0956941070459, 16.0193831990596, 15.7281742548459, 15.2139124988089, 
    14.7756380244286, 14.1041180008311, 13.9859157283261, 14.1708837777022, 
    13.8171965560778, 13.3843328423363, 13.7614337669119, 13.5607488139714, 
    13.2367366472139, 12.8932274939952, 12.7803978427082, 12.6753516515357, 
    12.5425965481997, 12.1910889697979, 11.8225219679276, 16.7188140567405, 
    16.5245726248579, 16.4538763077853, 16.3041639869534, 16.0864190938756, 
    15.771588610438, 15.356439627165, 14.9472970397149, 14.5200024584222, 
    14.3584778863135, 14.4178552705281, 14.0756709930582, 14.2199734934706, 
    14.2989542025996, 14.0271684622967, 13.3065029709532, 13.4371663865272, 
    13.4950121374036, 13.3333890803934, 13.1441206750444, 12.988656664193, 
    12.7460185731678, 12.5292432517153, 12.1494175362052, 16.7300635577496, 
    16.5436834087726, 16.4568011582953, 16.1557717219953, 15.7525870401325, 
    15.2677817742775, 14.7249988309498, 14.3465860961567, 14.1750027735782, 
    14.2034682447753, 14.2192341500746, 13.9764585609405, 14.3720956845641, 
    14.2584388842442, 13.6043954464768, 13.2759204937865, 13.4265866226213, 
    13.5299119133937, 13.280060650315, 13.1581632762731, 12.9514861568871, 
    12.4919342364582, 16.7049891553443, 16.5991421920483, 16.5180936387126, 
    15.9868261823303, 15.6313301606684, 15.0500460715044, 14.4305151128264, 
    14.1725141153666, 14.2437212192099, 14.2567477052139, 14.2753381102772, 
    14.2825541683321, 14.2486095747736, 14.0706668135876, 13.6468670100529, 
    13.3962281507287, 13.4980115009439, 13.3178916539748, 13.0108671843585, 
    12.8281795227425, 12.4178901860826, 11.9195534324931, 16.6053105307391, 
    16.7560590849887, 16.6278311907786, 16.0303497756032, 15.596204831518, 
    15.0107206987307, 14.3253629095287, 14.2773474196589, 14.3565219624368, 
    14.3312290387275, 14.1604005252306, 14.066480243615, 13.9858659931753, 
    13.7572039616853, 13.5652028081179, 13.4445037358096, 13.346616830902, 
    13.1696813123117, 13.0437838290975, 13.0928497206384, 16.6334596446216, 
    16.8476629922356, 16.6748390637419, 16.4899243824965, 15.9175783806432, 
    15.2136035971154, 14.3856745251139, 14.3365694175456, 14.3969036910189, 
    14.3413623870294, 14.1786349807428, 13.9010242239125, 14.038879392503, 
    13.7875285294146, 13.614507470473, 13.4972681052096, 13.3711415287768, 
    13.2819930352088, 13.0591091981935, 16.5873606019382, 16.761454587497, 
    16.7280351421303, 16.7168726160027, 16.2554820803626, 15.4719620891155, 
    14.6513916651933, 14.6809884874847, 14.5569368283555, 14.333943183744, 
    14.360946503741, 14.0093947096995, 13.9676200102836, 13.9907900234386, 
    13.7895188377358, 13.5017268086926, 13.4131499961355, 16.3164100550475, 
    16.2401937704721, 16.2725860025117, 16.5393135873723, 16.725716611869, 
    16.0214702952981, 15.3738766629061, 15.2373784638448, 14.9793359995479, 
    14.6661823047847, 14.321751816956, 14.0904965732883, 13.7694754009327, 
    13.7245521553629, 13.5807977811106, 13.572648520837, 16.1847385394, 
    16.0748054337595, 16.024335143151, 16.3823456522308, 16.8118326527244, 
    16.3699392506193, 15.9260525185825, 15.7886506458623, 15.4281771471194, 
    14.8878365459441, 14.3077153495391, 13.7690841473184, 13.1847433350907, 
    13.1594076251666, 13.0409295032732, 16.2690528538858, 16.1538982089965, 
    15.9747308077419, 16.162658046484, 16.5194054193891, 16.6167311055605, 
    16.284175239941, 16.0090311715527, 15.5386225855729, 14.6551199648494, 
    13.8978579227103, 13.6444438817727, 13.2323784850774, 13.0132140969171, 
    16.45835016866, 16.4179187229187, 16.0753180609453, 15.9472259525635, 
    16.208011810634, 16.5021913322433, 16.2139320318948, 15.7587078781068, 
    15.146412888221, 14.3554983315089, 13.7857308698429, 13.661100446579, 
    16.4942402878176, 16.4905494626294, 16.1687836069946, 15.8258694121971, 
    15.8400596576068, 15.9524772748147, 15.4790037079728, 15.004706249774, 
    14.8307272082626, 14.4592181800519, 14.0061477606446, 13.8023519821077, 
    16.4405286430494, 16.3842009987554, 16.0727174336037, 15.7844623971588, 
    15.577534294074, 15.4223109255067, 14.8393976177861, 14.5818585936996, 
    14.4979999007787, 14.1767797523979, 13.9890923244733, 13.7944905591849, 
    16.4230822084695, 16.235791255464, 15.9290829704911, 15.8543959072495, 
    15.726376746704, 15.4029071518788, 14.939046160404, 14.5899925483509, 
    14.4631478168193, 14.1783885865422, 14.0210461870322, 16.3641948706112, 
    16.0463773761801, 15.8928481158884, 15.8209582994797, 16.0343240877077, 
    15.7033513177627, 15.1670619530771, 14.8122727469001, 14.6163242101435, 
    14.4445871422715, 14.2808568942525, 16.2047486290228, 15.983093282988, 
    16.0721372299585, 16.1891288823514, 15.9936016590579, 15.5204953525012, 
    14.9626900992166, 14.9328295834212, 14.7463962978931, 14.5123093399964, 
    14.4471619956027, 15.9619049291403, 16.1314207288783, 16.1978123233374, 
    16.0568544486574, 15.7378853718079, 15.2901224310093, 15.1827935386068, 
    15.3680886263463, 14.9667811384298, 14.7302333270285, 15.8374415480355, 
    16.0080602860304, 16.1429407180737, 16.0746408115682, 15.8900029875236, 
    15.5916543551889, 15.609807967171, 15.8183269989463, 15.4990526408085, 
    16.2152056958065, 16.0445273645106, 16.1024661648189, 16.1127112161434, 
    15.8574848817857, 15.836532648011, 15.8625563040374, 15.938069710427, 
    16.1071103906274, 16.6816979888929, 16.564040157849, 16.3990912675518, 
    16.091865382421, 15.5442063457806, 15.8363635785793, 15.8947545622492, 
    15.2219256205235, 16.6817903726313, 16.6872296752444, 16.5724585722431, 
    15.841950017888, 15.4219807344811, 16.4274596878165, 16.3663907776182, 
    16.1947858981375, 15.38525878032, 15.6171659763143, 15.4651861397109, 
    15.4872820878052, 15.3695931108268, 14.9887936463017, 13.1219773445358, 
    11.1724806551414, 10.128639631279, 9.50431016378758, 33.3123124792657, 
    33.3006701839634, 33.2952443050418, 33.2800871059008, 33.2363166261495, 
    33.1805199998615, 33.3270137083095, 33.5632675822285, 33.8386930339166, 
    15.2674554356953, 15.2794483342085, 15.2456896392988, 14.9234733246897, 
    14.2047800247701, 12.8986687939224, 11.426766569333, 9.92538191501012, 
    9.07370170095552, 8.64474562771993, 8.15208317127087, 7.59173616550716, 
    7.07691570651543, 6.69379782518565, 6.55000861275002, 33.173543546319, 
    33.1689904605485, 33.1590103854622, 33.1377155600685, 33.1460856138357, 
    33.2354938729723, 33.4329800663649, 33.6264895398707, 33.8067475127655, 
    33.9376236089436, 34.0347795257609, 34.1307632290394, 34.2129291392609, 
    34.25720581029, 34.388646099678, 0.197824782840204, 0.180469218404196, 
    0.188445161974712, 0.165671756525717, 0.16772508692714, 0.16384638193536, 
    0.155979116967203, 0.177630497070844, 0.153907757222638, 
    0.182893488251502, 0.199703511571511, 0.157467286617847, 
    0.182906687823471, 0.215794980096309, 0.175261619447371, 
    0.179780248034664, 0.173740651357433, 0.218644747205691, 
    0.182937815125447, 0.205569575805032, 0.154462680350972, 
    0.172227728542468, 0.21629119835118, 0.176015521142883, 
    0.217967557208211, 0.135181802260459, 0.186463925477623, 
    0.201013199591387, 0.148285094151533, 0.179398914331211, 
    0.212655966751653, 0.135845030537645, 0.178783577268016, 
    0.185214258801659, 0.129119285242724, 0.191100327850558, 
    0.190874417236768, 0.146930918267874, 0.152295441180179, 
    0.173738709933567, 0.172172802738851, 0.128773528972439, 
    0.185880152822542, 0.171470609197178, 0.156569136432295, 
    0.131139156357613, 0.168992098352662, 0.17968397566506, 
    0.142507282343433, 0.166848819743709, 0.159969350932356, 
    0.127896152478534, 0.157593877852182, 0.128084789843262, 
    0.169525587780034, 0.185332751537195, 0.151554967267738, 
    0.150607171208192, 0.156830714972833, 0.146293684944379, 
    0.149686188395422, 0.135320477394655, 0.17839196472881, 
    0.178925278252492, 0.112661355024417, 0.151932304931423, 
    0.14744533785443, 0.156900004008598, 0.185639695205316, 
    0.142407761210167, 0.140845301677809, 0.184629072746856, 
    0.168219327230211, 0.129521425989896, 0.143473176252807, 
    0.151042166460657, 0.163809540929736, 0.196990676650072, 
    0.143625840902574, 0.113467410816279, 0.14127280447523, 0.180101368879, 
    0.16946047789137, 0.177136126804336, 0.13859427276836, 0.152621023925298, 
    0.170726531858965, 0.191194822830476, 0.144705712327298, 
    0.12082507056877, 0.137783377288317, 0.18089011848133, 0.176133139891099, 
    0.196758403859291, 0.140660395572506, 0.0971109385927634, 
    0.150563150740904, 0.172257957747298, 0.191594385937124, 
    0.142067282371772, 0.158521046133897, 0.135596259557086, 
    0.188464574968997, 0.177398719683198, 0.19205099911402, 0.14990662802171, 
    0.114494587676959, 0.149618928167001, 0.181579134567257, 
    0.198750234347173, 0.13959527149165, 0.179144830620356, 
    0.140219404672882, 0.195067787087067, 0.0819849346974468, 
    0.176772601803767, 0.1913762091523, 0.152992468852548, 0.140645430235169, 
    0.149781392043573, 0.195953230023696, 0.212894752396424, 
    0.142862225080266, 0.17920122055413, 0.148100619554691, 
    0.184681905256387, 0.106411544917241, 0.173912553518696, 
    0.197360782471481, 0.148040569515058, 0.157750165808681, 
    0.150907794489039, 0.198963547844185, 0.0866646286922883, 
    0.221442155161155, 0.147631977886687, 0.179880623845331, 
    0.156097016193785, 0.156049051515194, 0.127336797059606, 
    0.172029248608213, 0.212817376000852, 0.144573436511953, 
    0.165444728454005, 0.15273434330262, 0.190237834645961, 
    0.103256562338216, 0.222234568506599, 0.155589754043042, 
    0.185758760661454, 0.149608900728102, 0.128227248260673, 
    0.140028234382631, 0.169480408612148, 0.0982511308334105, 
    0.228937117075325, 0.141603185036857, 0.168234946017181, 
    0.155743268648235, 0.163916581463099, 0.105699364653471, 
    0.219102506008885, 0.166244441805238, 0.197382912277815, 
    0.142468798295114, 0.103753351620684, 0.146350807563333, 
    0.164686587916665, 0.108188736745062, 0.236637339937798, 
    0.14362360174084, 0.170076350094589, 0.146843258783122, 0.141751052174, 
    0.0973503269359525, 0.211128292513356, 0.176896757478306, 
    0.0914936480540682, 0.215488052152264, 0.131795046695744, 
    0.0830410962966557, 0.144158248245137, 0.158100789488289, 
    0.0962822381057229, 0.230801214623497, 0.145940645213365, 
    0.175818599881816, 0.13644929743568, 0.122601705310382, 
    0.0842721088999533, 0.202543855196771, 0.186501342837048, 
    0.104387833962062, 0.23082803929724, 0.13269103276157, 
    0.0614640116129389, 0.1399274219005, 0.146981742968096, 
    0.0771298291397016, 0.224754917419681, 0.155087600743821, 
    0.0742871147506459, 0.18737303743729, 0.126409667310517, 
    0.103077602769677, 0.0714469777287925, 0.189250054709799, 
    0.189147286673648, 0.0924208044432401, 0.229401766233471, 
    0.136148747963004, 0.0445485982453593, 0.142516703160276, 
    0.134507102544733, 0.0637301195496639, 0.219055361010554, 
    0.165410247514427, 0.0935026177426185, 0.19871785144332, 
    0.125052997604591, 0.0785105795537134, 0.0639491571776242, 
    0.173688540299109, 0.186461651870217, 0.0760506368655824, 
    0.231949624143609, 0.138748893068437, 0.0661167073182383, 
    0.0513346648848255, 0.15088665936919, 0.123142940011248, 
    0.0534763105744101, 0.209673181902769, 0.17789750009499, 
    0.0919647171918663, 0.201043340911983, 0.12102773971955, 
    0.0629239570887279, 0.0677094230681623, 0.152965179764553, 
    0.176720949665695, 0.0678816064128914, 0.233010968387332, 
    0.148107222237752, 0.0955950800678819, 0.0763235166350427, 
    0.159919569480722, 0.114613488288192, 0.0478543354118436, 
    0.191152463353281, 0.17832861487989, 0.0798976803145172, 
    0.20752606702799, 0.120763399884823, 0.0813539853672027, 
    0.0780468505441215, 0.0770507598814636, 0.123028694296881, 
    0.159060273856331, 0.0555796894274956, 0.223922279822993, 
    0.157757537092308, 0.0946366440102374, 0.0982125623324704, 
    0.164941749561767, 0.105075031959304, 0.0545604436954336, 
    0.163149639853416, 0.17595180450394, 0.0681065532240747, 
    0.215557382386743, 0.120506366324107, 0.103537708463377, 
    0.11132797141376, 0.0867522989650037, 0.0879223885526377, 
    0.128488308047946, 0.0492022473054462, 0.200417465881826, 
    0.15981006494434, 0.0748246175913295, 0.110474112072077, 
    0.172047235094264, 0.0968321358490775, 0.0963111991748489, 
    0.0709720012774257, 0.121678135960477, 0.162957627270869, 
    0.0579293486946612, 0.211427116060959, 0.120149369576415, 
    0.091451401120385, 0.130154699127226, 0.0940119084167084, 
    0.0509687304056438, 0.104775504522493, 0.0615345999897685, 
    0.169658498831303, 0.157077356156645, 0.0495623122867313, 
    0.121618726762697, 0.180518473369502, 0.0889853421703378, 
    0.107667259345634, 0.0780125317461478, 0.0723539575068216, 
    0.141280430754681, 0.05840327240229, 0.195054903077154, 
    0.114935965007168, 0.0625208222434172, 0.129610094183386, 
    0.10181736104095, 0.0255343561565831, 0.10899552518046, 
    0.108493601241531, 0.0800103528910831, 0.126155541404424, 
    0.152135306036473, 0.0471973546419739, 0.13046884826503, 
    0.179804817499404, 0.078364271653437, 0.0939089362891187, 
    0.077388559552295, 0.0182255891010092, 0.122035609408684, 
    0.0724969432042726, 0.16780755409588, 0.109547532197682, 
    0.0339372400660961, 0.129146165523854, 0.110058944000319, 
    0.0137704525780775, 0.11389050980412, 0.13157600808679, 
    0.0787484117557636, 0.0718647125009907, 0.146425321356015, 
    0.0542701003303134, 0.119905421925197, 0.171620855207666, 
    0.0670125647541317, 0.06557726378501, 0.0815982199004448, 
    -0.0166131140063076, 0.117333664467556, 0.121920020886245, 
    0.0863733707485529, 0.131415934913569, 0.110238574819389, 
    0.0305167306085061, 0.134168287560439, 0.115074802649157, 
    0.00520557258891455, 0.10299055767279, 0.125246191166709, 
    0.0699150263863239, 0.00830912923057501, 0.135183359918416, 
    0.0502053729175934, 0.085191734218716, 0.153839203663287, 
    0.0621498693889559, 0.0325387306167622, 0.0869904408005027, 
    -0.0261068464868015, 0.120729259413283, 0.127190517316589, 
    0.0793650973224091, 0.0871126368861764, 0.119708525516238, 
    0.0248187995868317, 0.125393910417287, 0.122767566630919, 
    0.00466012688519691, 0.0791541179498543, 0.0786087314843674, 
    0.0744979361925069, -0.0380764058073957, 0.111785870033452, 
    0.136573066851444, 0.0472548196038676, 0.0410722004019958, 
    0.125564570263381, 0.0657958361472153, 0.0155426113611453, 
    0.092722105882039, -0.0232561925283065, 0.111180985429292, 
    0.101642467969104, 0.0698962651574341, 0.0298123744547241, 
    0.128993888227404, -0.000604166052591523, 0.102007342088587, 
    0.111559546947973, 0.00780203245885554, 0.0433008691160239, 
    0.0342540759051337, 0.0783554023075168, -0.0499311901250606, 
    0.116807585607634, 0.121994589221166, 0.0538417932418814, 
    -0.00223110465193313, 0.0952716577554077, 0.0835477409542572, 
    -0.0178281963412341, 0.102475546428584, -0.0116533794573943, 
    0.09665230606368, 0.0347932326356882, 0.0802537351158717, 
    -0.0204693075196709, 0.0939050851389866, 0.128637855066544, 
    -0.0125706400411224, 0.0706205978136581, 0.0727442639831008, 
    0.0107934293153201, 0.00545009439236518, 0.0192767847881693, 
    0.0725788469167361, -0.0381028337996461, 0.108326697259131, 
    0.0624030098323537, 0.0696159701036483, -0.0442621325056721, 
    0.0552963846606241, 0.103210539584627, -0.0678037567254975, 
    0.0808416595338951, -0.00018693167126744, 0.0684701242266515, 
    -0.0255572282703349, 0.077112813712523, -0.0374030290712949, 
    0.10678419908946, 0.0992516414649681, 0.00363567702183817, 
    0.0333273659629242, 0.0554763492640275, 0.0253988998308493, 
    -0.0517341368790674, 0.0364670773981621, 0.066252016964961, 
    -0.0185635118402146, 0.101704638793362, -0.0248685907600982, 
    0.0858725399314155, -0.0693049736738438, 0.00838791616506327, 
    0.0860106737604705, 0.107374444164242, -0.0841665963832202, 
    0.0246838444778607, 0.00597833091820916, 0.0174409575256176, 
    -0.0494638188142967, 0.0445671777660303, -0.0248812387940585, 
    0.104455280592316, 0.0165198890186579, 0.0355423016822048, 
    -0.00650547952874952, 0.045477627157746, 0.0423810147731437, 
    -0.102982140364029, 0.0698059483584625, 0.0338820853936287, 
    -0.00328722759841097, 0.0842490969674024, -0.0912586370728233, 
    0.0717416827117808, -0.0626564658358226, -0.0139205329274623, 
    0.102024281761601, 0.0707996807262948, -0.0607619794721959, 
    0.00450824629702369, 0.0133912711318233, -0.056965925867107, 
    -0.037702806020758, 0.0112327361138424, -0.00497077206621099, 
    0.0996647870797813, -0.0767226391545804, 0.0630625857010647, 
    -0.0323922239023602, 0.0155579000275313, 0.0846486071569211, 
    0.0435322253035826, -0.108635471578698, 0.0985959463681969, 
    -0.025731773713639, 0.00332128963856508, 0.0475405366662102, 
    -0.115615911418036, 0.0149101644382705, -0.0396505750014735, 
    -0.00210333182667908, 0.100022756459037, -0.0136177463482409, 
    -0.0201029018887253, -0.00358610859118761, 0.0136631109942027, 
    -0.110970955857168, -0.00605185158718265, -0.0286444293620107, 
    0.00750840952516901, 0.0959821830999605, -0.132641335098517, 
    0.06298623811529, -0.0298397049005585, -0.00537449433660488, 
    0.0951674252428595, 0.018106848121067, -0.0792451196308446, 
    0.114028835236396, -0.0559131651070079, 0.000595148292594888, 
    -0.0199371283388362, -0.106797953838638, -0.0386191477847312, 
    -0.01921038100353, 0.0168437172635215, 0.0947236903355487, 
    -0.0966621444570293, 0.0232826842943154, -0.0323285188029712, 
    0.0792179167180163, -0.000593412502952617, -0.120509249241042, 
    0.0330441558520932, -0.0832180041052082, 0.00913035728870973, 
    0.0772714205134165, -0.149839356606014, 0.0300702533666021, 
    -0.0134126928839544, -0.000356342577619573, 0.0978580100251466, 
    -0.0215495581372432, -0.0378084744410209, 0.118948256285199, 
    -0.0696250078135141, -0.020132034595007, -0.0920200211174289, 
    -0.0755754901840457, -0.0617832674176476, -0.0082448131797074, 
    0.0281820399107155, 0.0917229771544796, -0.141141435923241, 
    0.052898168626909, -0.0501686135603817, 0.0885024365589548, 
    -0.0174398961359628, -0.0847719858104608, 0.0726743128981258, 
    -0.112633781931468, -0.00420115777186618, 0.0280560826871983, 
    -0.145154711285577, -0.00297471132505095, -0.00113081167338062, 
    0.0192091034444122, 0.0996732542591797, -0.0604005893676802, 
    0.0103358102952802, 0.106908632166106, -0.0980314798480189, 
    0.0623522503378745, -0.0518351007606106, -0.130952799256048, 
    -0.0315363534066212, -0.068658644040785, -0.00697505909501681, 
    0.0264809640761371, 0.0822985456045732, -0.158431702104869, 
    0.0561379900545804, -0.0419474697197503, 0.0894134188488235, 
    -0.0342728867203216, -0.0258395866349808, 0.103004955530429, 
    -0.117713265752617, -0.0392898394808664, -0.0453391773200696, 
    -0.115163598062492, -0.00624884322585139, 0.000408467964080562, 
    0.0367543396408667, 0.104257208974249, -0.0946714204203439, 
    0.0527297527913762, 0.0743853067001904, -0.120805484520764, 
    0.0794003242059902, -0.0685267168990564, -0.0974377494340046, 
    0.016168760487016, -0.0715763975854615, -0.0223888650071105, 
    0.00629378217995475, 0.0636053161403077, -0.163793049004419, 
    0.0469670193777119, -0.0195146785248184, 0.0922093754251162, 
    -0.049388747738115, 0.0261522337888257, 0.107051405362539, 
    -0.129116760055976, 0.049997332955198, -0.0849970746530434, 
    -0.102155786594791, -0.0683344067226991, 0.00807944073251035, 
    -0.00337161625831396, 0.0345882676473976, 0.0975331125345463, 
    -0.120606784798548, 0.0761886290318041, 0.0379444718021573, 
    -0.108087264599745, 0.0896494916383328, -0.0719474017295393, 
    -0.0272276508158435, 0.05252394840721, -0.0706531441372358, 
    -0.058752187272056, -0.037192866461458, 0.0237160171673353, 
    -0.139524523533831, 0.057831728820364, -0.00117513444715126, 
    0.107372352749523, -0.0682652521016206, 0.0655106513106432, 
    0.0764003145096563, -0.15329797484725, 0.0812592182590743, 
    -0.10513238311413, -0.0799523153144732, -0.024081462487053, 
    0.012043033654681, -0.0228001189376777, 0.0130806019138432, 
    0.0918964854872866, -0.138318020259272, 0.0826505617359634, 
    0.0152017672757655, -0.078155205008063, 0.0930398455847361, 
    -0.0673138111755421, 0.0283341013662697, 0.0640268564507554, 
    -0.0772359807290864, 0.0490377472432925, -0.0679020916316471, 
    -0.0912083798249367, -0.0274139758819804, -0.0881443470654018, 
    0.0798887817236574, -0.00134811840905976, 0.113291793453048, 
    -0.0915052258633234, 0.0918037601567904, 0.0399356335695772, 
    -0.144510066332566, 0.0954008295265828, -0.0966905957684143, 
    -0.0105090566601171, 0.0116198936729656, 0.00351330469126734, 
    -0.0598716410648921, -0.0233721229050675, 0.0856283775505911, 
    -0.136569452446415, 0.096987562005832, 0.00905332259121438, 
    -0.0600272868082408, 0.103092096860641, -0.0655618527797858, 
    0.0602530836353303, 0.0453689450291433, -0.103083596219196, 
    0.0842523460128031, -0.0482715505335043, -0.11397566232478, 
    -0.0167036529461182, -0.0413705554441875, 0.0833602304253528, 
    -0.0188496830365837, 0.106879750384306, -0.110557251276827, 
    0.103182179190992, 0.00977515519861518, -0.114662008298375, 
    0.100881544880542, -0.079744027335155, 0.0340717863688288, 
    0.0284235115896701, -0.0158322005565122, 0.0420757679898386, 
    -0.0742818203153039, -0.0632551137678942, 0.0639428962991272, 
    -0.100051739596406, 0.117496711447061, -0.0073432497422872, 
    -0.0564177031088453, 0.112669324537382, -0.0803666907776648, 
    0.077114556353783, 0.0187198855879233, -0.132855668008047, 
    0.0950042682326049, -0.0281646564010656, -0.0994237584189222, 
    0.0382453265770801, -0.0135259522426145, 0.0650392734462068, 
    -0.0398309889465307, 0.104841131749822, -0.117589518719626, 
    0.113206321266748, -0.00227770431742747, -0.0981133167912728, 
    0.0982347631451108, -0.0754335521313718, 0.0518690267202933, 
    0.0142529952401312, -0.0547255773862383, 0.0752263427131694, 
    -0.0591847023449188, -0.0895927841215088, 0.0538868717163064, 
    -0.0618512533696874, 0.117555804118673, -0.0377070412476621, 
    -0.0638688705831922, 0.106981276317816, -0.0988117484674845, 
    0.0835091584772625, -0.0103281435162814, -0.141631822573037, 
    0.101452596637041, -0.016422661719806, -0.0825500043218892, 
    0.0613090597891735, -0.000704843791443539, 0.0343347509875874, 
    0.038882747789301, -0.0548231163898809, 0.0996813985527662, 
    -0.090632295414521, 0.117901256595734, -0.0184767280005035, 
    -0.0963850540367854, 0.0998536291965039, -0.0863650132511894, 
    0.0601805357609448, -0.00319496790158467, -0.108796040324855, 
    0.0879696769171965, -0.0363534937906653, -0.081538017763848, 
    0.0673812273642971, -0.0430276542269201, 0.0931421932775464, 
    -0.0675094613402417, -0.0682203807602702, 0.107152004257099, 
    -0.108487390092754, 0.0862617459849318, -0.0181153702072858, 
    -0.130180324169167, 0.1031321262578, -0.0805395293163267, 
    0.055301822788147, -7.54264524629898e-05, -0.0115452076340512, 
    0.0541932409027647, -0.0720560271774864, 0.0777546376499775, 
    -0.0614512627164843, 0.111949218620945, -0.0355870235949172, 
    -0.0972878042154306, 0.100382186170154, -0.0988070453567965, 
    0.0639239237164491, -0.0197184817350712, -0.140009877872421, 
    0.0946652477975953, -0.0161039210940115, -0.0793081605891699, 
    0.0575883728399246, -0.0385876167201306, 0.0584292404508914, 
    0.0467819313151402, -0.0696610154328736, -0.06098986896913, 
    0.098426709618349, -0.0807779466155611, 0.0837320951048754, 
    -0.0178368707185857, -0.130627689595397, 0.097710021830818, 
    -0.0844458585383786, 0.04883994751507, -0.00746801624693884, 
    -0.073206753009286, 0.0716678804022971, -0.0710044712161665, 
    0.0612228987125767, -0.0589691853789323, 0.0935516758045084, 
    -0.0407239051509154, -0.0869433552805695, 0.0938021596223428, 
    -0.100759802939963, 0.0605128382555677, -0.0213042148575401, 
    -0.129263796429363, 0.0999932001699246, -0.0834881288831042, 
    0.0292195240266155, -0.0288668534610604, 0.016315702263604, 
    0.0501791181008257, -0.0593815828981834, -0.0563540328818078, 
    0.0781776637225016, -0.0689517145102897, 0.0753916979458979, 
    -0.0221955731664216, -0.122084322471166, 0.0939328190246347, 
    -0.0929538906952606, 0.0357471894882437, -0.0170789577049325, 
    -0.117902232534009, 0.0702174918277882, -0.0679109846539994, 
    0.0277234671243106, -0.0571825069055201, 0.0647711793252178, 
    0.0471221637329422, -0.0484650815191272, -0.0676507812575583, 
    0.0822054924807893, -0.0854962988234378, 0.0461120173966219, 
    -0.0141348791962477, -0.127565813484849, 0.0880215289646467, 
    -0.0794785208299254, -0.00404848224278003, -0.0224532383244457, 
    -0.033582065134644, 0.0710892868734594, -0.0320187054848985, 
    -0.0557300081127952, 0.0495990686634641, -0.0603378767062658, 
    0.0639586201989086, -0.0274951471911681, -0.0971165725402389, 
    0.0864827124825935, -0.0990706028453071, 0.00301178736756383, 
    -0.0112897607461152, -0.121870115914346, 0.0676537751777758, 
    -0.0691584809525931, -0.0180574780441316, -0.0504494338686029, 
    0.0290232597409756, 0.0568007850835576, -0.0452202974652739, 
    -0.0555390630230399, 0.0658232336121005, -0.0713494269655717, 
    0.0287269966138032, -0.0178677293712717, -0.120734706243175, 
    0.0796368336661697, -0.0812481634273068, -0.0470465920437626, 
    -0.0252082908578882, -0.0759192450565389, 0.0624877004789215, 
    -0.0471202659292922, 0.00241460655329929, -0.05436107170805, 
    0.0475060964984618, 0.049155117061932, -0.0433823815874364, 
    -0.0714158624335992, 0.0725646676603902, -0.0847077923030464, 
    -0.0465615989984817, -0.00891814215461339, -0.119396276007421, 
    0.0514203379057391, -0.0721383778560756, -0.0657498570976876, 
    -0.0446106021925089, 0.000998335283152322, 0.0731132890738868, 
    -0.0500095719025967, 0.03533333063488, -0.0615754504530556, 
    0.0171728208179039, -0.0974028191340982, 0.0728148638507482, 
    -0.0836646178787266, -0.105419377532353, -0.0296417320699298, 
    -0.0971177434337545, 0.0581718174676768, -0.0519021627863438, 
    -0.0529135656094993, -0.0561397027805151, 0.0210016687283105, 
    0.0702745378302381, -0.0604218868349775, -0.0597673345504333, 
    0.0584605154721147, -0.0698576167134751, -0.0883847401850046, 
    -0.026114279660936, -0.115474513852705, 0.0369261170935275, 
    -0.0660558874035855, -0.112903544496319, -0.0202023639042873, 
    0.0692794250548379, -0.0286197640227546, -0.0148408481284833, 
    0.00962863314258625, 0.0485884482531583, -0.073561513229887, 
    0.0592605827278156, -0.0708913365898888, -0.177398887253272, 
    -0.04466883814688, -0.102354719877034, 0.0407376483449258, 
    -0.0672103319938835, -0.0999895441768355, -0.0537403219592171, 
    -0.00446042609225242, 0.0787942102276466, -0.028941707658732, 
    0.0268263748814491, -0.0608172479901501, -0.104129910785735, 
    -0.0966964986321902, 0.0286303909145993, -0.0662130743191086, 
    -0.157127518044712, -0.0423423108847106, 0.0507253175458165, 
    -0.044753975758949, -0.0636217309852746, -0.00240951911272704, 
    0.0855866983578534, -0.0506182452512303, 0.0421595239260591, 
    -0.0635655752474932, -0.22946918742143, -0.0694169735011817, 
    -0.102837944660939, 0.0238795831244576, -0.0554127588133575, 
    -0.13062784318317, -0.0228574795534188, 0.0692605919687547, 
    -0.00541938326066506, -0.0181672120289473, -0.0972017906097432, 
    0.0516251344184608, -0.0751651038503324, 0.0184953020190385, 
    -0.0557232544416564, -0.21359030052173, -0.0630624050523438, 
    0.0386466295176329, -0.0648158067551656, -0.0886891288179956, 
    -0.0184723776064528, 0.0716689830161905, -0.0160001377404686, 
    0.00741837910621266, -0.236244821842444, -0.0952809374801659, 
    0.0114362001638408, -0.0424824403682042, -0.148458080119826, 
    -0.0367530222088243, 0.0460285301297086, -0.0105401528851748, 
    -0.0564297460340215, -0.0833816398333183, 0.0861159528957016, 
    -0.0426286405726109, 0.00304645002254792, -0.254511552938687, 
    -0.072340807099045, 0.0145961226634646, -0.0562848612599413, 
    -0.0926465945873809, -0.0309456372700791, 0.0586285925252524, 
    0.00822813509105014, -0.0334446166544686, -0.210622020404244, 
    0.0223381156474542, -0.0748727823747511, -0.0034816144453104, 
    -0.181344940847176, -0.0536026737647412, 0.0203659438010808, 
    -0.0409939458158773, -0.070963974982307, -0.0738789373029722, 
    0.0719947443670675, -0.00850696071887965, -0.023846236310894, 
    -0.250556127318046, -0.0809480459490109, -0.00715930707159253, 
    -0.0927509748479472, -0.0382426975014609, 0.0337337496509972, 
    -0.000968880079871908, -0.0625507709787322, -0.175470033883229, 
    0.0545249907233648, -0.045895807294083, -0.016629480297603, 
    -0.21443257686185, -0.0693713888569608, -0.00634871839575148, 
    -0.0537693868169251, -0.0765346701081802, -0.0694612799657539, 
    0.0452170708370209, 0.00357299776323336, -0.048562713961315, 
    -0.223233489900038, 0.00430553966898104, -0.0841959816486346, 
    -0.0310643008209794, -0.0986415316037823, -0.0483315126854629, 
    0.0108959778141638, -0.0293055155176645, -0.0737621184858437, 
    -0.140966216624027, 0.036741167109047, -0.0197744718909719, 
    -0.0293420850816303, -0.212136520005527, -0.0813121489861114, 
    -0.0463301065801525, -0.0802185529395972, -0.0642965682478415, 
    0.0166872222507796, -0.013841372174234, -0.0601369992560402, 
    -0.186364373012848, 0.00849603946848546, -0.0677421137951899, 
    -0.0412284223400225, -0.114875794041495, -0.0568482663280879, 
    -0.0242964958437264, -0.07719871570669, -0.115243664215599, 
    0.00472310191905038, -0.0115712843606115, -0.0409761656432697, 
    -0.190609443608362, -0.0467293865419344, -0.0797438206402577, 
    -0.0917725939168427, -0.0719568161672213, -0.0581606902707811, 
    -0.00652385570548141, -0.0768991651524869, -0.145397947025557, 
    -0.00451697650318088, -0.0489762108758736, -0.0431463428341811, 
    -0.118294150407074, -0.0595865435722586, -0.0691642884596539, 
    -0.0830576919430211, -0.105648215501015, -0.0180024311547911, 
    -0.0240003766782704, -0.0506757717732091, -0.164983927070531, 
    -0.0589526128439321, -0.0685266842221432, -0.107130688710555, 
    -0.0703274999568497, -0.0616368247855407, -0.0355385658345311, 
    -0.10321909145203, -0.121632008339662, -0.02777673853111, 
    -0.0412661567697594, -0.116458124493478, -0.0659873723402611, 
    -0.0685544950723135, -0.11814069509236, -0.0771634723213212, 
    -0.106915782891667, -0.0284933799125728, -0.0751518495933785, 
    -0.134390661588795, -0.0660228069832166, -0.0931866385018214, 
    -0.0781160717166113, -0.0616333454700405, -0.0839883739528231, 
    -0.12157475591958, -0.111601039474173, -0.0287694599715194, 
    -0.0472555736311969, -0.116129785316904, -0.0790971532248794, 
    -0.0594065615661515, -0.138569436023201, -0.0690696687051764, 
    -0.10343472067597, -0.0523152537949102, -0.115790552324815, 
    -0.120332741171116, -0.048661987642672, -0.070249105453187, 
    -0.0959554707423409, -0.0770762723828444, -0.0617121217887702, 
    -0.125797770393068, -0.131678443348544, -0.111370441670322, 
    -0.0329942275407319, -0.0795516791307446, -0.114759480734393, 
    -0.0833549548906338, -0.123482157916158, -0.0722690352088606, 
    -0.103332509266051, -0.0729293689649989, -0.147164935116262, 
    -0.112455539453923, -0.0269197057121412, -0.0615889676676278, 
    -0.109567357185855, -0.0869028647812218, -0.132594312348862, 
    -0.12055598167781, -0.114823044620836, -0.047529676557275, 
    -0.123999030874346, -0.121556947016169, -0.0615328180999083, 
    -0.0915542455703512, -0.0944064708449855, -0.0843811697512578, 
    -0.0816150974661932, -0.0833094184082009, -0.164902528380925, 
    -0.118359451823174, -0.0235432677017272, -0.0821892839983752, 
    -0.118247534137535, -0.093048555822593, -0.119643142198511, 
    -0.101583763716577, -0.0977330927997297, -0.0487457616437401, 
    -0.160454095902174, -0.129966197665839, -0.033458246133501, 
    -0.0747819627887568, -0.120114292594215, -0.0860319320896763, 
    -0.0815800399887233, -0.154042018401978, -0.102979461625567, 
    -0.018593628455446, -0.113655648936784, -0.119943718300179, 
    -0.0812954855194982, -0.0947526715398392, -0.11030784720067, 
    -0.0899469336960528, -0.0817177138189489, -0.0515963812181258, 
    -0.185407301879831, -0.122673872935495, -0.02309448178553, 
    -0.0796944830107206, -0.129865843544102, -0.0860891345178842, 
    -0.0727334250620392, -0.124899309956397, -0.0800275450607268, 
    -0.0080786125604891, -0.142257072838303, -0.131489542901961, 
    -0.0561786626988965, -0.0763604595925617, -0.138138116330798, 
    -0.0910519397492107, -0.0518114248058734, -0.181455608326627, 
    -0.087701536757687, -0.00762451085005495, -0.0935848582530283, 
    -0.123147571352191, -0.0829120682453386, -0.059206245874289, 
    -0.126799969377717, -0.0797145046500251, -0.00672650083834889, 
    -0.170728923950696, -0.121482751448679, -0.0316265072923497, 
    -0.0721822385341799, -0.148945227205642, -0.0786013979737313, 
    -0.0453823734775342, -0.150393775268043, 0.00371695004835826, 
    -0.110440370359635, -0.127400046621398, -0.0670101549812856, 
    -0.0553000443867498, -0.145805414323849, -0.0772166295013328, 
    -0.0175564256223142, -0.183674417825194, -0.0901429575770885, 
    -0.0067046277687526, -0.0755604418516661, -0.136316234224547, 
    -0.0691629063441363, -0.0374645789112584, -0.145512922830341, 
    -0.0712456048740546, 0.00720251591130018, -0.134907207205141, 
    -0.110763915962886, -0.0355528684188532, -0.0584979163483695, 
    -0.151701681813, -0.0639508349273413, -0.0181398730537901, 
    -0.16723203844872, -0.0660847914647359, 0.00343507249413638, 
    -0.0808170043780327, -0.117818863211862, -0.0525665254641549, 
    -0.043335517941283, -0.152655595450625, -0.0666264404748049, 
    -0.0061113244548608, -0.152794405716567, -0.0864891980280015, 
    -0.017579844008748, -0.0642042348539831, -0.136286345908191, 
    -0.0512288737966953, -0.0046632504781691, -0.159039566070318, 
    -0.0691569413759354, 0.00631689726863078, -0.0926124888798442, 
    -0.0775959239836538, -0.0293373426971533, -0.0601698400263351, 
    -0.158596276854665, -0.0546424594318017, -0.00692417276248846, 
    -0.149979350226192, -0.0697356304010354, -0.0106856414032948, 
    -0.0662078637314108, -0.106043771225692, -0.0383139468352047, 
    -0.0206967125785033, -0.150200664227624, -0.0615865740414356, 
    -0.00256998031825643, -0.106512164946063, -0.0209992627914822, 
    -0.0785868849816325, -0.136719516666095, -0.0440372700294277, 
    0.00195788430707247, -0.143721107371728, -0.0824851985624221, 
    -0.00719485388121289, -0.0688088015891233, -0.0660575174983281, 
    -0.0298121019626891, -0.0573614336585698, -0.146376654691869, 
    -0.0376184957600994, -0.00531934140319545, -0.110546687577191, 
    -0.0157865953394416, -0.0876615505143955, -0.108446203457838, 
    -0.0342659172284472, -0.0204371324975355, -0.13527017425524, 
    -0.0704703681577744, -0.00570347515536104, -0.0726004287833786, 
    -0.0261373692468077, -0.0941843951430659, -0.114530968570904, 
    -0.0173615388047911, -0.0147449253733534, -0.112909402192687, 
    -0.107250141929512, -0.0100504490786688, -0.0923639734549284, 
    -0.0638305683854409, -0.0300590190664406, -0.0575743750786816, 
    -0.123127747119445, -0.0441567135353028, -0.017069035264992, 
    -0.0787557992391475, -0.0233346363993694, -0.118181828221787, 
    -0.078509226304443, -0.0038528231602728, -0.0460009209386752, 
    -0.115116058248563, -0.0917894473478705, -0.00799657118194728, 
    -0.0888161668418773, -0.0255175403521269, -0.0975487611309868, 
    -0.090089120593266, -0.00332793945662242, -0.0463225274618994, 
    -0.0886372513362693, -0.0229896126396798, -0.118311159161342, 
    -0.035335705815576, -0.0133107742662127, -0.0828359871089737, 
    -0.106221273681862, -0.06405012795722, -0.021094705556474, 
    -0.0910675466873319, -0.0222481583889004, -0.124198672581914, 
    -0.0523653698179179, 0.00794480824257027, -0.0858296821957193, 
    -0.106579746942155, -0.0240166394733687, -0.108247182239625, 
    -0.0143496708127994, -0.0208894438797259, -0.116465361388034, 
    -0.0850255967082617, -0.0240889508511212, -0.0456770095624535, 
    -0.102931076408132, -0.0261275757700173, -0.124380409995597, 
    -0.0224561678758475, -0.00763584371972824, -0.125449036170306, 
    -0.114328644293948, -0.0324756699666607, -0.10581279821108, 
    -0.0205667936323163, -0.135644125049587, -0.0549787636872544, 
    -0.0226548172530696, -0.0838652815927264, -0.118526302303537, 
    -0.0318853958620668, -0.11528410885695, -0.0136748203442643, 
    -0.0187325873263117, -0.151580935415471, -0.105982656763789, 
    -0.0450475672687301, -0.112102237087257, -0.0231815925350353, 
    -0.134561542350225, -0.0340176727589627, -0.040715298063698, 
    -0.123615739128038, -0.129287427031865, -0.0387271351975653, 
    -0.106417597997201, -0.0171479283039326, -0.16094056649679, 
    -0.0883503848247964, -0.0674401174976842, -0.125291749517164, 
    -0.0318506194346686, -0.12279929558222, -0.0223014390312272, 
    -0.0442899900027966, -0.146914695246012, -0.121811044534296, 
    -0.0454312048481193, -0.107977299124889, -0.0233189563377509, 
    -0.150949056319115, -0.0693169884819871, -0.0907569924702268, 
    -0.131632165232603, -0.0352657693911014, -0.10711780653596, 
    -0.0338564997326372, -0.158442815197162, -0.107430116736109, 
    -0.056723519445573, -0.121427318371351, -0.0360043462976593, 
    -0.127615670890678, -0.0429715750369861, -0.112649460680275, 
    -0.13227368593517, -0.0386121511630419, -0.100752123510935, 
    -0.0339433999027049, -0.150347158443115, -0.0866829671001953, 
    -0.066459415049434, -0.129259946713764, -0.0392694574740972, 
    -0.098271093666532, -0.133314548556849, -0.124298253466755, 
    -0.0376942060289133, -0.118125857679452, -0.0572592383130539, 
    -0.128571793498194, -0.0607270612521056, -0.0884023966501706, 
    -0.128108516062197, -0.0388579301811208, -0.0865127764671347, 
    -0.136090593929539, -0.110788910752139, -0.0427905839288076, 
    -0.129403019806408, -0.0619291376449233, -0.0953130212900996, 
    -0.0399343349172051, -0.114956697493158, -0.117123900608121, 
    -0.0322171813601825, -0.106532029036017, -0.120175212810113, 
    -0.0847385908553114, -0.0756682093327001, -0.119760112275382, 
    -0.0562841099996622, -0.0823756173333665, -0.122467968121448, 
    -0.103067510348074, -0.0482217929536198, -0.12719352223715, 
    -0.0973590697640976, -0.0573688040756423, -0.107224236207367, 
    -0.0989040584908761, -0.0594503284664634, -0.101969284866044, 
    -0.11436693353483, -0.0745321973470854, -0.0906759375100115, 
    -0.126059417473664, -0.0963401713170288, -0.120864015328548, 
    -0.0808951415363263, -0.0832435069128563, -0.130209587492044, 
    -0.105970372879682, -0.0549269064065682, -0.125495229039548, 
    -0.103494056207457, -0.12015298838768, -0.133251529983318, 
    -0.0609956949755351, -0.110205034318651, -0.141828165434087, 
    -0.116933911441031, -0.149691049920651, -0.088224184480054, 
    -0.150193685792328, -0.150207051832446, -0.0607053792120137, 
    -0.126111853872532, -0.130711494917362, -0.139930309361984, 
    -0.172408875072853, -0.0840639722715747, -0.172157076538539, 
    -0.168563201339481, -0.141221418865046, -0.121035912618589, 
    -0.162460816383308, -0.188556391985054, -0.0892545594363845, 
    -0.159974521731953, -0.177184076062594, -0.166206147034097, 
    -0.112772539225609, -0.1770777439579, -0.193311711965471, 
    -0.14144049394208, -0.171011797197771, -0.181203762566385, 
    -0.105571440218385, -0.162893015151454, -0.190658446591471, 
    -0.133652518664192, -0.174371940985965, -0.182485332561959, 
    -0.10714066183861, -0.13889280906947, -0.183194026285502, 
    -0.122250462402696, -0.161125227583134, -0.176900616333244, 
    -0.126456816288834, -0.177055524323979, -0.108647697571604, 
    -0.137300223540572, -0.182668662351974, -0.117345976231731, 
    -0.162922320049961, -0.112802521837803, -0.17615036093817, 
    -0.103578027958075, -0.133972855541055, -0.0942009657626699, 
    -0.163067773865395, -0.0990325559268591, -0.124992684298091, 
    -0.0796279562724039, -0.088522796750679, -0.0823010938213834, 
    -0.0674849836486844 ;

 TLmodel_value = 0.0129475642349784, 0.0165106193302022, 0.0161768567059391, 
    0.00845917687262774, 0.00144598492044247, -0.00469607053658981, 
    -0.00917732737347004, -0.0114499794423909, -0.0108945254029229, 
    -0.00607913591930449, 0.00609682899330494, 0.0164196435446741, 
    0.0144586597746764, 0.00544364551715459, 0.0025746753963991, 
    0.00102657982486913, -0.00388666830755281, -0.0118299315240441, 
    -0.0321130984827399, -0.0471315622270155, -0.0467607830690525, 
    -0.0243162941450984, -0.0134499592145687, -0.00227827395656476, 
    0.0106331828904705, 0.0143043622588736, 0.0155639791427242, 
    0.0284389462583469, 0.0394734150010512, 0.0384180622417093, 
    0.0313483276184332, 0.0282094708790503, 0.0221639079608819, 
    0.0135871313844931, 0.01180955702443, 0.00296814287345927, 
    -0.0323101488591805, -0.0639173716010558, -0.0633604693374221, 
    -0.0292057070964465, -0.0113021168329487, -0.00243343296301705, 
    0.0106831120191575, 0.0218212348848981, 0.0253822160196539, 
    0.0255299204943983, 0.0220204190803165, 0.0165858322243792, 
    -0.0195803463548349, -0.0573386915897607, -0.0822376159223275, 
    0.0113934671903131, 0.015355940904662, 0.0139171479143563, 
    0.00627889784083509, -0.000604904591415537, -0.00706613905505197, 
    -0.0137359687676041, -0.0178660801456575, -0.0150161367155909, 
    -0.00747577595301868, 0.0101805150282223, 0.0210278508048071, 
    0.0136894647226743, 0.00422288722913621, 0.00437679277122181, 
    0.00628277622185621, 0.00118703865843427, -0.00460542044045161, 
    -0.0202277145674083, -0.0361173477368483, -0.0256622846740962, 
    -0.00817006774081234, -0.00603653384407431, -0.00176438576021712, 
    0.00776706187556328, 0.0108711116314019, 0.0106998822490019, 
    0.0251404612870845, 0.0387207148823234, 0.0388528918093286, 
    0.030646277548389, 0.0227217910170185, 0.015668899027112, 
    0.00537186090731584, 0.0067587235057983, 0.00211480012669141, 
    -0.0341369174241706, -0.0681928601626004, -0.0727035011892246, 
    -0.045020679196785, -0.0258881810631685, -0.0119350461256297, 
    0.00640320640791954, 0.0207225975622873, 0.0264977319557334, 
    0.0251355889078181, 0.0184013873253627, 0.00802734005277219, 
    -0.033345481996041, -0.0719998709574917, -0.0856568486949365, 
    0.0054896755339862, 0.00662617835284716, 0.00417394806311234, 
    0.00148831331277004, 0.000262088851135072, -0.00549131707493167, 
    -0.0174247204994815, -0.0227894119179215, -0.0184246741307631, 
    -0.00932872854099477, 0.0104650908725008, 0.0194111037625669, 
    0.0104340857006748, 0.00105720143332508, 0.00455716560733373, 
    0.0107230934602455, 0.00823253505997562, 0.00523241174391478, 
    0.00399933865311203, -0.00145953544101036, 0.00662630906461422, 
    0.00747241649543818, -0.00129111645344601, -0.00519633237527547, 
    -0.001438332189496, 0.000532784937403445, 0.00102326215286928, 
    0.0151230867661921, 0.0318340947002881, 0.0354296970423573, 
    0.0246678378784563, 0.0163214674940486, 0.00601762804542361, 
    -0.00294933800939869, 0.000212715213975072, 0.00142387457076507, 
    -0.0268622433125145, -0.0616637798663202, -0.0772169647542412, 
    -0.056287501219951, -0.0384598863103782, -0.0196857297378154, 
    0.00500177355424871, 0.0234892020064674, 0.0300598285169891, 
    0.0236074060102819, 0.0150874585659485, 0.00114804580440952, 
    -0.03995813910791, -0.0742603146412139, -0.0862567818947053, 
    0.00342054729648047, 0.000689136088553465, -0.000901490158534073, 
    0.00250378416171495, 0.00959705088980657, 0.00851401517032946, 
    -0.00563657051940054, -0.0142184784579181, -0.0163556473468997, 
    -0.0139918944198568, 0.00216159735097226, 0.00684411490865335, 
    0.00150969055698508, -0.00360885287054375, 0.000517803416261988, 
    0.00781026290218938, 0.00635532764964073, 0.00500619192286136, 
    0.0298494058967516, 0.0397782024519963, 0.0366442755851114, 
    0.0154842412313172, -0.00281533740835945, -0.0125021688539617, 
    -0.00908987657721713, -0.00786892336599511, -0.00819265408423681, 
    -0.00179804928312419, 0.0101374229720798, 0.0151651527012644, 
    0.0148455812289559, 0.00797650918779903, 0.000946809733788834, 
    -0.00918369340951409, -0.00579927687568265, 0.00329895764806925, 
    -0.0113444913774414, -0.0429403057099898, -0.0649748040444904, 
    -0.0563049366313329, -0.0377923727686887, -0.0161098316108583, 
    0.0188702866464066, 0.0469321113707809, 0.0522582653852993, 
    0.0362640818418104, 0.0216876209181327, 0.00741035280348333, 
    -0.0288744613592103, -0.0611848599029671, -0.072549458078201, 
    0.00690378074740777, 0.00331106263654485, 0.00218885587158616, 
    0.0103902668670909, 0.0248701471854608, 0.0328303433081331, 
    0.0186992816530009, 0.00316780821848342, -0.0107077650027795, 
    -0.0218330009998784, -0.0162650250895796, -0.0123451182586948, 
    -0.007279441731772, -0.00848016791796349, -0.00460225579589807, 
    -0.00161890129704578, -0.00226376910921221, -0.00206776039026571, 
    0.0227439297081961, 0.0312466116428749, 0.026463840572868, 
    0.0124796307887811, -0.00362336209242313, -0.0169616662459044, 
    -0.0131917665854747, -0.0110331318176266, -0.0153189562444262, 
    -0.0192297557138908, -0.0209037371450497, -0.0196042265862147, 
    -0.00110171051832336, 0.00360555726840892, 0.00167329135618752, 
    -0.00407133398554366, 0.00223303395904297, 0.0179929114668549, 
    0.019005284632277, -0.0035493612073566, -0.0403245216007888, 
    -0.0406607395115849, -0.0186005481710033, 0.0126590793016348, 
    0.0516996709009925, 0.079022708658339, 0.0776345034002721, 
    0.059177412516245, 0.0419733684492932, 0.020813041924492, 
    -0.0132485340136669, -0.0420618369884418, -0.0567274317267277, 
    0.0139385349303062, 0.0152125861844874, 0.0142770456395841, 
    0.0209251775813293, 0.0336884340554715, 0.0505386534885347, 
    0.0445235798908036, 0.0204407733544533, -0.0047942004195902, 
    -0.0299153092826184, -0.0379025920598244, -0.0295845259731171, 
    -0.0146589723430579, -0.0139701545378965, -0.0104532802526894, 
    -0.0119545038238812, -0.0155649449026583, -0.0069437354941451, 
    0.00819445138564081, 0.0129445306665883, 0.013442821724944, 
    0.0118264420152162, -2.97407407590923e-05, -0.0132128535245158, 
    -0.0118054592835071, -0.0123282168873556, -0.0199776053277562, 
    -0.0364014713909701, -0.0517230830289839, -0.0469438157623515, 
    -0.0116324189606076, 0.00457114151372095, 0.00889480625226098, 
    0.0100229934331757, 0.0192196982596914, 0.0363478686238908, 
    0.0433405888538712, 0.0194556914519504, -0.0128426843947555, 
    -0.0219820778826333, 0.000467419591722578, 0.0359706613024547, 
    0.0718539850602844, 0.0904450093746605, 0.0864573641400251, 
    0.0713162306474155, 0.0587376913806232, 0.036732500104029, 
    0.00654100909525372, -0.0203342507333758, -0.0330763709869003, 
    0.0174809966307294, 0.022082798457518, 0.0216057003564381, 
    0.0222003545347801, 0.0287579729480963, 0.0446662731205526, 
    0.049335221430364, 0.0291347752159554, 0.0017760658930104, 
    -0.0307489833058034, -0.0488394606913631, -0.0376394566243601, 
    -0.0213470821745245, -0.0190567882515956, -0.0160460567263761, 
    -0.0187508457079199, -0.0248605871530846, -0.0176857259565676, 
    -0.00195399999060133, 0.0078337629317834, 0.0122166804241589, 
    0.018986811605453, 0.00883038867472392, -0.0040696418110286, 
    -0.00952943511100932, -0.0145184703139767, -0.0251495826440291, 
    -0.0500018553556066, -0.0627208794403922, -0.0631579540839228, 
    -0.0178138383468983, 0.008132407796632, 0.0173771726136723, 
    0.0258537814130639, 0.0386652092297051, 0.0491676644151231, 
    0.0515896365080913, 0.0282802793016646, -0.00365136029901438, 
    -0.0143297165476289, 0.00578486852180446, 0.0382167596008135, 
    0.0643674818121121, 0.0681689204696115, 0.0666735043837832, 
    0.0682366188496421, 0.0756842620799685, 0.0624636137966362, 
    0.0274579816501769, 0.00177952595845731, -0.0121206220935169, 
    0.0156661786846244, 0.0195364377956798, 0.0183415421299047, 
    0.0132197456854685, 0.0185370911635313, 0.0281791336905617, 
    0.0425739811920124, 0.0332483337142457, 0.00953043512780304, 
    -0.0237121583788472, -0.0456833148044823, -0.0405008869910269, 
    -0.0285420154309446, -0.0246132237420192, -0.0223101028914105, 
    -0.0229519032317453, -0.0275460693981128, -0.0266265078511888, 
    -0.00502719869789706, 0.0150127018923675, 0.0227627688922427, 
    0.0283379316978949, 0.0133505789817595, 0.000629656280393354, 
    -0.00823282752746271, -0.0165941648580893, -0.0266734849184927, 
    -0.0377055980099184, -0.050083764830983, -0.0454372254938292, 
    -0.0114247862181275, 0.0117398468587167, 0.0209712685186232, 
    0.0321948777233255, 0.0410006904637385, 0.0444039761290757, 
    0.0306306675767807, 0.0156823916525372, -0.00985073791308424, 
    -0.0211943298717324, -0.00370885210969693, 0.0197892258951295, 
    0.035460148303662, 0.0388939925656542, 0.0382820159715218, 
    0.0461259872662147, 0.0661921963656539, 0.0762979618042441, 
    0.0487804045811943, 0.023642322856848, 0.0110850182799864, 
    0.0077679080899601, 0.0095548874770872, 0.0067568305170652, 
    0.00363640302687788, 0.00246411760415615, 0.00593176899270308, 
    0.0195299313004078, 0.0288398123979618, 0.0169020892332665, 
    -0.0127294592462036, -0.0336852627325574, -0.0379690590442505, 
    -0.0341095894967337, -0.0260035053299349, -0.0237430516095076, 
    -0.0260061589920986, -0.0294346296414378, -0.0289960512112291, 
    -0.00333636935207176, 0.0244272001822777, 0.0342213865460868, 
    0.0313474742299629, 0.00972452216838793, 0.000320594742222362, 
    -0.00619364441828548, -0.012549722968987, -0.0157036384838074, 
    -0.00687997374865421, -0.0155637151455192, -0.0134817310877881, 
    0.0054443679478983, 0.0156042428045388, 0.0198745607500763, 
    0.0236944323614337, 0.0296302601409606, 0.0303595791420308, 
    0.0189983925589404, 0.00425086164860308, -0.0176848981178398, 
    -0.0297930028903017, -0.0119110042271617, 0.00753736326700449, 
    0.0240712304141433, 0.0265948472868555, 0.0233749296781071, 
    0.0287527733652359, 0.0583711745998291, 0.0838774065684794, 
    0.0655109480143792, 0.0438087320438739, 0.0280959463958211, 
    0.00341576678058371, 0.00165186047301265, 0.000194924841096012, 
    -0.00209128180034057, -0.00280018687258358, -0.00665586994273493, 
    0.000770034792562939, 0.0186604277803028, 0.0163457266847248, 
    -0.00587789932444767, -0.0264247801338803, -0.0348102868353207, 
    -0.0341129034082657, -0.0257033330503638, -0.0226893927543929, 
    -0.0305232588290687, -0.035474947602734, -0.0308694192482048, 
    0.000830829593849185, 0.026719463846752, 0.0294984432531522, 
    0.016448473342497, 0.000411429182592849, -0.00186315539538456, 
    0.000519728039219338, 0.00101207591802331, 0.00572671089928378, 
    0.0225763849020675, 0.0274946583134947, 0.0217077913708437, 
    0.0205122597331276, 0.017861680506697, 0.00920294246100966, 
    0.0046590788100754, 0.00856836943364117, 0.010611632265603, 
    0.0117870766145983, 0.00804982460453102, -0.0150912008016744, 
    -0.0319148413575637, -0.0206358700523008, 0.00151048677105144, 
    0.0289579170296473, 0.0330708819686002, 0.0246906522032379, 
    0.0280613746258453, 0.0646386419606186, 0.0948568956926085, 
    0.0890450067603364, 0.0611642504979244, 0.0447689440681106, 
    0.00342732206750792, 0.00103399153744283, -0.00162682348405858, 
    -0.00371466520358258, -0.00511389566839983, -0.0128471223898916, 
    -0.0132847878263407, 0.00212920912542506, 0.0090752555469788, 
    -0.0013394881893866, -0.0156462308362861, -0.0228594945757044, 
    -0.0272938854515062, -0.0236902376958186, -0.0227253823077305, 
    -0.0354534988967704, -0.0388472434444725, -0.0234124340896317, 
    0.00801614297508932, 0.016985456278673, 0.00184334050959993, 
    -0.013030530852634, -0.0126968815988982, -0.00382219654179556, 
    0.00862369981880025, 0.0153173547038992, 0.0246066129578836, 
    0.0391762350465296, 0.0502511753552607, 0.0418268107065593, 
    0.0251401454869841, 0.00487222298492204, -0.0125221779011577, 
    -0.0180986966434051, -0.0129184291626326, -0.00270103383321589, 
    0.0149819484050582, 0.0193455975150179, -0.00455300761310167, 
    -0.0344239798081094, -0.0231409588393211, 0.00144491127134904, 
    0.036410240988245, 0.0378996946066784, 0.0326937464236158, 
    0.0458720027053735, 0.0860076662061786, 0.101549785240418, 
    0.0981237974118425, 0.0751188360822196, 0.0552174172562245, 
    0.00677488561460013, 0.00441311932807764, 0.00237427898072263, 
    1.52147926056152e-05, -0.00331919700255158, -0.00978071102011975, 
    -0.01861538447055, -0.0115053507255251, -0.00166797234829314, 
    -0.00290694602171444, -0.00831182858979115, -0.0107287628676275, 
    -0.0185409086333165, -0.0210094954855366, -0.0213506639937833, 
    -0.0278241262728567, -0.0247647573017312, -0.00884045730793848, 
    0.01184156368982, 0.00589692336190713, -0.0211836083336722, 
    -0.0316386133197963, -0.0187593900762189, -0.00498316056659306, 
    0.012441627872324, 0.0230236856418895, 0.0340986513915854, 
    0.0485065835230453, 0.0570361182878994, 0.0465481470370859, 
    0.0254950133313216, -0.00664649174245908, -0.0320090096206743, 
    -0.0370304863102454, -0.0307726679677585, -0.0124217451615055, 
    0.0182044475074968, 0.0259105116262974, 0.0048035972723017, 
    -0.0284124944393514, -0.0266037364318178, 0.000567218165616576, 
    0.0356067655854343, 0.0359650226339578, 0.0342446822924646, 
    0.0536679259872257, 0.0922724268565685, 0.112404533649337, 
    0.111057722347146, 0.0856071483846581, 0.0572235524305314, 
    0.00927826260248465, 0.00756911786295374, 0.00732652991274956, 
    0.00662673433084101, 0.00386335830078685, -0.000682123550826679, 
    -0.0123904980504654, -0.0121224179816383, -0.0040896903341683, 
    -0.00574794412110401, -0.00920299560546909, -0.0080656977883036, 
    -0.0140536200328477, -0.0174341344907934, -0.0192207827458868, 
    -0.0186663097410512, -0.0116842561176318, 0.00244952302029464, 
    0.0137549556104625, 0.00385345799183273, -0.016610487780556, 
    -0.0257413737211912, -0.0180822730612188, -0.00645602448645957, 
    0.010498653920577, 0.0223862794123551, 0.0325122298193509, 
    0.0491434889885665, 0.0571517672104694, 0.0589940473135955, 
    0.0218722936564283, -0.0225599734083633, -0.0580274667483809, 
    -0.0568419360116015, -0.0451177581260463, -0.0246238257579327, 
    0.00761307577497902, 0.0219885998932487, 0.0079887382983331, 
    -0.0189967222446323, -0.0191256065328361, 0.00109123350456461, 
    0.0258052735916922, 0.0226577763639221, 0.0213614806947424, 
    0.0418435278764544, 0.0755731603681277, 0.10757470080091, 
    0.110950357437125, 0.0860841072380247, 0.0551428056772616, 
    0.00939197461526537, 0.0071867287861017, 0.00836455189069008, 
    0.0104407036703558, 0.0110145148187988, 0.00864657631031133, 
    0.000551289186455307, 0.000400303804255862, 0.00664631072113169, 
    -0.00339674523298617, -0.0118827246165604, -0.00903832029125476, 
    -0.0102522866624849, -0.0117661605262872, -0.0153409258723349, 
    -0.0112696455106733, -0.00182350301069976, 0.00917116954077375, 
    0.0149553159188111, 0.0105898708856217, -0.00027063449196999, 
    -0.0141046045307703, -0.0174211542038801, -0.0060472879532331, 
    0.0120240799658134, 0.0200207969330159, 0.0276326980442932, 
    0.0383884234293313, 0.0464801492779009, 0.0479835081189202, 
    0.006998045405824, -0.045829026696483, -0.0879102287425313, 
    -0.0766692524255371, -0.0530607321650727, -0.0353901254149816, 
    -0.0128976673979652, -0.0113207695884555, -0.00289411089920606, 
    -0.0104545777567101, -0.00328237254867517, 0.0120715922204359, 
    0.0206150775846053, 0.0109944643712079, 0.00558230569041869, 
    0.0152514166012042, 0.0391168115736485, 0.0755388345799455, 
    0.0799626573763194, 0.067758394582155, 0.0430255651178998, 
    0.00454392040317296, 0.00275826909927398, 0.00281989349254602, 
    0.00212700603923236, 0.00364917935896708, 0.00717381124793255, 
    0.0116229579339459, 0.0167112558065219, 0.014952592735314, 
    -0.0138649383171576, -0.0283688899950972, -0.0193511823155518, 
    -0.0103635735202721, -0.00831835936175077, -0.0130967586041787, 
    -0.0107598736417642, 0.00079581485040214, 0.00760348321275486, 
    0.0146971554125201, 0.0181689068248266, 0.0107688865236787, 
    -0.00436239063091574, -0.0116912578775114, 0.000393211383661423, 
    0.0202017052683624, 0.0276877365534301, 0.0305257661249348, 
    0.0356545971859727, 0.0379231645731615, 0.035746053173377, 
    0.00092016257595778, -0.0433782484425901, -0.0792170417597627, 
    -0.068541018436788, -0.0506655270571042, -0.0379813458154999, 
    -0.0228178211712242, -0.019722218755358, -0.0136284934733308, 
    -0.00649281113656411, 0.00677963648640252, 0.0180507160139386, 
    -0.00609387326324608, -0.00793241677931823, -0.0051855433301815, 
    0.0132286256709435, 0.0370224907457541, 0.0601860638409389, 
    0.0368914567162854, -0.00278452250376164, -0.00274494904950311, 
    -0.00700523366433968, -0.0178697924529044, -0.0169736089722471, 
    -0.00265897578575876, 0.0127226665013669, 0.0201368009750786, 
    0.00381583574293082, -0.0377617453819132, -0.0475894764540773, 
    -0.0325209343627915, -0.0115768814481605, -0.00779136950093378, 
    -0.014685188034544, -0.0138652638634822, -0.00271996410488367, 
    0.0054054761391755, 0.0141332889476985, 0.0215592843673409, 
    0.0218389878681583, 0.010535868767885, 0.00343303666334622, 
    0.016378228389484, 0.0442572688321298, 0.0510350346564511, 
    0.0472654954159503, 0.0361933748152626, 0.0240176499806231, 
    0.0210940202834524, 0.00806230957306808, -0.0201072092569833, 
    -0.0418428529326409, -0.0388138547230306, -0.0239395254982172, 
    -0.0278629284503907, -0.0265319863574192, -0.027157958632166, 
    -0.016289348614159, -0.00738967643138168, 0.0121307211374826, 
    0.0186036743982244, 0.013282733251013, -0.00963567459259185, 
    -0.0175549084524954, -0.00940443884195132, -0.00151869729013109, 
    0.0109939548279927, 0.0122267789719302, 0.01182048927752, 
    0.00895239802806643, -0.0090643025820144, -0.00954595923902699, 
    -0.0218673104349321, -0.0434186819232165, -0.0400585796249053, 
    -0.0142197910619512, 0.00531460300511545, 0.00873363127697917, 
    -0.0117775333537237, -0.044462601164239, -0.0485144196482305, 
    -0.0292546787750713, -0.00559134308725506, -0.00213715403222542, 
    -0.0126502965431546, -0.0147295990272761, -0.00234850194716764, 
    0.0095800317270368, 0.0163544160515713, 0.0191182928801126, 
    0.023818489831417, 0.0296340361417287, 0.0364361747779065, 
    0.0523195706665105, 0.071070015054514, 0.0767725252069561, 
    0.06840711203447, 0.0302985907546373, 0.00962658448230681, 
    0.0143572949828874, 0.0182339842957475, 0.013130381365081, 
    0.0105638090143531, 0.00338079853438689, 0.0030092238207926, 
    -0.014496428194804, -0.0233149821177287, -0.0261728313893102, 
    -0.00852640353345037, 0.00504200979092365, -0.00421338889576795, 
    -0.0110505689819442, -0.0112008519156178, -0.00609374829826195, 
    -0.00413588496108117, -0.0129270001737714, -0.00692283608756185, 
    -0.00189723686828405, -0.0117350831565447, -0.0144643092950683, 
    -0.0325134111701351, -0.0596030075558191, -0.0559367370747474, 
    -0.0248552532096341, -0.00450817397828003, -0.00439773779642476, 
    -0.0187819041176587, -0.0370163341072038, -0.0450744228154234, 
    -0.0277075687647239, 0.00304827441042281, 0.00374657097190649, 
    -0.0152608417677291, -0.0228852926675865, -0.0031672416788427, 
    0.01241894328768, 0.0119672806696282, 0.0109537108308761, 
    0.0259001867258172, 0.0582419838976902, 0.0825136746068513, 
    0.0967107782176967, 0.091554723754509, 0.0757407653717114, 
    0.0461162858773317, 0.0151846401186391, 0.000954759727343828, 
    0.0230012001403819, 0.0274307676053356, 0.0230847429775132, 
    0.016947472750081, 0.0128009274099821, -0.00654406294952777, 
    0.00403168842464624, -0.000202067542492662, -0.00757500011896801, 
    -0.00832719265196047, -0.00627487501260269, -0.0103399701809884, 
    -0.0254369929193115, -0.0128856892873159, -0.00460350235627259, 
    -0.00831197648676329, -0.0102100835643328, -0.0281549862559122, 
    -0.0526656040932096, -0.0492266313055939, -0.0225718076631783, 
    -0.00666584723581684, -0.00628512106762314, -0.0163976105411464, 
    -0.0312661349877236, -0.0370540493033293, -0.0193608400968764, 
    0.0128321495971356, 0.00621131959291356, -0.0245096402214147, 
    -0.0361175113300135, -0.0133953032481815, -0.0024325930788629, 
    -0.0102631217458412, -0.00896045914763105, 0.0295333868567304, 
    0.102585071811664, 0.138138109650718, 0.142774884666001, 
    0.0972409771452812, 0.0736334933224253, 0.0434526877650775, 
    0.0150954984562939, -0.00695274442093267, -0.00752480564988792, 
    -0.00606199179057258, -0.0262933352560776, -0.00357733153509448, 
    -0.00374360397247155, -0.0163195795689394, -0.0291727717871949, 
    -0.030786879185098, -0.0155101840260784, -0.0063120457900467, 
    -0.0073681903179025, -0.0161439538906936, -0.0274073898952717, 
    -0.0262791023558714, -0.0110460723881269, 0.0184210167488464, 
    0.0143173030593707, -0.026335598541838, -0.0449140550137355, 
    -0.0290087574310148, -0.0300333017584297, -0.0469819244401624, 
    -0.0324610541872787, 0.0363192576981395, 0.127161976770385, 
    0.144242852986736, 0.134995215732687, 0.0728169583083678, 
    -0.0019716878063606, -0.00177270064568241, -0.00682338151949032, 
    -0.00941143290008758, -0.0110717749315886, -0.00499745889546071, 
    -0.00394179459198725, -0.00901242200753602, -0.0217191947806298, 
    -0.038506815761424, -0.0342010817495202, -0.0182999195707425, 
    0.0131266326768534, 0.018433600416998, -0.0149088273613222, 
    -0.046737139258009, -0.0508800460697094, -0.0531839601495364, 
    -0.0762093620116106, -0.0570936133903757, 0.0288450177170538, 
    0.133141388157411, 0.148340820048303, 0.129889838799783, 
    -0.00142781455124633, -0.00273572287575957, -0.00478836581552227, 
    -0.00506124494603441, -0.00266946325524058, 0.00251404823746733, 
    0.0021735655800455, -0.00286725572782698, -0.0148247987483694, 
    -0.0376605728785272, -0.0438540956213936, -0.0295741613131737, 
    0.000764068675123319, 0.0118655554882675, -0.0092626090203999, 
    -0.0375031849003154, -0.0569605712823823, -0.0806407591036413, 
    -0.0908940527311099, -0.0580912514955728, 0.0252145056879124, 
    0.0894953088673689, 0.000745945253960938, -0.00576442907786257, 
    -0.00815881104159044, -0.0052452896188772, 0.000259072770833597, 
    0.00758423093363399, 0.0106770500797866, 0.00828454995195933, 
    -0.00263837636494345, -0.0240778046828858, -0.0342649212424141, 
    -0.0265603620264035, -0.00076730060324682, 0.00932431164883643, 
    -0.000596366915745975, -0.0234868943585065, -0.0511715789320097, 
    -0.0799725086743557, -0.0855715662134497, -0.0496033550348955, 
    0.0256449593147183, 0.0720950400587209, 0.00050890191423292, 
    -0.0119590847786956, -0.0155047813462967, -0.00789350468061827, 
    0.00351112024776804, 0.0112549928226791, 0.0137899153843699, 
    0.0108476013256521, -0.00118598771448183, -0.0142221629005227, 
    -0.0159198703464269, -0.0105467429113662, 0.00593250612221352, 
    0.019757290766183, 0.0206363183211612, 0.00303636044969429, 
    -0.0297503180244244, -0.0724298523110727, -0.0783827610565814, 
    -0.0593119332853888, -0.00493677570571337, -0.0167272222258762, 
    -0.0158023377692203, 0.0014010215945876, 0.0122294665627447, 
    0.0147015190273771, 0.00773646603758951, -0.00550492040000248, 
    -0.0149537431605031, -0.0172546714694126, -0.00806729800116563, 
    -0.00085009549917822, 0.0149776889133026, 0.0352174906014049, 
    0.0393819410274141, 0.0277956919901732, -0.00778665124592094, 
    -0.0526798445818858, -0.0744724040624448, -0.00808667350850667, 
    -0.0103860442452962, 0.00257738891390541, 0.0316581215247254, 
    0.0323814363069329, 0.0195561104449284, -0.0054082226063498, 
    -0.0283383250711675, -0.0340175783373037, -0.0345904495311634, 
    -0.0209234205265561, -0.00646392179317921, 0.0128857907842564, 
    0.035433959130579, 0.0476038980515149, 0.0406505660653753, 
    0.0193050743379639, -0.00840998406569234, -0.000335095844687841, 
    0.0243873914994291, 0.0526027827666749, 0.0528884564717381, 
    0.0263843990085549, -0.0215224115355458, -0.0475506977401109, 
    -0.054145285702014, -0.0599548680006324, -0.0535525416894684, 
    -0.0375523314868667, -0.0254953993482878, -0.0057904739666609, 
    0.0205855102778888, 0.0377833246750138, -0.0104810508865621, 
    0.000235381978712366, 0.0258155234058673, 0.0469462870482117, 
    0.048737341730788, 0.0198015219978692, -0.03801048136928, 
    -0.0668752483775189, -0.0719813683326779, -0.0873254348124654, 
    -0.0859469568857848, -0.076746150211037, -0.0762885509652407, 
    -0.0579375238451794, -0.00755094316885137, -0.0108419503650548, 
    -0.0029531094011924, 0.0117644860946516, 0.0260320385466087, 
    0.0271315331687392, 0.00135805314073312, -0.0421713371303097, 
    -0.056031388036654, -0.0738815562034517, -0.104727087985557, 
    -0.103187460284842, -0.0951367546401218, -0.0910352657936312, 
    -0.0829061194575249, -0.0136568533881305, -0.012460615370042, 
    -0.0119876221863586, -0.00408337344973318, -0.00288620730735063, 
    -0.0148949862736827, -0.0273748012940083, -0.0259652214025892, 
    -0.0475150425711092, -0.0897706640906075, -0.0916850836414507, 
    -0.0716727617411929, -0.0186666492905766, -0.0211789304240224, 
    -0.0280350567634124, -0.0221853820851215, -0.0178409811735506, 
    -0.0223986210430083, -0.0233933125904582, -0.0123344188145091, 
    -0.0364704961591103, -0.0808671880768163, -0.0833326061311759, 
    -0.0596258947066549, -0.0285254254434115, -0.0331712556844121, 
    -0.0421177710292491, -0.0392952275862906, -0.0373213362261451, 
    -0.0443366053503318, -0.0378544268884025, -0.0227055245305056, 
    -0.0432052347061433, -0.0809635153481403, -0.0843549676948581, 
    -0.0535741039670215, -0.0350458750960181, -0.0363189306358851, 
    -0.0471176444335049, -0.0532818933431255, -0.036934439850489, 
    -0.0341713151633636, -0.0326853771104198, -0.0267583602732337, 
    -0.0479415089674478, -0.0776338772137229, -0.0801923308136426, 
    -0.0322523695370024, -0.0460955751474211, -0.056537336739774, 
    -0.0472282087776092, -0.0123058831219398, 0.00620725790191012, 
    -0.000231418800773645, -0.0117986510233602, -0.0383059250262704, 
    -0.0706878352552045, -0.0694048533881801, -0.0265352905200085, 
    -0.0424830275216618, -0.0489604973892249, -0.0235756220150489, 
    0.0214731438177261, 0.0425857622170224, 0.020840907782395, 
    -0.00700993429458213, -0.023974194848949, -0.0443725629112998, 
    -0.0503401903657027, -0.016811976788888, -0.0377273139437221, 
    -0.039387961650773, -0.00484477150334412, 0.0271896948491072, 
    0.0342111799404695, 0.0091055851702194, -0.00965037994344112, 
    -0.0078552527195103, -0.00809885793103826, -0.00681389938112683, 
    -0.0276652797696658, -0.0289031824411395, -0.00240102545857706, 
    0.015841807508794, 0.0150438494444683, -0.00519697299952048, 
    -0.0118112507477169, -0.00524144042564615, -0.00331950045032903, 
    -0.0193322906953633, -0.0198816505047994, -0.00144175247711782, 
    0.00753203547190269, 0.00474381889582491, -0.00754966423526364, 
    -0.00758358892631241, -0.0048178841686109, -0.00391831179919112, 
    -0.0161789463534969, -0.0145666632905065, -0.00374686685758645, 
    0.00191174523124971, 0.00159155812788246, -0.00261530561204123, 
    -0.00237811708903899, -0.00625032216212012, -0.0188495483181722, 
    -0.0159587500417869, -0.00744179172629591, -0.000159722548936052, 
    -0.00993852200150385, -0.0176447781409628, -0.0142722707729867, 
    -0.00885558442706843, 0.00441477532871353, 0.00377461572342738, 
    0.000510099071995149, -0.00451547331490963, -0.00377271777315985, 
    -0.00205884740257123, -0.00083811089268248, -0.000977429645338066, 
    -0.00025331323824276, -1.50585506126048e-05, -8.19470932997056e-05, 
    0.000167572606011072, 0.000281230269323909, 3.60240466386104e-05, 
    5.15286063503576e-06, 4.37348396245356e-05, -4.16739086632757e-06, 
    -0.00644222245226954, -0.00143927386226674, -0.000208266855641955, 
    -0.000164338168794069, 5.58639913581871e-05, 0.000466279068392992, 
    0.000310298459049644, 0.000437308362897762, 9.76117469744712e-05, 
    -8.31928149970467e-05, 2.9798791225816e-05, -4.29699884385249e-05, 
    3.29930715674726e-05, 5.19630857432846e-05, 1.58421651755011e-05, 
    3.3216892048751e-05, 2.88855262022329e-05, -2.05290518508915e-06, 
    -7.87984179056558e-06, 0.000504406796763657, 9.01820977477984e-05, 
    -0.0107809359145911, -0.0102196094437012, -0.00642644423902163, 
    0.00321558407710288, 0.0105231188894632, 0.00953100143956294, 
    0.00366412559393877, 0.00281973010395942, 0.0018712250363919, 
    0.000682448426082365, 0.00110539397899561, 0.00139494859021734, 
    0.00124335368127894, 0.000425016947917689, 0.000477815108873476, 
    0.000267263655599067, 0.000102825233525356, 0.000211295627869387, 
    -3.62603499720598e-05, -0.000211823198183143, 0.00266897814518906, 
    0.00262268609044026, 0.00180559306444059, -0.00122181190622904, 
    -0.00299014391756674, -0.00381521536555691, -0.00209985879934873, 
    -0.00120139560886189, -0.000675602860242856, -0.000255692903440251, 
    -0.000186312502509954, -0.00026510592029442, -0.000279731978504, 
    1.0664092287454e-07, -3.54536298844296e-05, -2.27607122690693e-05, 
    -1.23142904216059e-05, -4.23014563549295e-05, -8.61219464357903e-06, 
    1.03987196373955e-05, 0.0123610609792234, 0.0164579295089536, 
    0.0158002461730109, 0.00861253678842856, 0.0023850235872657, 
    -0.00312048577532759, -0.00802315092294955, -0.0130209342182779, 
    -0.0125965016156499, -0.00749342012147224, 0.00469793464265366, 
    0.0132042305598417, 0.0140620609779031, 0.00735442241246228, 
    0.00246662642078306, 0.000826341891006821, -0.00454521552346237, 
    -0.0132968750884342, -0.0296343047445258, -0.0421589746868298, 
    -0.0509301784045145, -0.0237495177641578, -0.0170887944232747, 
    -0.00867928910376683, 0.00479025832427871, 0.0109294315758013, 
    0.0143192558872805, 0.0298333167829121, 0.0398962445853942, 
    0.0369985706744855, 0.0296572203838496, 0.0277134630409104, 
    0.0229037486616385, 0.0148234007241317, 0.0125650139202444, 
    0.000872697098399822, -0.0323970261784474, -0.0622579471022477, 
    -0.0660481992518822, -0.0345643528550157, -0.0151807470400514, 
    -0.00552981238358994, 0.0103353366116871, 0.0225974774349126, 
    0.0245783427365449, 0.0253357029411169, 0.0211504317201422, 
    0.014248603677714, -0.0189148905279399, -0.0442631861048264, 
    -0.0751977968057208, 0.0109958846445372, 0.0146123527625537, 
    0.0146012177527087, 0.00685976851316352, 0.000341382392982961, 
    -0.0043642619260276, -0.0128625885979807, -0.0189252586472544, 
    -0.0167278373865533, -0.00968348038779403, 0.00918376169536931, 
    0.0184620291426995, 0.0121870585099065, 0.00592717380813795, 
    0.00370978973184232, 0.00521083978765899, -0.000524077328250382, 
    -0.00465845836377426, -0.014757379420826, -0.0429424537824622, 
    -0.0431803370177967, -0.00815909895146293, -0.00489228895791607, 
    -0.00410015664584092, 0.00185438889224776, 0.00493540753558684, 
    0.00788100702621426, 0.0282949393202707, 0.041075334750061, 
    0.0365003173492476, 0.0288905975382237, 0.0233862745718554, 
    0.0163905747642494, 0.00545557263538707, 0.00862260622546789, 
    0.00418020670514466, -0.0284393667352405, -0.062310942835939, 
    -0.0742600704953825, -0.055274609072126, -0.0358451089166944, 
    -0.0176576737386015, 0.00718626936534111, 0.0231681277477493, 
    0.0278183274040587, 0.023366235955747, 0.0152632378837544, 
    0.00306186858377455, -0.0360390842038251, -0.0635582556430062, 
    -0.0808563006462154, 0.00565292710823213, 0.00753265194128524, 
    0.00518350847503108, 0.00186080863837397, 0.00215474992854538, 
    -0.00333618502942216, -0.015781808389591, -0.0222578386734927, 
    -0.0192857968585992, -0.0123314581411662, 0.00722223701924301, 
    0.0139398338350491, 0.00999981927421628, 0.00285984070982572, 
    0.00480549281329699, 0.00989987001273641, 0.00729943879097593, 
    0.00647113924740269, 0.00653800891732174, -0.0287951926572987, 
    -0.016233895482078, 0.00957637876613321, 0.00363090652195793, 
    -0.00415834287291656, -0.00482652455376791, -0.0032589429363557, 
    0.00292555164517655, 0.0249130093337994, 0.0372520451598647, 
    0.0327044781137124, 0.0213369391871326, 0.014844671676785, 
    0.0048920267219297, -0.00273947870027401, 0.00206622877683592, 
    0.00292847380766988, -0.0215029066096657, -0.0542440725292413, 
    -0.0744753116937512, -0.0613747077631643, -0.0438754410702999, 
    -0.0213245848919605, 0.00926905259696337, 0.0277776991505186, 
    0.033395932481381, 0.0198345733957382, 0.0115652339121589, 
    -0.0014557760680425, -0.0459612436346839, -0.0734816986879982, 
    -0.0851454846187384, 0.00403331584526618, 0.00131031258796713, 
    -0.000343728630610459, 0.0029589342985664, 0.0125664739331382, 
    0.0108318165061741, -0.00426884636926912, -0.0131587530712994, 
    -0.0164892297697963, -0.0171017901360558, -0.00431644500045416, 
    0.000461187093210636, 0.00384552412863111, -0.00117135188972983, 
    0.00205012082179993, 0.00894441597526794, 0.00611651160026452, 
    0.00965324015265905, 0.0277381310836677, 0.0277805855583376, 
    0.0332686723000725, 0.023328294639949, 0.00375456012961352, 
    -0.00935278088528122, -0.0104362982224827, -0.00875210143893252, 
    -0.00358856753293267, 0.0102619262877112, 0.0186923394716113, 
    0.0130636906509659, 0.0143586321282171, 0.00857398663763385, 
    3.49709335155808e-05, -0.0084367761829682, -0.00320780618019269, 
    0.00291187415170974, -0.0130067494033508, -0.0390030692527425, 
    -0.0615831983617025, -0.0553167934533821, -0.0308724974328158, 
    -0.0140672895172157, 0.0211193638362684, 0.0549826445895195, 
    0.0580199141960372, 0.0368274247637808, 0.0244001120918479, 
    0.00915173863721863, -0.0298543216784698, -0.0655049716603865, 
    -0.0706698050477358, 0.00771179744170651, 0.00334798847644134, 
    0.00212704069546357, 0.0102594919122599, 0.0275791981333697, 
    0.0354125371079757, 0.0180699099741378, 0.00208898715529341, 
    -0.0129256917575657, -0.0251678735050479, -0.0224557460848499, 
    -0.015185212296828, -0.0043511549988865, -0.0064441863108455, 
    -0.00332337559993836, 0.000187999614102943, -0.00247249916996956, 
    0.00582539967578795, 0.0294810686709372, 0.0268503810837738, 
    0.0216917411101316, 0.0145555722436563, 0.000519554867772509, 
    -0.0147078120303692, -0.0138886147881387, -0.0118547742510384, 
    -0.0114675448554276, -0.00988608697047365, -0.0172829839916259, 
    -0.0219860958332473, 0.000181857311775362, 0.00326726866593179, 
    -0.00038609950869961, -0.00220315457771942, 0.00878149874662831, 
    0.0231531603664387, 0.0212951192943391, 0.00831715069461479, 
    -0.0406998738799023, -0.0390875410153756, -0.0089820144362805, 
    0.0168897620179954, 0.0493674833657135, 0.0843374973714301, 
    0.0804036018550698, 0.0622456343952438, 0.0416038239481051, 
    0.0153129498615382, -0.0238796456114158, -0.057468528568815, 
    -0.0599031407887576, 0.0133609154619451, 0.0139007872957274, 
    0.0132326953486817, 0.0191021229330116, 0.03248147485629, 
    0.0498350661913423, 0.0409922334523081, 0.0153589857964073, 
    -0.00844143014164101, -0.0324014311460508, -0.0398184122488461, 
    -0.027048274078298, -0.0117976373865432, -0.0125208793777652, 
    -0.0109140442060973, -0.0119480773413055, -0.0164322827614318, 
    -0.00161128161315199, 0.0112474171598215, 0.0084328260803863, 
    0.011177160623503, 0.0138697477881088, 0.00153325705258528, 
    -0.0143175144523233, -0.0119091081074786, -0.0124876813700258, 
    -0.0184082437643194, -0.0343544315364121, -0.0565246979246205, 
    -0.0476843929198345, -0.00831468593433625, 0.00550127203636222, 
    0.00774647517091035, 0.0133373189686165, 0.0287973190163636, 
    0.044405875295672, 0.0467714655352595, 0.0253963365043625, 
    -0.0111501770331468, -0.0206131360824899, 0.00645261740964399, 
    0.041112422572392, 0.0688243193904797, 0.0902605043173049, 
    0.0828120809598148, 0.0692871959894115, 0.0541036831141722, 
    0.0274990021897954, -0.002691974902106, -0.0309114804455105, 
    -0.0372409622644815, 0.0157656657574286, 0.0206062319920304, 
    0.0202568117542539, 0.0205253630264785, 0.0262148289291302, 
    0.0422986958157145, 0.0438682931272722, 0.0236104746194913, 
    -0.00134240353465378, -0.0336290987479479, -0.0476727286169865, 
    -0.0334967684015352, -0.0183364862842753, -0.0175981555654125, 
    -0.0171253138879115, -0.0222614572448685, -0.025827729136246, 
    -0.0107740900363005, -0.00383231383618993, 0.00898124063481147, 
    0.0161737239786907, 0.0223514087299203, 0.0101496875503062, 
    -0.00592754759171167, -0.0097449415983582, -0.015805554422642, 
    -0.0265699269674958, -0.0507493850028307, -0.0567876565515128, 
    -0.0632889727174049, -0.0142230365576826, 0.00947484061354198, 
    0.0167890985605338, 0.0274802652675004, 0.0441869406152939, 
    0.0509244003261041, 0.0404169004633139, 0.0264895249230769, 
    -0.00168601651220209, -0.0154130121396848, 0.0051845124215497, 
    0.0385389239438676, 0.0674535393746199, 0.0670757016705437, 
    0.061704614151258, 0.0649343540832139, 0.0749857195059143, 
    0.050292747662834, 0.019991652040157, -0.00240028934035333, 
    -0.0149235479501055, 0.0147295148475701, 0.0161840557409246, 
    0.0180920796172721, 0.00985759643033279, 0.0163984988014882, 
    0.0264517073941991, 0.0408130398767775, 0.0298900867245962, 
    0.00586282464729472, -0.0279921165312195, -0.044672428682212, 
    -0.0368349222879272, -0.0256541018962891, -0.0225314166321884, 
    -0.0217351726463178, -0.0253043692161667, -0.0298660509587491, 
    -0.022910241039649, -0.00808205736820168, 0.0173440342902296, 
    0.0280942486567719, 0.0302516166556098, 0.0151058375679496, 
    -0.000108391564694693, -0.00979306177436712, -0.0217025187544996, 
    -0.0303389476163214, -0.0299317766318745, -0.0370036370379306, 
    -0.0303792618127551, -0.0106754897473822, 0.00841352536734229, 
    0.0196906495872737, 0.0336615009695309, 0.0419683661436667, 
    0.0386560785628011, 0.0170020847425731, 0.00723766715414559, 
    -0.00805356543284047, -0.0189150321290397, -0.00645379139208346, 
    0.0168535133698623, 0.0354768152573642, 0.0397308618549599, 
    0.0358583891768628, 0.0407392390661075, 0.0660467685154047, 
    0.0709243674124898, 0.0444248363275769, 0.0296971787280247, 
    0.0119008014471561, 0.00602293915750914, 0.00825307769635472, 
    0.00670527594819154, 0.00320638834471543, 0.00190706925515843, 
    0.00498875111110271, 0.015898381541517, 0.0262681731467029, 
    0.0125236447689897, -0.0210294703201598, -0.0373926895251342, 
    -0.036433596443501, -0.0292617844005433, -0.0242111908436477, 
    -0.0225309930498734, -0.0248703670114624, -0.0305980423439393, 
    -0.03061693035452, -0.00542215866793172, 0.0217971334796933, 
    0.032879700281965, 0.029100347889282, 0.0101951907667264, 
    0.000186825161888736, -0.0100420976512573, -0.0228101728466077, 
    -0.0234757047128734, 0.00846156060851283, -7.8756527381017e-05, 
    0.0038968842504157, 0.0100276590089587, 0.0133435361793128, 
    0.0190807055121918, 0.0261585423690528, 0.0309744779245904, 
    0.0300146527819916, 0.0147690317513264, -0.000750620070941608, 
    -0.0180205636337403, -0.0291516853018662, -0.0146697275528704, 
    0.00628762866222783, 0.0237794782213751, 0.0274787526692709, 
    0.0236902765856256, 0.0260269817139355, 0.0577689560968447, 
    0.0791664332140285, 0.0571283497094981, 0.049714458075764, 
    0.0248764921950487, 0.00296529684059243, 0.000723558804441289, 
    -4.70616851080147e-05, -0.00232670544825368, -0.00267737762700323, 
    -0.00705480179856433, 6.21070332395735e-05, 0.0184322796176141, 
    0.0121260305304303, -0.0154161927433667, -0.0340408814156369, 
    -0.0348639043327941, -0.0276084492105327, -0.0213609522091978, 
    -0.0217701753894882, -0.0295589666745226, -0.0339645418601483, 
    -0.031990433053796, 0.00149743604418219, 0.0162687514430421, 
    0.0165006937225684, 0.0103520511983938, -8.03094057034703e-05, 
    -0.00251939409752146, -0.00644741818401939, -0.0158506414538326, 
    -0.0113158829537717, 0.029050877682954, 0.0353031607296941, 
    0.0315035401502085, 0.0212195949721265, 0.0169251015327925, 
    0.009738341974743, 0.0110260576579349, 0.0143778126647237, 
    0.0146789153319344, 0.0113336454916653, 0.0113675144997554, 
    -0.0165731921609747, -0.0287999042034279, -0.0208190278497629, 
    -0.001369446976522, 0.0252513575794833, 0.0344570603580397, 
    0.0290224071558848, 0.0281658778391802, 0.0628078609983508, 
    0.0931308654546957, 0.0905023012391209, 0.0649758848022841, 
    0.0460622895132567, 0.00394710545835058, 0.00138627290930944, 
    -0.00142929484967247, -0.00366857162778249, -0.00459002498101119, 
    -0.0118054406700408, -0.0123206097234233, 0.00335770476251509, 
    0.00907977792765262, -0.00695815412080423, -0.0228449291709474, 
    -0.0248660174610517, -0.0244890530764933, -0.02292710955924, 
    -0.024564849652579, -0.0357438829263867, -0.0364442215110115, 
    -0.0182779285938789, 0.009921832763495, 0.000850279358549977, 
    -0.0142088206157983, -0.0154834733243788, -0.0104869866761657, 
    -0.00271347760995614, 0.00300178111710324, -0.0022925566159203, 
    0.00975872651324024, 0.0401780185970868, 0.0544378373063183, 
    0.0425741652154204, 0.0201241214051508, -0.0033469263953904, 
    -0.0148167513995617, -0.0108722515394761, -0.00746729705972192, 
    0.000847389199513291, 0.0166896435940198, 0.0187137337747243, 
    -0.00989261886448128, -0.0364521122060302, -0.020158050916819, 
    0.00392318260530508, 0.0391174041048685, 0.0374573051578792, 
    0.0339293542053461, 0.0496924660554478, 0.0882412122435964, 
    0.0993015992473384, 0.101611753155608, 0.0745854480080178, 
    0.0549865853069268, 0.00722290427790179, 0.00421759373773351, 
    0.00333526585696116, 0.00158377538062621, -0.00324346750581035, 
    -0.00970041676509201, -0.0188773774993062, -0.00923274414625247, 
    0.000111446666546113, -0.00339904750375535, -0.0111848771160188, 
    -0.012502570834722, -0.0173770246415368, -0.0209080072933623, 
    -0.0221271939342213, -0.0311496405412286, -0.0297314516077604, 
    -0.0074075522293568, 0.0101978545835093, -0.00973437401708763, 
    -0.0305149369634949, -0.0276718073874432, -0.013755264309796, 
    -0.00157632587105576, 0.0106280183246589, 0.0118118272241629, 
    0.0248867600988776, 0.04599988418001, 0.0601503222661441, 
    0.045281968095564, 0.0233630669430528, -0.0119407890650169, 
    -0.0332575897403153, -0.0311520676551934, -0.0271733975713642, 
    -0.0100479888240294, 0.0165094075463229, 0.0219891783694236, 
    -0.00193051702598284, -0.0303474538031633, -0.022142365448897, 
    0.00578784638208503, 0.0356555130513533, 0.032986624592918, 
    0.0358520566965215, 0.058385869764981, 0.094835003619047, 
    0.110602504858718, 0.113155983620243, 0.0878822316631212, 
    0.0576580170707086, 0.00901258511014578, 0.00713442353771564, 
    0.00798841761313044, 0.00809342067765439, 0.0031176720951681, 
    -0.00143204783600236, -0.0154133735644303, -0.0139708923954794, 
    -0.0050930826347541, -0.00583122725595172, -0.00924067075706123, 
    -0.00842590608901404, -0.0123950796772744, -0.0161116864786163, 
    -0.0188949087941101, -0.0223785043613159, -0.0197084292516329, 
    -0.00186115106667, 0.0120192249418577, -0.00262814408934944, 
    -0.0183270184681208, -0.0212300826239562, -0.0156399027557393, 
    -0.00437295442063403, 0.0112322132912564, 0.0212292064653555, 
    0.03142652933665, 0.0476729585941816, 0.0535536310856736, 
    0.0592023661841266, 0.0171050023496239, -0.0211582882113549, 
    -0.0581388538367963, -0.0535324731712119, -0.0448812157362497, 
    -0.0264779227502042, -0.000210797782276273, 0.0207144677779532, 
    0.00471341504644234, -0.0195805238636902, -0.0137211060275018, 
    0.00411402591206054, 0.0240417307420105, 0.0207545142032041, 
    0.0242282156286434, 0.0486319660459029, 0.0735151812701682, 
    0.106214857059577, 0.108205974088448, 0.0880122454367313, 
    0.0539996638005609, 0.00855855269318943, 0.00670674394571659, 
    0.00862527913208692, 0.0103514171669755, 0.00967504619849252, 
    0.00752210493292437, -0.0049058664593592, -0.00764197175004767, 
    0.0024461915723482, -0.00305954524358108, -0.011363545331851, 
    -0.00971999248828735, -0.0099559071416046, -0.0109555221188932, 
    -0.0153834800209446, -0.0141269520106705, -0.0078127267056661, 
    0.00738469276927201, 0.0151804808459843, 0.0134032521983598, 
    0.0044800567851348, -0.00984884026330727, -0.0142903774154437, 
    -0.00309249559892259, 0.0137721150498689, 0.0211873567820239, 
    0.0280146126313695, 0.0372438128765268, 0.0450872037032029, 
    0.0469846896080498, -0.000806737600411939, -0.0479586427019185, 
    -0.0870214613938601, -0.0743195246265181, -0.0523922844574024, 
    -0.0386740212828352, -0.017742645609821, -0.0121117786749852, 
    -0.00156100450991561, -0.00968354815925352, -0.00191116538075868, 
    0.0124517927846486, 0.0202039195262102, 0.00852668265781462, 
    0.00122079424516501, 0.0127461247745295, 0.0384193458699123, 
    0.0758101527549309, 0.0823690982947969, 0.0689481199484988, 
    0.0456888506094185, 0.00324568522117163, 0.00168613606450722, 
    0.000650797708029329, -0.00258981085547046, 0.0010851088394249, 
    0.00603469502589858, 0.00811876493913796, 0.00833018892383202, 
    0.0143843157439903, -0.0122964746458981, -0.0274252873397242, 
    -0.0207578835214157, -0.0106037868373004, -0.00834433908088461, 
    -0.013092510690903, -0.00994829519183376, 0.000978644644515721, 
    0.00800857552070739, 0.0155150624663255, 0.0208163381636139, 
    0.0174195848857266, 0.000718570191715623, -0.00982905713216437, 
    0.00368518634776329, 0.0198841343648467, 0.0236234327996355, 
    0.0248948918963002, 0.0343963890094878, 0.0383139101710094, 
    0.0349398042003924, -0.00325882189749238, -0.0450230959161509, 
    -0.0756772568929402, -0.0666555778503114, -0.0506534446389463, 
    -0.0364096594085256, -0.0248183965552678, -0.0196192480495323, 
    -0.0135380634633447, -0.00630540100588323, 0.00649203861457668, 
    0.0180289546952504, -0.00624035039021809, -0.0101108933522518, 
    -0.00697551357186144, 0.00680221850707323, 0.0307061260002996, 
    0.0579019526731551, 0.0374471319766955, -0.00389204706462031, 
    -0.0049201340526142, -0.0128528212760949, -0.0252948590562124, 
    -0.0202578612375223, -0.00319267157190565, 0.0117255788090527, 
    0.0178847880264536, 0.0124499139502914, -0.0317935061949967, 
    -0.0472140485357127, -0.0338770930096479, -0.00940813477299099, 
    -0.00760866103568387, -0.0147978426256103, -0.0101876596501412, 
    0.00143199812403989, 0.00764930290334431, 0.0157711111388569, 
    0.0229514830075045, 0.0246178137976564, 0.0184079641811616, 
    0.00644262800232732, 0.0217717674702961, 0.0435434328848126, 
    0.042618564187683, 0.0373503305577608, 0.0378051287141803, 
    0.023655158936531, 0.0213383050692362, 0.00791800565024266, 
    -0.0248844409571308, -0.0357181985431526, -0.0439653967962481, 
    -0.0207005388673042, -0.0244629713423097, -0.0264728952137347, 
    -0.0257249775363761, -0.0149643505614729, -0.00810005060158427, 
    0.011415625063507, 0.018200437107743, 0.0131987435218938, 
    -0.00997836489907146, -0.0174924891925526, -0.00707949666943056, 
    -0.00529948838496466, 0.00854347020355303, 0.0109549749006364, 
    0.0100773676044689, 0.00870109902856375, -0.00984235721977989, 
    -0.0139469979108812, -0.0307583849427784, -0.0503539363254843, 
    -0.0398276196566671, -0.0135867963712318, 0.00464721800822211, 
    0.0142625069287142, 0.00312858123825323, -0.0335068047016003, 
    -0.0443429667597485, -0.0294813105442875, -0.00380239779507439, 
    -0.00368620991217761, -0.0142519699019373, -0.0112859080804787, 
    0.00109171051877533, 0.0106662170834016, 0.0169454040434187, 
    0.0183608670190453, 0.0251676740701056, 0.0391218117530561, 
    0.0447912015846162, 0.063211077241276, 0.0676435245846113, 
    0.0643748863473372, 0.0675875358091235, 0.0329548529781519, 
    0.0126688758631784, 0.0123984024827489, 0.0169945243524288, 
    0.0124462579396059, 0.0156093507865797, 0.00143143187213969, 
    0.00427149270385539, -0.0138034677159175, -0.0227290724099552, 
    -0.0253360598693861, -0.00906171697721608, 0.0044880088182207, 
    -0.00197137747374535, -0.0091959159023291, -0.0121245577376524, 
    -0.00654764145370976, -0.00453042953586825, -0.0151257461550762, 
    -0.01086196700453, -0.00390089005884144, -0.0110310712174129, 
    -0.0139265094567777, -0.0315862023195985, -0.0576866074677785, 
    -0.0522486795408954, -0.022072795481559, -0.00527008932291592, 
    0.000251717097737601, -0.0107620196226734, -0.032005106371696, 
    -0.0433755635641729, -0.0239838937525538, 0.0047240072536717, 
    -0.00520964801688316, -0.0222780683265067, -0.0197786171457797, 
    -0.00261181640923481, 0.0115224223063326, 0.0102399864690465, 
    0.00699917533974656, 0.0230861237761397, 0.0674778896842708, 
    0.0924538907548773, 0.112742823972242, 0.0915225770062972, 
    0.0731638706177969, 0.0524917776935987, 0.0197114840790081, 
    0.00367359566040241, 0.0228325565595263, 0.0289478023215203, 
    0.0224936804259704, 0.0179699067849205, 0.0136226984071948, 
    -0.00803542344397633, 0.00265278055001651, 0.00288509169329816, 
    -0.00611241936499688, -0.00776727853452111, -0.00757425036862025, 
    -0.0121919214693194, -0.02711970187834, -0.0132398971519017, 
    -0.00402625559493886, -0.00672349684261944, -0.0055745558174591, 
    -0.0178568958293057, -0.0424208578630364, -0.0446790040397828, 
    -0.0193815294232531, -0.00643743341035793, -0.00585025538893316, 
    -0.0151008730987586, -0.0300867422422827, -0.0389527353867808, 
    -0.0154311443964605, 0.0119789622758653, -0.00551369615141385, 
    -0.0333824849058537, -0.0361175407587929, -0.0157635548065259, 
    -0.00522884093877277, -0.0139771999005611, -0.015473888111732, 
    0.0224655114855327, 0.100106513781064, 0.140351996574854, 
    0.1431750620152, 0.0947489717912541, 0.0753670389005912, 
    0.0511831726661592, 0.0216404750547465, -0.00654489169788272, 
    -0.00779375710078482, -0.00698073165509227, -0.026811026901715, 
    -0.00283612027101297, -0.00126741227526062, -0.00882944454037951, 
    -0.0224636407370705, -0.0285455468384978, -0.0160265086618378, 
    -0.00593529970765077, -0.00985499941421424, -0.0199485418343057, 
    -0.0296635157358533, -0.0267978386038141, -0.00911286742491078, 
    0.0189600263342119, 0.0126305102516011, -0.0259562711123956, 
    -0.0437263859930805, -0.0297077195150066, -0.0310344433874658, 
    -0.0533368078193225, -0.0399581783695847, 0.0285409162768668, 
    0.122451541514318, 0.145004572520701, 0.132896546645157, 
    0.0731049545069171, -0.00151580431280475, -0.00184900983460665, 
    -0.00532455168119875, -0.00855860952566953, -0.010641891070289, 
    -0.0052613461366105, -0.00788775710277442, -0.0180182709461846, 
    -0.0294012925184101, -0.0384482836712446, -0.0291518799586765, 
    -0.0140853217742921, 0.00814967008771999, 0.017854063424587, 
    -0.00774360625398549, -0.043426296385424, -0.0521760458963638, 
    -0.0501181687306996, -0.079859069294785, -0.0735024375927214, 
    0.00646279896709412, 0.124590874148857, 0.147823352866937, 
    0.126436290327959, -4.1374527638143e-05, -0.00313207909139559, 
    -0.00507643592325533, -0.00443713376358691, -0.0027261325698113, 
    -7.22427799961706e-05, -0.00417757452321218, -0.0100121338780843, 
    -0.0157258470277169, -0.0343815490427062, -0.0405163136964057, 
    -0.0281923909846342, -0.00283232065104689, 0.00988522042624632, 
    -0.00970343811198974, -0.0356765992254925, -0.0569393421781021, 
    -0.087620676873971, -0.085709965448368, -0.0513463673166596, 
    0.0276119410225075, 0.0841477121617177, 0.00196686005895379, 
    -0.00614169188396948, -0.00813864132854042, -0.0037741416510496, 
    0.00133857893406591, 0.0060484806121137, 0.00564100309031284, 
    0.00496487344952359, -0.00191750550355653, -0.0217924150306363, 
    -0.0294571497125062, -0.0225028975285868, 0.00101600636586129, 
    0.0104586298377216, 0.000712277796798405, -0.0217407783810915, 
    -0.0535092831284942, -0.0816026370389952, -0.0712628485603124, 
    -0.0230489376002763, 0.0408865169398146, 0.0737902025551134, 
    -0.000524765766437771, -0.0122086753127873, -0.0142483340738841, 
    -0.00772092871141403, 0.00161641604791481, 0.0101668826336512, 
    0.0135217750658157, 0.0104480516886597, -0.00492063038050844, 
    -0.0148659547860543, -0.00944246496355359, -0.00510760691230395, 
    0.012781020134998, 0.0251678713473691, 0.0236969561979199, 
    0.00382490136972111, -0.0293065275920988, -0.0726250668373122, 
    -0.0733826835978016, -0.0577043469168009, -0.00793113500085236, 
    -0.0165755946841135, -0.0118367951586865, 0.0037341983270906, 
    0.00628709642967677, 0.0126734605116133, 0.0113244672723101, 
    -0.00505698795482501, -0.0182876194209186, -0.0220841562169151, 
    -0.0081698636285583, 0.00264779560962879, 0.0229411632469492, 
    0.0415725743913535, 0.0411972723333602, 0.0279481826786138, 
    -0.0131159733432911, -0.0484378004049246, -0.0702961343241744, 
    -0.00895808333866516, -0.00523069711431023, 0.0133140910445611, 
    0.038816664504107, 0.0236486588590704, 0.0179670003483401, 
    0.00191880162494297, -0.0253805754015777, -0.035238706429571, 
    -0.0409585526380898, -0.0286728550560301, -0.00783797385827718, 
    0.0101203961578317, 0.0348290956582818, 0.0437240287867484, 
    0.0369971278104227, 0.0170998017052101, -0.00531409692719813, 
    0.00852006686532344, 0.0322321133387217, 0.0510755097870108, 
    0.0469782599063721, 0.0311255005493034, -0.00673369289874253, 
    -0.0404165249481499, -0.0552708755240506, -0.066920646674351, 
    -0.0641730414812002, -0.0443100695557266, -0.0313028607573568, 
    -0.0155438263128351, 0.00696216306138257, 0.0351816247400442, 
    -0.00725578203739818, 0.00588382315921131, 0.0242899597500075, 
    0.034384448134386, 0.0451563399799534, 0.0339472960777689, 
    -0.0164253958174576, -0.0585813191343392, -0.0717770155953744, 
    -0.0911407635734816, -0.0895948427247212, -0.0770356145140772, 
    -0.0821856210811707, -0.0678569685360819, -0.0171806569231358, 
    -0.00941085607648738, -0.0042425765435943, 0.00166376222752734, 
    0.0065049425993526, 0.0149480426592947, 0.0134052748706434, 
    -0.0328984435015033, -0.0527971318981953, -0.0664931396259918, 
    -0.102026883689559, -0.10152942002116, -0.0937039078850271, 
    -0.0925481118821919, -0.0859465620665076, -0.0153934522875511, 
    -0.0188724327858383, -0.0255548911563259, -0.0210381639648036, 
    -0.0138639859353798, -0.0127616080134774, -0.030617988321667, 
    -0.0257265573798571, -0.0459523343740555, -0.0867118199796698, 
    -0.0908642335593132, -0.0698827501210436, -0.0215520276747471, 
    -0.0265375487373593, -0.0384141331699972, -0.0342154562828392, 
    -0.0274724707736705, -0.0216701470859825, -0.020189595720032, 
    -0.0118183755959292, -0.0382843935130609, -0.079357936198331, 
    -0.0842247266131019, -0.0611438555396144, -0.0307245973170921, 
    -0.0351051395333744, -0.0460427194596119, -0.0453993492659526, 
    -0.0416239116355991, -0.0415701722012592, -0.0313402287525077, 
    -0.0236248842583811, -0.0473294462641887, -0.0805725675479424, 
    -0.0815204471491519, -0.0508759886750857, -0.0351233291504198, 
    -0.0398842228397678, -0.0502653257847133, -0.0499456291846109, 
    -0.0282387142218557, -0.0331075240887595, -0.0328699260022792, 
    -0.024930243020255, -0.0430073550484853, -0.0759893923819473, 
    -0.0817599694469444, -0.0321404621126467, -0.0469292178596535, 
    -0.0552093489067155, -0.0384317296343241, -0.000969886743121945, 
    0.010530935414228, -0.00210473626033571, -0.00840696363868607, 
    -0.0294785344186545, -0.0671351697290764, -0.0714840603936897, 
    -0.028233345375127, -0.0444865624676434, -0.044901345179987, 
    -0.0101982934821306, 0.0314593228135904, 0.0429961041406322, 
    0.0170960539263598, -0.00750480431893709, -0.0189768412660489, 
    -0.0439460720315647, -0.0527625704654941, -0.0239564116105772, 
    -0.0409068478493075, -0.0309476994653602, 0.00716603018119585, 
    0.0282831593837237, 0.0283054924933171, 0.00539925825922784, 
    -0.00961635674705976, -0.00587081858277216, -0.0088077376924871, 
    -0.0122713513110694, -0.0296854157503556, -0.0239033794505264, 
    0.00400086991417553, 0.0130532955931777, 0.00714299649442039, 
    -0.00656741179944016, -0.0104227131983774, -0.00472296929931649, 
    -0.00412838486168937, -0.0183677099830041, -0.0176898674671224, 
    -0.000397820970418622, 0.00561226414951842, 0.00257973866980847, 
    -0.00686932271839843, -0.00477443766442028, -0.0038832638117445, 
    -0.00343138727383189, -0.0150308440286868, -0.0148731301217866, 
    -0.00476790327153682, 0.00217039514734206, 0.00260046989682835, 
    -0.00150713356154028, -0.00140484186853836, -0.00624344690469078, 
    -0.0187784208235269, -0.0172311336977931, -0.00921997744068727, 
    0.000234727545149809, -0.01012008708788, -0.0160559471621392, 
    -0.0138438841402205, -0.00944193620416069, 0.00939874858741466, 
    0.00938544242335415, 0.00973174653462426, 0.0153988500471782, 
    0.0260765438008861, 0.0330674977010336, 0.0394598331358816, 
    0.0357696555218787, 0.0222178332937801, 0.012615272021835, 
    0.00291393973847537, -0.00229521451818253, -0.00247965346862399, 
    -0.00124966834621031, -0.0026977406545054, -0.00268445334538435, 
    -0.00212486507745284, -0.00201618433835483, -0.000860174993006748, 
    5.85330027129508e-05, 0.00054740824325609, 0.000504003200546854, 
    -6.10632275503112e-05, -0.00375129655308521, -0.00366083821178191, 
    -0.00231953045398949, 0.00226334853667964, 0.0063560145862741, 
    0.00618523666003412, -0.000394093511172144, -0.00673266900322799, 
    -0.00695345874663732, -0.00466790052980686, -0.00123293422705612, 
    0.000678363417706826, 0.000829783978380876, 0.00126332810930015, 
    0.00161197514592203, 0.000571438729049213, 0.000145398862564207, 
    9.22012908221222e-05, 8.14323118930599e-05, -0.000182385132235097, 
    -0.000387443611594562, -0.00038841343166561, -0.000170751098005313, 
    -0.00712151947050094, -0.00668047852269124, -0.00490949382111152, 
    -0.0011962510340937, 0.000857995917709038, 0.000392981259184617, 
    0.00267205251559942, -0.000598604327337183, 0.00333393796316395, 
    0.00551679102761013, 0.000914806252745588, -0.00102358629859664, 
    0.000179808662969059, 0.000363113127145606, 0.00039475991932671, 
    0.000222495545422506, 2.90283038841732e-05, 7.06854013601823e-05, 
    0.00012473677729299, 6.38875173775998e-05, 2.61066012095779e-05, 
    3.08673822021094e-06, -1.93367127416973e-05, -0.0013650417717806, 
    -0.00124916767872812, -0.000706300483624707, 0.000644336283216715, 
    0.00183442613629016, 0.00233194845372159, 0.000951536869157445, 
    -0.000288249636626607, -0.000714447479535732, -0.00109666195234618, 
    -0.0004174585022754, -0.000203550832825688, -0.000161683189719927, 
    -0.000212118461190355, -0.000203739258067454, -3.89573467861957e-05, 
    4.73526818841873e-05, 2.57349103130409e-05, -1.31004866853991e-06, 
    -8.11140404510059e-06, -1.16794963960197e-05, -1.82315333433943e-05, 
    -1.63600890662674e-05, -0.00345050184644121, -0.0077821187067063, 
    -0.000416581749801136, -0.0136665292824357, -0.0138301496933767, 
    -0.0148379258826094, -0.0202851601434395, -0.0212065788656745, 
    -0.0159222283499325, 0.000979394451906968, 0.0075455971970464, 
    -0.00650809412779267, -0.00163047815175185, 0.000145787898927099, 
    0.0018583629838416, 0.00238718389215246, 0.012334109652096, 
    0.0164050576541998, 0.0146251243193777, 0.00807594252226356, 
    0.00309382391236832, -0.00163674028747339, -0.0069575860533185, 
    -0.0137259765231129, -0.0138649499580657, -0.00770911243418054, 
    0.00501089273738206, 0.00912377120806369, 0.0134798099646605, 
    0.00936057107853355, 0.00292271869327141, 0.000561165052438765, 
    -0.00596635680699085, -0.0146241196528327, -0.0275993409374118, 
    -0.0334249432463335, -0.0473560656829578, -0.0202600476287102, 
    -0.0184134643174014, -0.0116845036315779, -0.000696632135777607, 
    0.00602990985231446, 0.0122125531565268, 0.0310724159112397, 
    0.0396986047782759, 0.0358338132531728, 0.0285713424323505, 
    0.0269650916013883, 0.0243115154775857, 0.016378001998227, 
    0.0127461038010652, -0.00211635169043248, -0.033894297452557, 
    -0.060438423166982, -0.0680778712131342, -0.038301675628211, 
    -0.0177416256859712, -0.00986788920929595, 0.00796446168719113, 
    0.0223787730352732, 0.0236180599658587, 0.025287195211993, 
    0.0196232941075925, 0.0118761009723588, -0.0196300983728431, 
    -0.0376605664685419, -0.0689652460418013, 0.0111402408440278, 
    0.0146541135653461, 0.0149422637359028, 0.00740977823775836, 
    0.001284080504806, -0.0025950615158852, -0.0112852201667282, 
    -0.019094400224621, -0.017632852664506, -0.01024271891034, 
    0.00941081062401785, 0.0157234183298296, 0.0128146110834956, 
    0.0082989409235702, 0.0036144849107774, 0.00394776141854348, 
    -0.0023733156188502, -0.00502634566650348, -0.0110646307582193, 
    -0.0358358670886967, -0.0505706538041059, -0.0112378348134175, 
    -0.00309386787801001, -0.00510676565271754, -0.0012626191931171, 
    0.00125018235489418, 0.00590099599543875, 0.0310610120159441, 
    0.0415974683047031, 0.0332117970260216, 0.0282682705509161, 
    0.0251052677568531, 0.0167196476873858, 0.00541011028052978, 
    0.00997424302038228, 0.00557521416330813, -0.0227423866479986, 
    -0.056266436460136, -0.0733868552813857, -0.0608733350706587, 
    -0.0436853663028577, -0.0249982282899371, 0.00492587277943951, 
    0.0239224354895916, 0.0274872333591337, 0.0227265382734313, 
    0.0126259027069125, -0.000799630252083944, -0.0386186661193793, 
    -0.0561486306375177, -0.0703516543030713, 0.00584659048451277, 
    0.00847069576081169, 0.00664216314028962, 0.00223391471794964, 
    0.00286617536365497, -0.00221696683166707, -0.0144133674296155, 
    -0.0219388967317684, -0.0200445059038878, -0.0132252530517721, 
    0.00314569748768313, 0.00729042119013558, 0.0112790535563593, 
    0.00509106559434032, 0.00520560822697874, 0.00886610642080973, 
    0.00739924226305445, 0.00719292187991404, 0.0100552471671449, 
    -0.0402348914056974, -0.0416935540515174, 0.00275073041461074, 
    0.00773477051727923, -0.000393862224328268, -0.00557882701786812, 
    -0.0047380924955317, 0.00706877210691417, 0.0327781815281473, 
    0.0372747298852126, 0.0270342643286349, 0.0187797281446856, 
    0.0144346649422551, 0.00328708491388056, -0.00298139863662582, 
    0.00333655684867928, 0.0050368601221094, -0.0150143806519736, 
    -0.046480664778716, -0.070624125456991, -0.0627781779499903, 
    -0.0456037249270805, -0.0247615799498561, 0.00983689826541969, 
    0.0291097662565605, 0.0362613198888728, 0.0166730020163564, 
    0.00813207560424613, -0.00131372965647393, -0.0477510527640101, 
    -0.0752634269476704, -0.0824198560545533, 0.00416371311219802, 
    0.00184950876513355, 0.000218756375370311, 0.00257238603432961, 
    0.0135524971800437, 0.0109365605267675, -0.00311451829049571, 
    -0.012690089451704, -0.0165923759502282, -0.018791733012041, 
    -0.0104897634024544, -0.00289926250159522, 0.00691462890441032, 
    0.00135414997491056, 0.00414031253682649, 0.00963318350421554, 
    0.00948819342216477, 0.0135995162342039, 0.0261265241327451, 
    0.00145795394426433, 0.0144583484467756, 0.0260157082404638, 
    0.0115912268351961, -0.00404222237876997, -0.0106468963558756, 
    -0.00870158483094087, 0.00313669949848873, 0.0206903360980501, 
    0.0182405060850313, 0.00690974729274762, 0.0138116036786341, 
    0.00768483115617258, -0.00147901916241296, -0.00725906655743717, 
    -0.000868752914050001, 0.0031441187905829, -0.0131318341432999, 
    -0.0371593021727649, -0.0605568414657853, -0.0534913486945782, 
    -0.0231249162838162, -0.0148853808985572, 0.0211606342289531, 
    0.0568641838508499, 0.0605212565130717, 0.0375557485170599, 
    0.0249064482143214, 0.0106811595595861, -0.0305708043446497, 
    -0.0689792179959022, -0.0670169517316159, 0.0076462091545449, 
    0.00315437691192962, 0.00128219817984721, 0.00927303821237106, 
    0.0291346552026881, 0.0356751264214176, 0.0161008177205214, 
    0.00046155655007885, -0.0144092875905888, -0.026933873473503, 
    -0.0276594139631954, -0.0174233412177534, -0.000670535298919567, 
    -0.00364525728730633, -0.000790255840146602, 0.0032932641630234, 
    0.0027258174939165, 0.0151365480508799, 0.035610928731062, 
    0.0232854736835259, 0.0190247478852131, 0.0158270472464319, 
    0.00537910861296864, -0.0102386574356191, -0.0141814106911023, 
    -0.0117868766868717, -0.00404020858986763, -0.00307192943078893, 
    -0.024390799203353, -0.0262676693795395, 0.00213739833851067, 
    0.0020462170753873, -0.00207652769827268, 0.0015511223187134, 
    0.0150599556478641, 0.0298593287894323, 0.0205417641857933, 
    0.0123327989924781, -0.0427505806641702, -0.0357767661686599, 
    0.00148199615623103, 0.0169615025609933, 0.042531736457, 
    0.085843153242122, 0.0817839148871866, 0.0642629043116274, 
    0.0387939710903704, 0.00837212952554389, -0.0359224544538554, 
    -0.0686783605702204, -0.0583201659605734, 0.0126276794170485, 
    0.012045944744606, 0.0109363960553206, 0.0169417724663278, 
    0.0296290831904517, 0.0481170451372188, 0.0369111140796701, 
    0.0106243672981888, -0.0110750792601529, -0.0342528391542028, 
    -0.0408869948870174, -0.0251607602815097, -0.00926216322145084, 
    -0.0106517152590082, -0.00999046056803017, -0.00945155930522555, 
    -0.0111042556402501, 0.00716880261076216, 0.0143337814293332, 
    0.00632695502739724, 0.0103999115755675, 0.0157056320346183, 
    0.00433399608597575, -0.0134614035674798, -0.0121224706334607, 
    -0.0110583511212164, -0.0116856509132323, -0.0301074824718448, 
    -0.0605091354564181, -0.0494661372089817, -0.00571689501836449, 
    0.0045183553664292, 0.00586613667623056, 0.0164805914621003, 
    0.0355187997870224, 0.0495454877297174, 0.0472701483280652, 
    0.0283996434189786, -0.0171140246098715, -0.0197259571473385, 
    0.0155748048678624, 0.0432266680781974, 0.0607150769667978, 
    0.0909266474258928, 0.0802777668692184, 0.0665132696523336, 
    0.0483389332546979, 0.016303532068711, -0.0158569775287696, 
    -0.0440664803223394, -0.0450751005033664, 0.0145880195903019, 
    0.0188104783978511, 0.0182066186070226, 0.0188083679147405, 
    0.0236371546897215, 0.0400702889883097, 0.0413141019220872, 
    0.019581820571641, -0.00481910170336543, -0.03654634798661, 
    -0.0467374618233172, -0.0306701806261398, -0.0161179397114542, 
    -0.0165415529747153, -0.0184467978950446, -0.0246824548906602, 
    -0.0243998152924819, -0.00406560639141231, -0.00611763112195431, 
    0.00749790631944238, 0.0178077286329995, 0.0243530730266088, 
    0.0123881836942552, -0.00797234353103071, -0.00936430076537046, 
    -0.0153373175139191, -0.0264636151631701, -0.0472837884157539, 
    -0.0455762014918103, -0.0629548918086589, -0.0131417164470411, 
    0.00944443120480266, 0.0152385804469677, 0.0280084781296638, 
    0.0473204323381695, 0.0466036268667937, 0.0317960781630926, 
    0.0233553284878009, -0.00312586136702472, -0.0146182385876421, 
    0.00685255709948926, 0.0409487913284329, 0.0695277555684837, 
    0.0725899058971273, 0.0618622564540393, 0.0632491047006376, 
    0.0747741298413111, 0.0407088101432353, 0.0142678996989786, 
    -0.00662088630496221, -0.0213051939583181, 0.0128826460131416, 
    0.0144974478916745, 0.0179225805301479, 0.0083442720813137, 
    0.0142080648763972, 0.0256072202646306, 0.0397186181673853, 
    0.0273025958513546, 0.00157474986153798, -0.0323886068178666, 
    -0.043499505837265, -0.0342185643277199, -0.0231815075124204, 
    -0.0209632828240616, -0.0217074283517288, -0.0281133297098934, 
    -0.0313400842902912, -0.0154831519565146, -0.011250403236554, 
    0.0131207644245579, 0.028521809970853, 0.0316937538917541, 
    0.0176360322064866, -0.00138993327357574, -0.0102131662176345, 
    -0.0230461294252227, -0.0291444993586911, -0.0117287512130403, 
    -0.0176332278923306, -0.0171488732262284, -0.00942452329065003, 
    0.00591322881616464, 0.0175866376588183, 0.0332448079148446, 
    0.041106755598637, 0.0323317342987007, 0.0109135485586756, 
    0.000964096739093842, -0.00625014593604514, -0.016235785914822, 
    -0.00691022193236074, 0.0175098725403017, 0.0400428369750654, 
    0.0444549153341857, 0.0380441434254035, 0.0366057127791431, 
    0.0624547980163146, 0.0632599797208455, 0.0427143426837508, 
    0.03579509948369, 0.0103363368586803, 0.00453421288741817, 
    0.00722454154369185, 0.00686290063331998, 0.00295859521116906, 
    0.0019241395635907, 0.00539206547868816, 0.0147373688471621, 
    0.0252667960784277, 0.00889058043380437, -0.02840095752765, 
    -0.0388519909536644, -0.0339994475239602, -0.0250182750520923, 
    -0.0226372497288417, -0.0226064496404153, -0.0254537489342881, 
    -0.0314294405875878, -0.0281305917414624, -0.00777535510815817, 
    0.0152547230928868, 0.0292704778335624, 0.0284283761781806, 
    0.0120420928432093, -8.83188979925049e-05, -0.011948806836698, 
    -0.0253472308577713, -0.0219883776724751, 0.0228698328136405, 
    0.0164490550796165, 0.0192019196860823, 0.0124581157038936, 
    0.0100819186902411, 0.0169597773176338, 0.0280503481250155, 
    0.031653698477675, 0.0299352045355173, 0.0122288609164239, 
    -0.000456719915876219, -0.0164733829603632, -0.0277469007462479, 
    -0.0149385822821357, 0.00730605445631651, 0.0238723055916035, 
    0.0296343461187023, 0.0257504868623303, 0.0232014340966982, 
    0.0512436994566199, 0.073272679705913, 0.0503612258436497, 
    0.0530970284759963, 0.0201497347743174, 0.0026035243517032, 
    -5.46001401684932e-05, -0.000326556241759197, -0.00253251200452039, 
    -0.00253055848142491, -0.00684266429741075, 6.40024080919431e-05, 
    0.0182265438760031, 0.00887439805127215, -0.0240967748582722, 
    -0.037143941248514, -0.0311584086607699, -0.0222955137994039, 
    -0.0186751254578064, -0.0206443771812782, -0.0287014767102682, 
    -0.033837437085844, -0.0360140415335848, 0.00109374525931584, 
    0.00599008998357883, 0.00878142284386831, 0.00849827965966255, 
    0.000545736654815517, -0.00325301218325524, -0.0134021293331676, 
    -0.0247944570948041, -0.0197279933922091, 0.0294130487780227, 
    0.0450094883822578, 0.0379604809044244, 0.0204746680129091, 
    0.0158025908798385, 0.0113317448211624, 0.017236275051512, 
    0.0185002271111295, 0.0187777850378442, 0.0120916069816616, 
    0.0149391165832436, -0.016571850006328, -0.0269858986364192, 
    -0.0194514774030765, -0.00341904456842854, 0.0203046353610831, 
    0.0344535761102532, 0.0309093280742746, 0.0264864083983354, 
    0.0543810465624877, 0.0865260347252552, 0.0855742161821912, 
    0.0687229755402967, 0.0449124981265959, 0.00386816674580851, 
    0.00144698214862707, -0.00171729038683024, -0.00387131240580374, 
    -0.00458513728662095, -0.0110741862474326, -0.0115865539488241, 
    0.00360201861732534, 0.00806348961900681, -0.0135162646675836, 
    -0.0279361468202983, -0.0248304914064819, -0.0228200235058042, 
    -0.0230635430198612, -0.0241980559662076, -0.0336333751697952, 
    -0.0338463201416348, -0.0178395652640375, 0.00882919166623188, 
    -0.0107750880854896, -0.0201063050242543, -0.0133365316356501, 
    -0.00822436653805257, -0.00308601738069507, -0.00488682460800825, 
    -0.0182297963743737, -0.00656330928848406, 0.0364829006870078, 
    0.0573194705928078, 0.0412111873602238, 0.0161070177373172, 
    -0.0083732841925286, -0.0130695786570124, -0.00307934807344482, 
    -0.00237788094740281, 0.00346991392979221, 0.0180392280125839, 
    0.0176222414393227, -0.0137570917202799, -0.0356306196186051, 
    -0.0179857578291544, 0.00858163015150877, 0.0411740606633541, 
    0.0365516419144333, 0.0340965895140095, 0.0488608764573181, 
    0.0840611886708711, 0.0973785643124282, 0.102752785864926, 
    0.0756650614479656, 0.05546017760219, 0.00699306128335316, 
    0.00373755407939866, 0.00358283545481008, 0.00267247577985242, 
    -0.00361557569610229, -0.00999124435571196, -0.0186988811321971, 
    -0.00759624279399842, 0.00184657866801939, -0.00491296622741065, 
    -0.0144082538653243, -0.0138991497940248, -0.0160382534479779, 
    -0.0202334327617867, -0.0227025364814964, -0.0325035362825145, 
    -0.0329001712513032, -0.0100035858874344, 0.00672626453635588, 
    -0.0191910068487716, -0.0330556009352071, -0.0222088173292285, 
    -0.0089468377334547, 0.000744252151069349, 0.00616942877992229, 
    -0.00561723530713553, 0.0100804615341321, 0.0409881447782826, 
    0.0593132391418359, 0.0478042804517596, 0.021422996241051, 
    -0.0153163071645419, -0.0327993163199823, -0.0267777594356043, 
    -0.0243969085926121, -0.0118053163168549, 0.0116839954462292, 
    0.0209683784165664, -0.00631024711586117, -0.0316038084955046, 
    -0.0191314751741569, 0.0107939001202807, 0.0357904446887144, 
    0.0321701443919123, 0.0386388664343593, 0.0627163514306933, 
    0.0971582328094002, 0.10774273141287, 0.113012999135202, 
    0.0894130832553424, 0.054042348222641, 0.00845073036685038, 
    0.00700960355351067, 0.00845642263149425, 0.0091723888056703, 
    0.00209566367482219, -0.00341674999761608, -0.0179365465795228, 
    -0.0131332478656849, -0.00447799535756953, -0.00589887859580396, 
    -0.00976105572682882, -0.00889095422379317, -0.0111028371665229, 
    -0.0140860284126648, -0.018008453278241, -0.0256477162312127, 
    -0.0270625017141993, -0.00862534538280188, 0.00996374458242292, 
    -0.00718882561609814, -0.0175720354172514, -0.0173127313887036, 
    -0.012694756502278, -0.0017890232345586, 0.0110295423466785, 
    0.0115429637730947, 0.0263112886980799, 0.0462936776485848, 
    0.0524565277614689, 0.0579365855865485, 0.0109430338199124, 
    -0.0182781740903455, -0.0587793991337848, -0.05132264274368, 
    -0.048242984754464, -0.032795837123627, -0.00982565484825998, 
    0.0173610400088633, 0.00350351142514889, -0.0198983981629532, 
    -0.0116161089047517, 0.00720581239330484, 0.0231587924391879, 
    0.0188488158531198, 0.0257935070942199, 0.0546787250336963, 
    0.0737157156515331, 0.10693086890883, 0.108455785500949, 
    0.0870347530579739, 0.0511849437063898, 0.00728543982537772, 
    0.00597940755876277, 0.00844455938535936, 0.00922479833249716, 
    0.008597035451759, 0.00584941902609572, -0.0111157059860317, 
    -0.011812282801145, -0.00130480075782286, -0.00337775805732022, 
    -0.0108181874093184, -0.0101378714187394, -0.00997925625597843, 
    -0.010094480790527, -0.0150378427552684, -0.0168761435938176, 
    -0.0157492972847202, 0.00181444390159487, 0.0147443047280663, 
    0.0143437246133958, 0.00720714630976093, -0.00721182744312572, 
    -0.0114754038456132, 0.0005377327736886, 0.0150461813957905, 
    0.0207329438612899, 0.0304591903692364, 0.0380750495468533, 
    0.0457500909360469, 0.0463394020605235, -0.00308737582550166, 
    -0.0443086660028351, -0.0851729535354595, -0.0741964032572985, 
    -0.0547087485505656, -0.0408808816600169, -0.025627777809835, 
    0.000461090296281638, -0.00862002788276406, -0.00444955282748367, 
    0.0112892988496758, 0.0201634286300532, 0.00831593608315519, 
    0.000403323691839105, 0.0112380928817423, 0.0374797971663154, 
    0.0762954621070507, 0.0795648662845796, 0.0641948837143891, 
    0.0449458856742374, 0.00155874307180865, -0.000154959222096639, 
    -0.00331707360662, -0.00837082258346115, -0.000416996933463017, 
    0.00567427576414486, 0.00299936729695442, -0.000804936255963914, 
    0.0121993272383779, -0.0103403485549356, -0.0251284224027966, 
    -0.0219629514346108, -0.0102151668609101, -0.00817910111047566, 
    -0.0127721752537151, -0.0104365388410302, -0.00143638869551779, 
    0.00747507781360345, 0.0159085245030846, 0.0222111315819924, 
    0.0212644615598021, 0.00326224548178784, -0.00968653349571057, 
    0.00593731911491949, 0.0194955509084443, 0.0223289056790947, 
    0.0229310730648557, 0.0340879922429451, 0.0393403167084415, 
    0.0339440487336921, -0.00441355573444749, -0.0442878203981453, 
    -0.0712389803733993, -0.064476271121632, -0.0483790799370624, 
    -0.0334949595550116, -0.0258436235511613, -0.0179808713008376, 
    -0.0108742566777258, -0.00863253409832324, -0.0013840179359831, 
    0.0169004782975923, -0.00292230139374728, -0.0126528350173417, 
    -0.00808802956547723, 0.00206262673968533, 0.0279422738625419, 
    0.0568005052456633, 0.0353602833293981, -0.00581938159210118, 
    -0.00881030734861891, -0.0211663115252162, -0.0327827542509795, 
    -0.0224721316350837, -0.00320900468742467, 0.00993667246922884, 
    0.0117053976626997, 0.016930988575474, -0.0232056853949006, 
    -0.0451802270776502, -0.0352415466505701, -0.00764516167437329, 
    -0.00774618891030274, -0.0145013475238949, -0.00786738812211912, 
    0.0032453687605572, 0.00960476043314446, 0.0173193157804615, 
    0.0242078967320134, 0.0266670742570978, 0.022958630102796, 
    0.00584708962513591, 0.0244551823925018, 0.0417935364836423, 
    0.0338862973777075, 0.030042391086575, 0.0390322655278863, 
    0.0238667555117004, 0.0217125966294981, 0.00831202654600124, 
    -0.0282416504129751, -0.0336140584006227, -0.0503743160439596, 
    -0.0228066042152366, -0.0204459674590798, -0.0258681758701464, 
    -0.023906845106119, -0.0140333515686766, -0.00814358914012495, 
    0.00830995925993101, 0.0173363989006531, 0.0138403111835047, 
    -0.0124117410210956, -0.01745988077752, -0.00794538944319229, 
    -0.00739106316947924, 0.00724887310752534, 0.0125633654711901, 
    0.0096298290496014, 0.00960689858757181, -0.0116106115224982, 
    -0.0188788833018826, -0.0387100697274504, -0.0539873129323738, 
    -0.0390116759294634, -0.013275782375441, 0.0037827702482459, 
    0.0146446458096933, 0.0147934241911398, -0.0203546692198335, 
    -0.0424702207464672, -0.0316858397424973, -0.00286231420350638, 
    -0.00671468614272245, -0.0145930018037061, -0.00736423057829895, 
    0.0037918059979308, 0.0114818792516781, 0.0179797498728842, 
    0.0184692259555076, 0.0251116978557391, 0.0433621484067718, 
    0.0437461955438061, 0.0669593170905113, 0.0639819190859364, 
    0.0542626281909975, 0.0646931363471602, 0.039202223836426, 
    0.0185083571947354, 0.0118259687376311, 0.0146141084476649, 
    0.008513973385369, 0.0207159644340146, -0.00276247249819027, 
    -0.000651576759601075, -0.0229682004807556, -0.0237843125794133, 
    -0.0114223933458574, 0.00624062981748244, -0.000642474540572308, 
    -0.00744644312800812, -0.0113350795022117, -0.007313353958453, 
    -0.00359072892531735, -0.0137465085351731, -0.0119021411876124, 
    -0.00666914112102903, -0.00994483177681676, -0.011757289631226, 
    -0.0285422052657857, -0.0537008212584313, -0.0480167129592673, 
    -0.0215836690052727, -0.00606829892865549, 0.00449769577006032, 
    -0.00120314961916763, -0.0245007909979012, -0.0408131400162044, 
    -0.0231639271967852, 0.00320353482169132, -0.0139942663210969, 
    -0.0262015561435998, -0.0157964073009108, -0.00186667613641844, 
    0.0110563670937955, 0.0101837870468551, 0.00514968240219729, 
    0.0192897284073661, 0.0714187111220215, 0.0916007532925164, 
    0.116444196408612, 0.0893830152390311, 0.0684075731169816, 
    0.0617536195206987, 0.0278962958862707, 0.00666990447839573, 
    0.0211033940294663, 0.0266887207153524, 0.026536294170931, 
    0.0164182449673599, 0.00164663481315417, 0.00603341487826909, 
    -0.0032682313441029, -0.0073357365747703, -0.008156799091027, 
    -0.0111053290582874, -0.0267795975901705, -0.0154296269473529, 
    -0.00448930487715649, -0.00524641931486664, -0.00250164916241119, 
    -0.0094202131636004, -0.033027358709946, -0.041531284041193, 
    -0.0198449433876228, -0.00618100135723596, -0.00397843345966772, 
    -0.0126736865244469, -0.0295869009787129, -0.0396762287340061, 
    -0.0137845021911689, 0.00964367570020448, -0.00914199150245678, 
    -0.0349149650939953, -0.0357246952210443, -0.0190864736910554, 
    -0.00704327915018401, -0.0157127377643733, -0.0185765927150633, 
    0.0166171332987807, 0.0944647358690676, 0.139425184142885, 
    0.138610544578553, 0.0922333609626918, 0.0774286252510146, 
    0.0586169332540385, 0.0268907186095098, -0.00534786618812276, 
    -0.00710609028900483, -0.00704907224900966, -0.0258721312536261, 
    -0.00257022338507085, -0.000815473543119745, -0.00448162652635405, 
    -0.0160735318683972, -0.0255804001260676, -0.0173890267477736, 
    -0.00644119518690238, -0.0130650874464634, -0.0233805133449683, 
    -0.0315925308796778, -0.0292401072174847, -0.00864716405126567, 
    0.019098924055886, 0.0158571487382524, -0.0181118942248182, 
    -0.0425309977912115, -0.0307706703232187, -0.0298168207982897, 
    -0.0545790130111923, -0.0502767601290563, 0.0169543042319664, 
    0.116333117893922, 0.144858062814083, 0.131229270858592, 
    0.0745783258877361, -0.00154554248611457, -0.00253267413207353, 
    -0.0049997289638512, -0.00832767143141807, -0.0108052498042783, 
    -0.00683418498639948, -0.0124292290337033, -0.0234196201948033, 
    -0.0311400509974457, -0.0359684654358679, -0.0253886944960691, 
    -0.0106907350669359, 0.00474065539103557, 0.0158480211295924, 
    -0.0019857149208606, -0.0388645495170534, -0.0516282385006743, 
    -0.0519909435350016, -0.0754972957684705, -0.079781131306371, 
    -0.0112833923725542, 0.124587354440976, 0.147755235207491, 
    0.124459765684401, 7.68072166739207e-05, -0.00400909648461009, 
    -0.00542221597472438, -0.00429510693372833, -0.0034663625989435, 
    -0.00337334322530977, -0.0097763964925327, -0.013999255105948, 
    -0.0122763989733017, -0.0309824018050673, -0.0360251561939782, 
    -0.0255550540543553, -0.00456198347167049, 0.00923305742001168, 
    -0.00924575319887842, -0.0324935521499557, -0.0553811879356959, 
    -0.092571155809548, -0.0723119045048706, -0.0388295974996164, 
    0.0296992232045436, 0.0905916911128568, 0.00204887774631173, 
    -0.00664674135985386, -0.00833723150903529, -0.0026443045377936, 
    0.00151841561814256, 0.0027323970665367, -0.000457383584164818, 
    0.00249360772334538, -0.00199953164785608, -0.0196016296481891, 
    -0.0250060522597753, -0.0205055264007138, 0.00172969381914913, 
    0.0110843984148026, 0.00438518688125227, -0.0193204974558199, 
    -0.0567802642962344, -0.0815025256955038, -0.0527677869237745, 
    -0.00034974881048135, 0.0509089901425514, 0.0767076529221483, 
    -0.00167614951542341, -0.0125502816808164, -0.0136417537577443, 
    -0.00821342798783786, -6.46934195444134e-05, 0.0083956127682767, 
    0.0108269729724917, 0.0107697717375844, -0.00841250765523044, 
    -0.0154139189618171, -0.00527401667296601, -0.0030838117275234, 
    0.0164818287793327, 0.0296457752658429, 0.0281500550671649, 
    0.0114304476768862, -0.0249262693304009, -0.0705113160977596, 
    -0.0709377389903205, -0.0543577663369967, -0.00998598863678194, 
    -0.0153891076905535, -0.00782630204150542, 0.00572624563802288, 
    0.00306402506693515, 0.0109628398101019, 0.0133683711984449, 
    -0.00198159641317828, -0.0206927986128153, -0.0267267540489941, 
    -0.00906028983680388, 0.00518743832481233, 0.0253526669985368, 
    0.0432363377032003, 0.0438563399694488, 0.0328689826844188, 
    -0.00616230472237645, -0.0449305047146374, -0.0675464971668309, 
    -0.00810510007069498, 0.00163675810978609, 0.0217319019531007, 
    0.0445771502301594, 0.0187022345887818, 0.0152366513449615, 
    0.00723372144485136, -0.0198872077377487, -0.0352539531944011, 
    -0.0464352901670943, -0.0365664533746285, -0.0111140614062492, 
    0.00627526704687054, 0.0306946396856911, 0.0357597683120182, 
    0.0365465863203626, 0.0218502467175809, -0.00124502645063524, 
    0.0150696840961415, 0.0335061502607096, 0.043080135732849, 
    0.0410613274527296, 0.0298806778104353, 0.00447496030401988, 
    -0.0312671967546805, -0.0535694770104856, -0.0701323899681978, 
    -0.0731146328768334, -0.0529040240004883, -0.0330091442002197, 
    -0.0242254674959423, -0.0121980039718745, 0.0233355439893022, 
    -0.00457934009810946, 0.00512893489448895, 0.0131019146329657, 
    0.0185457265208518, 0.0425432167361791, 0.0407278901560466, 
    0.00371109629601828, -0.0454883220181525, -0.0667717120064033, 
    -0.0907571262794418, -0.0930344620541249, -0.0791547705470429, 
    -0.0841488514786039, -0.0801473766099443, -0.0309864889122157, 
    -0.00949167988200174, -0.0103865367202421, -0.0136634530231694, 
    -0.0113300205215569, 0.00634268146397268, 0.026572029742578, 
    -0.0114001145396655, -0.0460481801039627, -0.0617451597263708, 
    -0.0975972286464301, -0.101271084547476, -0.0929334681231005, 
    -0.0911104622979937, -0.0876516285632269, -0.01707895157933, 
    -0.0235306165836043, -0.0351760813756058, -0.0316383159715508, 
    -0.0188397835860576, -0.00167298363505112, -0.028741076078886, 
    -0.0282634275910428, -0.0429496893036658, -0.0841517214679107, 
    -0.0909145817037919, -0.0697353317291694, -0.0235510079193944, 
    -0.0293903929463359, -0.0419496846459284, -0.0400391424598289, 
    -0.0307561119828788, -0.0157107166173105, -0.0207241178259553, 
    -0.0118297332733618, -0.0343947407903304, -0.0733936943619098, 
    -0.0851943176363519, -0.0641385012675962, -0.0314786017889861, 
    -0.0368957186854618, -0.0470988025296978, -0.0467122306531165, 
    -0.0397820526924877, -0.0334209004191362, -0.0235604525461461, 
    -0.0195378083897229, -0.0443881304278162, -0.0774262651184172, 
    -0.0845284650186253, -0.0551323077327592, -0.0339950063380101, 
    -0.0422759359609364, -0.0517983227623206, -0.0433420323587538, 
    -0.0190958267811687, -0.0351495691198013, -0.0327485974155821, 
    -0.0239980947844179, -0.035792273345462, -0.0714912868819972, 
    -0.0833602017497619, -0.031412866079, -0.0467049821631947, 
    -0.0525277180745058, -0.0260952408219816, 0.011743958964335, 
    0.00640141456625232, -0.0109793741586243, -0.00743529084085304, 
    -0.0224778976838466, -0.0658202816911261, -0.0743671044616815, 
    -0.0288812060837289, -0.0455601105552784, -0.0370492775097002, 
    0.00833638860519872, 0.0405573509924383, 0.0400891591911629, 
    0.00925391795125212, -0.00737248971966453, -0.0179599488113565, 
    -0.0496035238926846, -0.0569582962140048, -0.0295502437986857, 
    -0.0391152570103407, -0.0186254588832559, 0.0169909308208121, 
    0.0262287463211731, 0.021258761636517, 0.003636563570466, 
    -0.00940717000230746, -0.00739273190471248, -0.0154173036498627, 
    -0.0178357419148946, -0.0301412253188871, -0.0194323375618795, 
    0.00537212118344022, 0.00862242393937163, 0.00290730841118415, 
    -0.00704118251248416, -0.00981794961205366, -0.0049184514878712, 
    -0.00526608015469866, -0.0166200599953328, -0.0164252579138375, 
    -0.00098182901168627, 0.00375187031545143, 0.000936770202128781, 
    -0.00504745477968676, -0.00245500936947012, -0.00319215479454177, 
    -0.00167266570335989, -0.0129318258319151, -0.0152699116055383, 
    -0.00719132460112898, 0.000963601180595613, 0.00317965575507436, 
    -4.11703825898448e-05, -0.000387321338612753, -0.00525357811806353, 
    -0.0181290514840271, -0.0188570755295027, -0.0116888797480124, 
    0.000368210838538406, -0.00905113717618071, -0.0138274131100391, 
    -0.0130576067719807, -0.0111702567637104, 0.0275194350890226, 
    -0.015450344041293, -0.0153103411499433, -0.0129965177297422, 
    -0.00078712515346125, 0.0160447825168, 0.0186597758715017, 
    0.00316414228271283, -0.0115724486058388, -0.0128829201694039, 
    -0.00540977248061675, -0.0179253645400841, -0.00739583769822009, 
    -0.00520171975161639, -0.0102888528140418, -0.00972106022425084, 
    0.00839272072562335, -0.00902284725945642, -0.0105914218032903, 
    -0.00823384121012228, 0.00471076964876003, 0.00481285085479296, 
    0.00776008605521411, 0.019001421201585, 0.0298183722062962, 
    0.0299294416034073, 0.0390075676184443, 0.00105658624759106, 
    -0.000112402698724327, -0.000665694514823892, -0.00122260414009563, 
    -0.00243264987336668, -4.67128737366188e-05, 0.00272837326168464, 
    0.00200343112704378, 0.00196999638215141, 0.00193037809229351, 
    0.00178267048757663, 0.000278492707156097, -0.00235184598707008, 
    -0.0039403513430058, 0.000682877751391891, -0.000366746590150273, 
    -0.00107148251842871, -0.00163507790558471, -0.00320504931789987, 
    -0.00435972960512583, -0.00104745011747997, 0.00357150382918226, 
    0.0086382218858973, 0.001345147796071, 0.00128542924171454, 
    0.00115680352651835, 0.000432143979786632, -0.00109967762528735, 
    -0.00274060087743346, -0.00410404656198105, -0.00411411163944707, 
    -0.00362822319030658, 0.0128028483309819, 0.0164331313082528, 
    0.012689617625582, 0.00703759172383848, 0.00319045279334799, 
    -0.000576352125312588, -0.00546125651922615, -0.013763032464316, 
    -0.0145771361935667, -0.00721118366286466, 0.00517107930570088, 
    0.00630268374851145, 0.0111861537068683, 0.00978396468193023, 
    0.00326239048412197, 0.00032494509890357, -0.00790934248842374, 
    -0.0160193117677353, -0.0264088203683366, -0.0263967276165063, 
    -0.0393688037050638, -0.0153440328008889, -0.01845129881993, 
    -0.0138356237946182, -0.00472389962575095, 0.00123217375332215, 
    0.00998434503822589, 0.0321581490510027, 0.0383379834740756, 
    0.0343407287632171, 0.026500737048638, 0.0258251054266721, 
    0.0253129561909318, 0.0179773608524344, 0.0106797838055399, 
    -0.00829305317924332, -0.0372303529554375, -0.0569612018100132, 
    -0.0676328175678623, -0.0379332673998106, -0.0172001382030422, 
    -0.0112699581841051, 0.00713160445244045, 0.0225098897884182, 
    0.0225420947141304, 0.0255840606012125, 0.0194755271873576, 
    0.01141830736316, -0.0183020505264032, -0.0342842318611635, 
    -0.059778347560614, 0.0119006474002198, 0.0152024006953033, 
    0.0146346028826208, 0.00772882966045449, 0.00195719736629828, 
    -0.0012265542734313, -0.00941432062349631, -0.0182876603061853, 
    -0.0181819017789849, -0.0099266663222131, 0.0102494387379423, 
    0.0142319084451364, 0.0122644395308606, 0.0100589492978681, 
    0.00390883293420178, 0.00288822473878117, -0.00418532763054179, 
    -0.00655573867927312, -0.0135663831324153, -0.0283967288562545, 
    -0.0461906563883289, -0.0123960721993366, -0.000788489777894993, 
    -0.00586409613247293, -0.00284052379326423, -0.000819735137455452, 
    0.00449615172056249, 0.0328180302324548, 0.0398694093246921, 
    0.0305005041214167, 0.0283606672395468, 0.0255612045373301, 
    0.0183574107086532, 0.00704715133369283, 0.0114157134292412, 
    0.00380451563596544, -0.0205009872349739, -0.0490576756684775, 
    -0.0707645103168617, -0.0623226488588461, -0.0482555876640512, 
    -0.0310684213361126, 0.00219979419299884, 0.024934468119887, 
    0.0261402835395646, 0.0230924626652786, 0.0124590299359894, 
    -0.0021267615342487, -0.0349554720377343, -0.0466053877307458, 
    -0.0586316452752793, 0.00666335810294913, 0.00957559391294511, 
    0.00839549145263867, 0.0029615668706024, 0.00351082886838881, 
    -0.0017563160753009, -0.013523797044719, -0.0202353630292335, 
    -0.0202066181337241, -0.0133935677930022, -0.000318636245548972, 
    0.00304656718324639, 0.0130525309252466, 0.00803792634526955, 
    0.00556773674045941, 0.00855181751925643, 0.00817759405223349, 
    0.00993129255823663, 0.0141280122551018, -0.0358856978875022, 
    -0.0498264402453455, -0.00530106530563014, 0.00961484820348707, 
    0.00102121289555455, -0.00515126581863772, -0.00429419815853418, 
    0.0113876810733614, 0.0365086386867298, 0.0335056582471116, 
    0.0219352228588972, 0.0185470313495665, 0.0147351202662473, 
    0.00316357741585132, -0.00228757823708533, 0.00535766657709928, 
    0.0064283827980045, -0.00989880860095101, -0.0403588866739041, 
    -0.0662423184027192, -0.0636388858687975, -0.0458520709384398, 
    -0.0284340850405642, 0.00823413900806283, 0.031057339356627, 
    0.0343840626266007, 0.0123937715192943, 0.00640887399023234, 
    -0.00265133660787818, -0.0475706466367521, -0.0755728688807697, 
    -0.0737625660894113, 0.00406752951759171, 0.00241484802970826, 
    0.00124134118196829, 0.00269424736325589, 0.0148104235251958, 
    0.00999562475584795, -0.00431364300526067, -0.0116590245858825, 
    -0.0164076845139849, -0.0186242611620575, -0.0148117596699331, 
    -0.00536161725175397, 0.0104217723883733, 0.00455590803949232, 
    0.00650056430531585, 0.0099836053749006, 0.0133423870392048, 
    0.0215656460848951, 0.0146012607711186, -0.0188468953055038, 
    -0.00779485905047494, 0.0217514717855543, 0.016371153872445, 
    -0.000518680279259108, -0.0101100572625838, -0.00657710556669245, 
    0.0113083479578907, 0.0268584836474815, 0.0153528813851234, 
    0.00354392543439351, 0.0137011877198447, 0.00770467900294417, 
    -0.00231601829247459, -0.00649106548507602, 0.000975609136700331, 
    0.00373521026538574, -0.0116345541987268, -0.0352399138273738, 
    -0.0603729502844508, -0.0501094306967934, -0.0162196221612614, 
    -0.017348900254687, 0.0230193640868186, 0.0562110954618086, 
    0.0570838208141852, 0.0316159189279432, 0.0217441703490728, 
    0.011355415744344, -0.0326762872320134, -0.0707088851602557, 
    -0.0622474489360094, 0.0075143140839182, 0.00261298431966122, 
    0.000720078168540891, 0.00871262361204638, 0.0319426838085331, 
    0.0348431709317497, 0.0100798543180955, -0.00194489523429967, 
    -0.0166476593878052, -0.0280452283582166, -0.03027491416254, 
    -0.019302742160346, 0.00412672769099458, -0.000182285304402509, 
    0.00269108324493703, 0.00580804047860591, 0.00729426954559818, 
    0.0255628055477274, 0.0352670441041239, 0.0176142036246919, 
    0.0157816591730359, 0.0161093413447974, 0.00873909647803521, 
    -0.00575898655963715, -0.0132042691797512, -0.0100012831149936, 
    0.00501997961338954, 0.00392873828488084, -0.0277600982163556, 
    -0.0275057628896712, 0.0043223069317185, 0.000786910306468855, 
    -0.00342296076084166, 0.00478984065168933, 0.0196391052382142, 
    0.0315863444061797, 0.0173600006088339, 0.0109994023065821, 
    -0.0417586456355865, -0.0299382189526895, 0.00912165293219176, 
    0.0115194197244253, 0.0382756928728147, 0.0848889701682124, 
    0.0805973417343272, 0.0629427640535856, 0.0329032544775445, 
    0.00254381435398876, -0.0411110863954013, -0.0708058753806993, 
    -0.050739437762583, 0.0121990180518439, 0.00995158162345953, 
    0.00786128902047748, 0.0154130248675144, 0.0284721289691027, 
    0.0481177731045347, 0.030799695979272, 0.00569364701426749, 
    -0.0138599900972532, -0.0357782541968711, -0.0395064873063454, 
    -0.0225263901423796, -0.00556211449655084, -0.00798052942878366, 
    -0.0079730986560422, -0.00535606944356535, -0.00407209002445302, 
    0.016619100759896, 0.0170518747501979, 0.00514927296943583, 
    0.0110181051693845, 0.0165067080084515, 0.0045296933459733, 
    -0.0113831684159211, -0.0118877714210621, -0.008693681081939, 
    -0.00111677829385897, -0.0188917478769452, -0.0567443455142581, 
    -0.051318204193636, -0.00393025261784523, 0.00209509478159004, 
    0.00343532341545074, 0.0187057573130403, 0.0385981727655425, 
    0.0508339821108857, 0.0453344703155693, 0.0295269585604223, 
    -0.0221529172384437, -0.016635928839373, 0.0215320812182319, 
    0.037995658249005, 0.0507095855469091, 0.0891942410937664, 
    0.0780651140496717, 0.0621948903727955, 0.0390238614767951, 
    0.00413537844497346, -0.0302952600165958, -0.0497216490637996, 
    -0.0488424929555232, 0.0140360237337995, 0.0170028289403267, 
    0.0156519652991149, 0.0176761543581501, 0.0224796243760622, 
    0.0412680506122599, 0.0369063614572206, 0.0142628326446045, 
    -0.00956941601534018, -0.0397103379435682, -0.0441767652000579, 
    -0.0265430837706373, -0.0135430689922036, -0.0154089976580197, 
    -0.0201739122343756, -0.0243349156874186, -0.0182382651199346, 
    0.00261718006411312, -0.00720123569271801, 0.00715108161434572, 
    0.0185736716231818, 0.0243805374956499, 0.0119178383150474, 
    -0.0102904226941145, -0.0084945732538392, -0.0118229456410843, 
    -0.0183054701310666, -0.041168244814792, -0.0318264708706566, 
    -0.0620580536164327, -0.0125755133685199, 0.00826516058844572, 
    0.0124716991234701, 0.0291564696143353, 0.0485643639018603, 
    0.0413688285920408, 0.026303673350552, 0.020338405152714, 
    -0.00512309885646461, -0.0127925257540788, 0.00980689523139371, 
    0.0459663755991607, 0.0657358266115696, 0.0799526579054938, 
    0.0646605767203694, 0.0657078455988932, 0.0737570041336911, 
    0.0309239982614513, 0.00482726264042417, -0.0053715672193343, 
    -0.028187044381026, 0.0110985564035164, 0.0126868291524613, 
    0.017788350548921, 0.00676262341723369, 0.0136749809345635, 
    0.0264631237818887, 0.0395030668159039, 0.0235763017749382, 
    -0.00402872911916823, -0.0363250899080169, -0.041277116691169, 
    -0.03072752573548, -0.0202169552949542, -0.0194943488747693, 
    -0.0236203996953897, -0.0324848625911605, -0.0292197959482672, 
    -0.00796883788199505, -0.0111691124019228, 0.0104013538016779, 
    0.0285907775718887, 0.0314635990598565, 0.0186338661040807, 
    -0.00435847713828003, -0.00945014545455703, -0.0191957821108209, 
    -0.0224763370604669, 0.00187314301810396, -0.00540632207768953, 
    -0.0153530945568744, -0.0087850601999293, 0.00491335029226408, 
    0.0154057841881426, 0.0324692007639873, 0.041709479765067, 
    0.0272130866064671, 0.00697399286289181, -0.00194692523228734, 
    -0.00451682271387573, -0.01489438040729, -0.00717598736595517, 
    0.0206991006125327, 0.0482137672489031, 0.0540675297706107, 
    0.0420664861566202, 0.0365439576614748, 0.0610913748329797, 
    0.0543865551540287, 0.0361274138138433, 0.0414046068240281, 
    0.00462399841097702, 0.00358662400694561, 0.00643348151960942, 
    0.00716328342591015, 0.00285377973512684, 0.0024595447959244, 
    0.00715925155809197, 0.0164571733125317, 0.0244431582776099, 
    0.00325335872737399, -0.0344991493345949, -0.0371847398685277, 
    -0.0291439684191628, -0.0204729460216894, -0.0212020451783615, 
    -0.0225020117440482, -0.0271837575640448, -0.033425645019433, 
    -0.0210127351050879, -0.00493252395088929, 0.0094023918395456, 
    0.0253718244741573, 0.0273181859283768, 0.013784938690907, 
    -0.00111603755505764, -0.0109867137849122, -0.0223511261472378, 
    -0.0206251082555562, 0.0270130732267461, 0.0244604869266383, 
    0.0265255980360071, 0.0126506356375083, 0.0071623950478045, 
    0.0138961132793896, 0.0282664393725701, 0.0336855999496124, 
    0.0304636998101253, 0.0114061848825735, 0.000595238936169242, 
    -0.0133517769503387, -0.025581779890742, -0.0145512564935654, 
    0.00951719675305487, 0.0265242970772593, 0.0328111280398661, 
    0.0290615176485742, 0.0228343262680341, 0.0478256122886361, 
    0.0668039362708531, 0.0422087184571, 0.0530729874161603, 
    0.0137281592240804, 0.00289999241590856, -0.00029173357001305, 
    -6.09094632275665e-05, -0.00267521410880872, -0.00234152889344493, 
    -0.00573347660838137, 0.0016231894367178, 0.0190075979568475, 
    0.00494329917340309, -0.0305786355943248, -0.0348948073414764, 
    -0.0256908645953897, -0.0181340882312891, -0.0152747283052024, 
    -0.0196063566441032, -0.0305437121348242, -0.0369971614028526, 
    -0.0368453569880986, 0.00281419940969908, -0.00492073730923765, 
    0.00254361523747403, 0.00597480648234873, 0.00203585950420525, 
    -0.00301155286977442, -0.0141060354989204, -0.0246742814736783, 
    -0.0237042848030796, 0.0185603297899686, 0.0463360538754512, 
    0.0408971516442983, 0.0205795240350741, 0.0153639466466159, 
    0.0127901690264918, 0.0216758064648779, 0.0236454730199163, 
    0.0250259335882227, 0.0132938810089297, 0.0159691192262795, 
    -0.0147615701520974, -0.0250836595111992, -0.0172041513889409, 
    -0.00291552918554062, 0.017221953308729, 0.0338686632821374, 
    0.0309503749660143, 0.0250621267479354, 0.0439761950743746, 
    0.0776206467448372, 0.0692474374793615, 0.069506621505277, 
    0.0379698171079339, 0.00418198597986479, 0.00171205674997459, 
    -0.00168794510831637, -0.0035894900653406, -0.00440887575234762, 
    -0.0104257602464863, -0.0103629174355676, 0.00438947243481737, 
    0.00653323027667487, -0.0201105406275419, -0.0303294083705763, 
    -0.0236510095502994, -0.0214952696993347, -0.0219572404037828, 
    -0.0218923928244906, -0.0327257889029278, -0.0327161998184844, 
    -0.0192034290679899, 0.00429837668306374, -0.0215701625495317, 
    -0.0221709299253036, -0.0108616981984505, -0.00661765024143121, 
    -0.00407292699971052, -0.0111193673330494, -0.0252515288927594, 
    -0.0213312461914573, 0.0243889032238178, 0.0545978364811707, 
    0.0429920191344374, 0.0135572789261756, -0.00768503833442793, 
    -0.00580649676244465, 0.00706125916000313, 0.00681705262735321, 
    0.0104489886393246, 0.0160429395100395, 0.0179279968517565, 
    -0.0150765374981226, -0.0333247878212231, -0.0167080351073114, 
    0.012307852391161, 0.0405180884755099, 0.0365719288701844, 
    0.0321391197991712, 0.0434965773325601, 0.0705395369705015, 
    0.0911580539893319, 0.0988771498793674, 0.0781504060804055, 
    0.0519375708263939, 0.00678319451957826, 0.00347430200754506, 
    0.00397029729372583, 0.00393206221525261, -0.00432650993147803, 
    -0.0105303284601562, -0.0179532900433046, -0.00537287332381075, 
    0.00383741159340242, -0.00759378410651246, -0.0179046590832172, 
    -0.015305102662819, -0.0142870533993878, -0.0186048148286773, 
    -0.0219559501492088, -0.0317127525987842, -0.0322032003575197, 
    -0.00730034830452099, -0.000782343620078069, -0.0281747810177386, 
    -0.0306646397997902, -0.0153812596276152, -0.00459166814946604, 
    0.00152956556455495, -0.000113660100631023, -0.019570633872161, 
    -0.00655425079174033, 0.0327852334803935, 0.0557866985009753, 
    0.0522874845070565, 0.0196647031810109, -0.0164487543392876, 
    -0.0279331819096001, -0.0167270833622286, -0.0166749103481213, 
    -0.011556277576853, 0.00631940146531015, 0.018374572519149, 
    -0.00927707572903206, -0.0327125095707294, -0.0149474876031037, 
    0.0143892380588363, 0.0362132133425768, 0.03234958109757, 
    0.0401800850150889, 0.0620762439822972, 0.0935586178615282, 
    0.102652413506364, 0.109264973580894, 0.0927802612550892, 
    0.0529654883479437, 0.0082313837306419, 0.00744538954604356, 
    0.00925461099802745, 0.0100008900249169, 0.000405352948057786, 
    -0.00545110654341324, -0.0190603634834275, -0.0107173405121931, 
    -0.00198724709917439, -0.00627934914854562, -0.0111121864230184, 
    -0.00970961748587714, -0.0101915841231901, -0.0119465466929689, 
    -0.0165207693163187, -0.0268835156244378, -0.0306531021807265, 
    -0.0135451584622629, 0.00572891963916221, -0.0114947403410253, 
    -0.014662865100962, -0.0141948917938338, -0.00995689471624472, 
    0.00083507933931898, 0.00850649605323021, -0.00342995888835605, 
    0.0150445916499444, 0.0416882825381001, 0.0523927950617295, 
    0.053913291064563, 0.0158262893449779, -0.0127858996933218, 
    -0.0504570971630082, -0.0464850495723148, -0.0436869255106341, 
    -0.0350080305739143, -0.0167001141094461, 0.0118178615870363, 
    0.00101930183108039, -0.021415633455972, -0.0117685129923573, 
    0.00877236136310563, 0.0220882747913344, 0.0175558848545312, 
    0.0275343758508988, 0.061168412996335, 0.0775153769694999, 
    0.105970421390416, 0.102711934092057, 0.0906713586072919, 
    0.0504176971458954, 0.0067205892132708, 0.00610568752224735, 
    0.00863566168836446, 0.00807104921430327, 0.00784538906339811, 
    0.00345039127252423, -0.0161742176893415, -0.0120613901095376, 
    -0.00302866854711718, -0.0037262649791415, -0.0102319582574557, 
    -0.0102732966031301, -0.00962282177236429, -0.00898378131714697, 
    -0.0140970655914966, -0.0190429828256277, -0.0225109775170308, 
    -0.00656141363300918, 0.0119622050486564, 0.0127900206428409, 
    0.00783940790615438, -0.00507791331799505, -0.00799885523080437, 
    0.00402417296860876, 0.0138042955484907, 0.0154280576715931, 
    0.0307397073651113, 0.0386377699541541, 0.0463590772894522, 
    0.047775357133578, 0.00137274427465753, -0.0340548502834507, 
    -0.0753033366013621, -0.0744857756257735, -0.0562817821380531, 
    -0.0428536954870401, -0.0255846771177438, 0.00776761270366889, 
    0.0181607059868058, 0.00905896752090931, 0.00188293520749302, 
    0.00963462349393275, 0.0386994201957126, 0.0756166791383854, 
    0.0824048600154837, 0.064171157506996, 0.0463499318313911, 
    0.000407392093102377, -0.00171543648544116, -0.00703096630220622, 
    -0.0133166171977154, -0.000710398767622828, 0.00587160568711912, 
    -0.00356636412782522, -0.00732651824732336, 0.00730427423467322, 
    -0.00911785458319704, -0.0225232303602221, -0.0223746077727014, 
    -0.00932689874742797, -0.00756184193332628, -0.0120382529443011, 
    -0.011754515948621, -0.00698197998365319, 0.00425290575203526, 
    0.0151017262449316, 0.0222706856466878, 0.0223568484383152, 
    0.00512019086845092, -0.00859487589249044, 0.00865644416419101, 
    0.0198489792543703, 0.0213088300023684, 0.0242375262508162, 
    0.0342358712999953, 0.0389571311651702, 0.0319852285202298, 
    -0.00101162102841136, -0.0340525381058959, -0.0715927149627602, 
    -0.0624922124850011, -0.0520128214765316, -0.033251721117001, 
    -0.028004913725409, 0.0136550918462444, -0.0011804618687984, 
    -0.0132671620978765, -0.0109186066390111, -0.000299229949142841, 
    0.0270847849206062, 0.0474402203004205, 0.0349182017505012, 
    0.0332870506559228, -0.00719654722925159, -0.0123135838667409, 
    -0.0276509921509918, -0.037252653315823, -0.0223302059558721, 
    -0.00223293633888167, 0.00720331746265841, 0.00338915729172237, 
    0.0152298419368916, -0.0161762355174275, -0.0421895769277306, 
    -0.0356723518230772, -0.00602558737191074, -0.00805408673298851, 
    -0.0136441730479974, -0.00668076177173641, 0.00304652618828626, 
    0.0103344244683919, 0.0179033634777298, 0.024845953470556, 
    0.0279161029419158, 0.0265407755851237, 0.00837102770415844, 
    0.028816098517187, 0.0407107339052151, 0.0280397185885289, 
    0.0247150935297689, 0.0383737430098026, 0.0254735000219565, 
    0.0232267170353276, 0.0121954522569055, -0.0471407377268875, 
    -0.0311039350274055, -0.00844404143336849, -0.0181881679606327, 
    -0.0104898844583473, -0.0105739940078828, 0.0036855444563562, 
    0.0129817930533577, 0.00915841165886431, 0.0134013537765165, 
    -0.013252129272815, -0.0229577788233153, -0.0441232695151897, 
    -0.0533846078964767, -0.0360728177456733, -0.0120435078554524, 
    0.00403845115978231, 0.0104127537362452, 0.0194636085542223, 
    -0.00763846009949291, -0.0370651019695369, -0.0332512055720357, 
    -0.0023381541951229, -0.00920859279550463, -0.0128718576310739, 
    -0.00358839211647315, 0.0063793854601595, 0.0124992607004313, 
    0.0182738434765293, 0.0194500792170122, 0.0237956120158261, 
    0.0453210144252167, 0.0432427789514976, 0.0756473987728032, 
    0.0624467442798292, 0.0458461551778421, 0.0538102248269793, 
    0.0438765492965938, 0.0267256270814906, 0.0111597378398305, 
    0.000123856847014114, 0.0192616806108263, -0.0227606205416934, 
    0.0014724888867141, -0.00494914907119347, -0.00938750376715823, 
    -0.0082786442952605, -0.00227819352582926, -0.0105426368067811, 
    -0.0136830803948912, -0.00887208721555331, -0.00856681037890865, 
    -0.00893111699570747, -0.0248197270289509, -0.0486827508984497, 
    -0.0442822383690874, -0.0209030185246952, -0.00603078842137916, 
    0.00746839742231889, 0.00922137577276272, -0.0137173556199875, 
    -0.0360880535916041, -0.0238784772439559, 0.000178759989525479, 
    -0.0190825270072989, -0.0247860822808853, -0.00955623969846873, 
    0.0013406431859151, 0.011677691031586, 0.0116509033219886, 
    0.00675843200154501, 0.0144685941233125, 0.0696687162554213, 
    0.0942618231335083, 0.124329759100194, 0.0888572441128162, 
    0.0615576077842493, 0.0618255704320499, 0.0338736103149769, 
    0.0138457207750097, 0.018597094657779, 0.0192025603509168, 
    0.0192616806108263, 0.00831164484821362, 0.000920472178626135, 
    -0.00600964385026229, -0.00722015756518257, -0.00656491286148152, 
    -0.0215003792543803, -0.0210135636202031, -0.0079255232279946, 
    -0.00405022841160003, -0.000994754542053304, -0.00328812140087814, 
    -0.0231124939251479, -0.0380270150298341, -0.0205746772521207, 
    -0.0055428626781629, 0.000436845081895836, -0.00682170129658567, 
    -0.0270501583966611, -0.0394605356008928, -0.0152773648583908, 
    0.00679487678499105, -0.0102616857586944, -0.0336380720818386, 
    -0.031305523061025, -0.0183044939750999, -0.00673495382710083, 
    -0.0125217680403112, -0.0173540569670299, 0.00677070096768501, 
    0.0795217546959291, 0.136740091822143, 0.1357215198004, 
    0.0874736326062566, 0.0759570235207383, 0.06502913853431, 
    0.035616039323398, -0.0033934350392687, -0.00585090559299326, 
    -0.00655979105964695, -0.0211260735536414, -0.00255103487930843, 
    -0.00118307920535475, -0.00234217024292302, -0.0103517944317908, 
    -0.0224584737380551, -0.0177024787535376, -0.00662565532827319, 
    -0.0145906917761599, -0.0251343861344687, -0.0327043230941285, 
    -0.0325979410998924, -0.0100254502629045, 0.0178939809639228, 
    0.0187650176943096, -0.00943204912353045, -0.0397734416764733, 
    -0.0310301667456716, -0.0258381791991676, -0.0499855936081137, 
    -0.0571986564288387, -0.00266667500130411, 0.0992545357226099, 
    0.141930564902665, 0.132595409933371, 0.0817052736246357, 
    -0.00188357743537337, -0.00312742240111613, -0.00489678476597774, 
    -0.00788292661513704, -0.0109853161941018, -0.00892541027875276, 
    -0.0145890401471326, -0.0260414808598861, -0.0300960518567528, 
    -0.0333299489736994, -0.0233637612490654, -0.00783477816924506, 
    0.00463752673120286, 0.0138101480580311, 0.00197996048954653, 
    -0.0339593107088243, -0.048603584568792, -0.0491003604918359, 
    -0.0678067085746868, -0.0815138804873369, -0.0388255814984436, 
    0.108105723267919, 0.147050575192368, 0.120301863795371, 
    5.57163654696293e-06, -0.00424814457793934, -0.00545183675256468, 
    -0.00393081424371508, -0.00469520292446278, -0.00613601411727611, 
    -0.0136666382919076, -0.0165487810946258, -0.00951041968376994, 
    -0.0285274429271107, -0.0320345312375711, -0.0207182726063283, 
    -0.00479023151099038, 0.00922617999354573, -0.00865338968448534, 
    -0.0299055507978351, -0.051851785947818, -0.0918475641583077, 
    -0.0659443068246157, -0.0334094036854208, 0.0161982052967629, 
    0.0895952723069557, 0.00182810185860088, -0.0068653843385873, 
    -0.00821724746526028, -0.00133144253478664, 0.00108219356607376, 
    -0.00121025426327461, -0.00647960792194922, -0.000233854372007205, 
    -0.00315394009054549, -0.0180863104843786, -0.0224341163047035, 
    -0.0201859450922384, 0.00277840792584509, 0.011367569886541, 
    0.00503172716280129, -0.0197500983296369, -0.0601357560295251, 
    -0.0780315947573565, -0.0388768499711245, 0.0170678883551574, 
    0.0551036540422312, 0.0775311626872967, -0.00269664790395226, 
    -0.0128293209745384, -0.0128030016627743, -0.00832971252246472, 
    -0.000638908009287298, 0.00588322896897686, 0.00540978691307335, 
    0.0108902408160909, -0.0103813251220628, -0.0155280747584604, 
    -0.00266004799607931, -0.00218223174343919, 0.0198488213983175, 
    0.0319116965694774, 0.029046146408334, 0.0131627260842316, 
    -0.0286617710373165, -0.0705131860137361, -0.0701718088432905, 
    -0.0476735469161481, -0.0113832548630147, -0.0135172612584363, 
    -0.00374848863320508, 0.00746169341099235, 0.00118932938810291, 
    0.00916026258662488, 0.0126429006227724, 0.00368746337878717, 
    -0.0209410624697076, -0.0296025852366231, -0.00853053232775489, 
    0.00868314349488605, 0.0265977736589409, 0.0425433440242539, 
    0.044969365273449, 0.0320949690460489, -0.0045266952084375, 
    -0.0417397707685099, -0.0618029536223104, -0.00627161310786416, 
    0.0079324687991406, 0.0290441303975929, 0.0469872782725788, 
    0.0159960654087696, 0.0132405546459396, 0.0109421944658999, 
    -0.0128092117025386, -0.031937890465419, -0.0483951690621848, 
    -0.0413895915140284, -0.0124619118004737, 0.00310756703015654, 
    0.0244136590233284, 0.0296598811856853, 0.0343205383156539, 
    0.0228519405052135, 0.00167571648928136, 0.0176212198629917, 
    0.0297314210312193, 0.0318796105136713, 0.035141731659206, 
    0.0255450771839177, 0.0101767110400185, -0.0210083532920597, 
    -0.0470727647544277, -0.0679928222523704, -0.0749026758848411, 
    -0.0576427784126955, -0.0383022376804794, -0.0315317721478384, 
    -0.0219693539512942, 0.0159803770832575, -0.003696675505524, 
    -0.00137150677496884, -3.74219335603102e-05, 0.00568267128615313, 
    0.0425879115466891, 0.0406529341094391, 0.0163514668171301, 
    -0.0291535651149026, -0.0599840451390911, -0.0861664122818378, 
    -0.0947375752537718, -0.0807153223866156, -0.0850204309430759, 
    -0.0860995018189225, -0.0396914723904302, -0.0106686869495175, 
    -0.0186253702410875, -0.0258101823167729, -0.0235619482755255, 
    0.00109902120030821, 0.0329386282427133, 0.0103769263983747, 
    -0.0340802351617308, -0.056647932483425, -0.0936961569522142, 
    -0.102817212987843, -0.0948531853351016, -0.0904089672014072, 
    -0.0883029079910348, -0.0181864950003632, -0.0265018214533613, 
    -0.0386408439426552, -0.036850311478373, -0.0204505289321319, 
    0.0136550332118881, -0.0170903377029351, -0.0298428335066809, 
    -0.0392844724447549, -0.0826884035106959, -0.095953285597031, 
    -0.0778540289559931, -0.0238114765361401, -0.0302865093959929, 
    -0.0415060762518454, -0.0413697982706129, -0.029935523810573, 
    -0.00444141505464476, -0.0212242780499696, -0.0131769174792596, 
    -0.032348213631755, -0.07269304013597, -0.0918750230325262, 
    -0.0768010966024683, -0.0306612072523872, -0.0378888872187086, 
    -0.0471547528455138, -0.044838654130548, -0.0346574912098389, 
    -0.0232351077230511, -0.0201011705524105, -0.0162817457135128, 
    -0.0416554435898281, -0.0793783459016295, -0.0905912198703666, 
    -0.0622744414736518, -0.0321202045840913, -0.0429852067873637, 
    -0.0514719005780817, -0.0371273270394001, -0.0148416689577499, 
    -0.0355242399007912, -0.029795032512114, -0.0221305267740898, 
    -0.0265731847250768, -0.0683142451293984, -0.0856775302140503, 
    -0.0305892221127973, -0.0449423462233471, -0.0486888779471562, 
    -0.015750874019129, 0.0193961396430662, 0.00147010622855225, 
    -0.0154805299745481, -0.00569161121681714, -0.0138323101470431, 
    -0.0601001764043958, -0.0750174606921586, -0.0286493887664333, 
    -0.0452110414667074, -0.0287363512024866, 0.0217877642815158, 
    0.0448938486337153, 0.0390945736389724, 0.00905914529465221, 
    -0.00414242134270819, -0.0136542438074651, -0.0469284407162887, 
    -0.057236362116914, -0.0319726525867227, -0.0345186274128623, 
    -0.008633737718377, 0.0220724957282351, 0.0241219961805006, 
    0.0186601790619964, 0.00757548688004357, -0.00702631487844509, 
    -0.00570560345466444, -0.0160133377646671, -0.0230938896102376, 
    -0.0300396269402365, -0.016151956810541, 0.00622229463938042, 
    0.0073425012601865, 0.00377036323935396, -0.00406723831231907, 
    -0.00638948589811802, -0.00280007228833936, -0.00736465038038016, 
    -0.0157750202369211, -0.0159962871726602, -0.00129591049674853, 
    0.00535981378399521, 0.00240534430940441, -0.00284015275037584, 
    0.000365478557537923, -0.00118506496973186, -0.000108327532655536, 
    -0.0108061881219819, -0.0147452790945193, -0.00805749973927781, 
    0.000613079865692656, 0.00369233649671585, 0.00196420471139804, 
    0.00109279279899831, -0.00415191788225323, -0.0177057457062547, 
    -0.0190113113737106, -0.0141403938438814, -0.000296816044061772, 
    -0.00810459906996503, -0.0112334994104617, -0.0120998893418018, 
    -0.0133941047074377, -0.00380006579728723, -0.00538305207505429, 
    -0.00648485293896903, -0.00793154960216934, -0.00891703120079369, 
    -0.00235539664261422, 0.012828251853988, -0.00459656092204621, 
    0.0188316785773089, 0.00023784934756851, 0.000158234773162403, 
    1.41730825151717e-05, -0.000824254665866152, -0.0032759606947799, 
    -0.00637358744427489, -0.00731911092026709, -0.000254815275514717, 
    -0.00520650987762456, 0.0316769078871881, 0.0298282775899446, 
    0.0275935458830989, 0.0196499064884754, 0.0018172071563311, 
    -0.0226650059963922, -0.0438632789104233, -0.0195600833104082, 
    0.010122787530335, 0.00481899023803944, -0.00809265456397766, 
    -0.0128611952115703, -0.00400890544775553, 0.00539863758846812, 
    0.0097026374963774, -0.00033635129711107, -0.000287331780476874, 
    -0.00014363960803333, 0.000350322007553322, 0.00143600790209114, 
    0.00257016581271709, 0.00407916643092403, 0.00242901097151264, 
    -0.0031702353892736, -0.00248400592598298, 0.00499777202091538, 
    0.00507136811492454, 0.000516567453760777, -0.0023000831350506, 
    -0.00398843038766028, 3.52833042918999e-05, 0.000153807251760707, 
    -1.13236700795415e-05, 0.000177424273580186, 6.24414854882071e-05, 
    0.000111427360299987, 4.84704444380315e-05, -3.20490906204464e-05, 
    -1.2689048354568e-05, -0.000365102171731211, -0.000205276049929494, 
    -0.000109645816839928, -0.000213761420313626, -0.000227889009557918, 
    -0.000392456970149639, -0.000297850470763114, -0.000152009599610536, 
    -0.000154660244449684, -0.00024398480157139, -0.000374533714248185, 
    -0.000240707171808502, -0.000361929196221472, -0.000149281523567453, 
    -0.000177339446052449, -0.000307727894882926, -0.000368362563128193, 
    -0.000230822828630256, -6.96392069159083e-05, -0.00024536480601124, 
    -0.000259278051044483, -0.000246176024280063, -0.000481976361800194, 
    -0.00019086451200277, -3.98892649991304e-05, -0.000329676482292816, 
    -0.000145980746366846, -0.000136030621533574, -0.000531520894104355, 
    -0.000202582858002925, -6.33851559849362e-05, -0.000145450413312089, 
    -0.000378895125715102, -0.00013585079916989, -4.29891945499635e-05, 
    -0.000479795852368762, -0.000175911842594023, -0.00013746201617966, 
    -6.54757513885355e-05, -0.000397701796190541, -7.49416749664025e-05, 
    -4.36582532087739e-05, -0.000125242457184629, -0.000394407093941916, 
    -0.000167086249517442, -0.000155938830875121, -7.06229333869721e-05, 
    -0.00039410840606806, 2.34213157536796e-05, -0.000115550744665772, 
    -9.06637466579455e-05, -0.000303358063595298, -0.00019361780623984, 
    -0.000134922791681646, 3.25970671317002e-05, -0.000259248085763168, 
    -0.000368153785059076, -6.03988253181687e-06, -0.00012624667212328, 
    -6.34008974246635e-05, -0.000217489692792227, -0.000247902895675972, 
    -7.64707875717018e-05, 0.000130226125321585, -0.000216817955231565, 
    -0.000338911180963664, -0.000117433074272558, -0.00010731451242128, 
    5.04511437871674e-05, -0.000151753293723521, -0.000479388826801867, 
    -0.00034196482123897, -9.5871214838825e-05, 4.59211602289182e-05, 
    -0.000172399624106104, -0.000282589196882527, -0.000255639621896268, 
    -4.1231418041097e-05, 2.25895092429651e-05, -1.78050393863156e-05, 
    -0.00044096231479464, -0.00037942085325148, -0.000143628107411225, 
    -0.000129123619918295, -7.80256683783406e-05, -0.00027337732605584, 
    -0.000552909517503363, -0.000390169318846557, -1.81162586254737e-06, 
    -0.000124672061195987, 0.000137779737867611, -0.000341323814009181, 
    -0.000424150002903149, -0.000149505024763343, -0.000308708312273323, 
    -0.000140921338107518, -0.000196593610304857, -0.000612693978817788, 
    -0.000486023876192254, -9.70273879009505e-05, -0.000334239130735154, 
    0.000171789301827474, -0.000260246586378714, -0.000433444166908791, 
    -5.63414219901256e-05, -0.000466374539888781, -0.000431457821075749, 
    -0.00026445876712471, -3.59459609181879e-05, -0.000513395579360911, 
    -0.000538982993989842, -0.000134088365729468, -0.000477089251364577, 
    8.9366612753695e-05, -0.00027075168368198, -0.000424678514832509, 
    6.03177314025119e-05, -0.000620063841136608, -0.000536871505215361, 
    -0.000476524188230129, 0.000165538545689951, -0.000418851949252742, 
    -0.000524418916576768, -7.28084981553844e-05, -0.00035121039577482, 
    -0.000495608374764462, -4.83771620379764e-05, -0.000347007791676251, 
    -0.000371597689494057, 0.000203174580296783, -0.00059635863596221, 
    -0.000589563321074743, -0.000583958237086751, 0.000149938013158753, 
    -0.000375927059039775, -0.000528364946678734, 6.16787101293204e-05, 
    -0.000568750907118967, -0.000464527033230498, -0.000166130239899486, 
    -0.000538929442389189, -0.000181131578624659, 0.000267167438236234, 
    -0.000541175524570889, -0.000578433994106001, -0.000294709369306, 
    -0.000568806238635162, -2.23431389184738e-05, -0.000437759625773047, 
    -0.000519025963115481, 0.000182333011898819, -0.000707236048429981, 
    -0.000458714088616116, -0.000234178757653977, -0.000643176544563052, 
    -3.5740629751034e-05, 0.000220650889074839, -0.000526143568694435, 
    -0.000581399936145199, -0.000574891324826365, -0.000427316000775003, 
    -0.000196268760027314, -0.000540947265011995, -0.000462372750404243, 
    0.0001735003200469, -0.000785078914968647, -0.000577597410551377, 
    -0.000266470056040895, -0.00026118422239581, -0.000672425593685422, 
    7.84985746827231e-05, 9.3239763808337e-05, -0.00055703354270173, 
    -0.000627114458925831, -0.000807480926791471, -0.000322570011586395, 
    -0.000301846345063691, -0.000613367591336351, -0.000317427342453827, 
    -1.97402098150372e-05, -0.000795100131849231, -0.000703833427949915, 
    -0.000280122667322366, -0.000605721606875707, -0.000508554003343059, 
    -0.000184670937805901, -7.61614559202717e-06, -0.000592645972620378, 
    -0.000634051665308833, -0.000849586838197811, -0.000526650570657568, 
    -0.000332975545856796, -0.000273815557953317, -0.000653210601696342, 
    -0.000148337479561274, -0.000256387334379808, -0.000760798962644263, 
    -0.000861345601910931, -0.000266590969299481, -0.000820712232817117, 
    -0.000355264693880155, -0.000332745353437689, 0.000114806064080952, 
    -0.000612736104322636, -0.000555855023721135, -0.000838846198398667, 
    -0.000731752969256527, -0.000346218535638738, -0.000538519888067864, 
    -0.000528579430664304, -0.000179771322046329, -0.000368324368300897, 
    -0.000683712894953724, -0.000909936586511416, -0.000223194364400131, 
    -0.000810153485720889, -0.000466841533428369, -0.000381664118494812, 
    -0.000312968091440602, 0.000170091826843088, -0.000618440106397183, 
    -0.000454413317457163, -0.000783792753521709, -0.000889948209559202, 
    -0.000343850576483328, -0.00070367970976762, -0.000400938213735222, 
    -0.000206302776315118, -0.000108449495107139, -0.000619034917057168, 
    -0.000910867669888277, -0.000264891592778861, -0.000773755266315711, 
    -0.000578847257336765, -0.000391316542256264, -0.000475839686267036, 
    7.31846842764698e-05, -0.000529752589853627, -0.000394336364521128, 
    -0.000649571645613419, -0.000876613175935174, -0.000310622614493959, 
    -0.000703145193131083, -0.000325924279959988, -0.000282223428026001, 
    -0.000365284349777302, 0.000116263578963999, -0.00060460550142309, 
    -0.000817506859487439, -0.000420919358245623, -0.00072273010716831, 
    -0.000678811879305592, -0.000417318472998208, -0.00057077950808577, 
    -6.2087127724598e-05, -0.000392374846927456, -0.00034672949501141, 
    -0.000636106129404435, -0.000834708856305299, -0.000237792966426079, 
    -0.000707682503460307, -0.000289254731359325, -0.000317379988252214, 
    -0.000464491390210248, 5.74382528612678e-05, -0.000449732901877247, 
    -0.000763937375866289, -0.000490037415954565, -0.000707682015527112, 
    -0.000606419932797507, -0.0004632072741422, -0.000600187868501308, 
    -0.000131974481786436, -0.000298335354291911, -0.000304132495184692, 
    -0.000299272866317809, -0.00055621650328445, -0.000743120880765991, 
    -0.000232217083768171, -0.000705598071682127, -0.000293295717542475, 
    -0.000381923892418348, -0.000512140904750135, -6.8838021356201e-05, 
    -0.000353921965851691, -0.000645856887824598, -0.000511232538726263, 
    -0.000655051762639657, -0.000577171723371498, -0.000401914670680096, 
    -0.000562391536910414, -0.000162846988210023, -0.000166552965962404, 
    -0.000285121600887483, -0.000374372903001393, -0.000387081399894848, 
    -0.000594092642052477, -0.000276838968967494, -0.000668400685496237, 
    -0.00032706810889747, -0.000470562145103732, -0.000528994829448581, 
    -0.0001266952463422, -0.000122149897177968, -0.000543901356081648, 
    -0.000248983805904829, -0.000454715242061745, -0.000470809305512923, 
    -0.000593547823227547, -0.000239663854402288, -0.000432536223499104, 
    -0.000161730081047078, -0.000140044635734815, -0.000366767971537891, 
    -0.000462083133277197, -0.000297038465667887, -0.000452773364491123, 
    -0.000336335629769535, -0.000590624404992465, -0.000434851587955851, 
    -0.000488600357057816, -0.000461035051538279, -0.000146915884425878, 
    0.000140529383076143, -0.00042179865204477, -0.000313219423838123, 
    -0.00035538592586833, -0.000425798161001411, -0.000401126317017434, 
    -0.000204748712704451, -0.000403622395899629, -1.07141720580022e-05, 
    -0.000160590601900297, -0.000430841657432317, -0.000545884628946866, 
    0.000140200775654962, -0.000431157531636978, -0.00011528771223538, 
    -0.000342490760888407, -0.000513393478412608, -0.000588849494674811, 
    -0.000324610282030992, -0.000391058069254056, -0.000132559912107045, 
    0.000279187638409311, -0.000366133389115143, -0.000378449532622894, 
    -0.000222216919798913, -0.000169370963368646, -0.000270425402734961, 
    -0.000265158775057896, -0.000426913335091547, 0.0003548338927251, 
    -0.000394818550090573, -0.000394183449826114, -0.000503229004988157, 
    0.000424702612060486, -0.000441881397413265, -0.000114040339809834, 
    -0.000317291359649345, -0.000516588006357062, -0.000469369311706276, 
    -0.000156832351955827, -0.000378908556203026, 0.000117909221735583, 
    0.000239824709390642, -0.000233272162257628, -0.000452559176629442, 
    -0.000124400744061603, 0.000377617736725825, -0.000277576778075669, 
    -6.5290796435185e-05, -0.000218781541520397, -0.000537652763460228, 
    0.000431458571387539, -0.000690821581522462, -0.000201854720440813, 
    -0.000409048165565249, 0.000727317838921503, -0.000349429829260176, 
    -8.55378821518238e-05, -0.000220256680359038, -0.000220948510894071, 
    -0.000344419556839926, -0.000119278606659744, -0.000402195991667733, 
    0.000552508265286207, -0.000263834522776431, -0.000112272363297714, 
    -0.000435156177182347, -5.73466583636618e-05, 0.00105805081363903, 
    -0.000420648066209472, -2.52604177431084e-05, -0.000241369756128926, 
    -0.000842623146060887, 0.000106391127381893, -0.000663447689667465, 
    2.23227734541264e-05, -0.000301589994381497, 0.00060954213500827, 
    -0.000170946112762948, -9.20161714467473e-05, -0.000154420441174397, 
    0.000480372691195914, -0.000347584071176242, -3.10923049717836e-05, 
    -0.000146164169051164, -0.000561736973477922, 0.000463444676331912, 
    -0.000984309782098559, -0.000134565496748699, -0.000354235690601011, 
    -6.24647275962237e-05, 0.00150356935234561, -0.000362530989056045, 
    5.44173489790496e-05, -0.000298824927992069, -0.00108933213611822, 
    -0.000214921800837672, -0.000585324349462594, 5.66833826031647e-05, 
    -0.000325649563798869, 6.79020123158926e-05, -3.71029170369277e-05, 
    -8.51712306706713e-05, -9.95873732541124e-05, 0.00157002775693827, 
    -0.000498233516021206, 2.86880605433072e-05, -0.000356479831632572, 
    -0.000866250592131899, -7.36610480992363e-05, -0.00108332949047761, 
    -1.78744186523136e-05, -0.000239920780246683, -4.45265118728346e-05, 
    0.00135689015856596, -0.000225062025006474, 6.95156776442026e-05, 
    -0.000244395347448267, -0.000444192525630826, -0.000266294947557254, 
    -0.000569581029953838, 2.50564663022267e-05, -0.000134710010425299, 
    -0.00053705171044229, -0.000808501029881113, -0.000188314258618663, 
    -3.28150649837462e-05, -3.83378642412669e-05, 0.00215569145836544, 
    -0.000454805054369884, 0.00013338809102392, -0.000440198893552002, 
    -0.00137461505405756, -0.000468239165608041, -0.00126969527369829, 
    -5.2481827435823e-05, -0.000272187993809919, 0.000173336052243076, 
    0.000818124066112343, -7.05427775574879e-05, 8.17784000040073e-05, 
    -0.00016381810790958, 0.000604003277230219, -0.00017147285830181, 
    -0.00060607749209495, 0.000109624015405381, -0.000445383177044416, 
    -0.000768513295597175, -0.00116070872468602, -0.000221870103130855, 
    -3.63051391717996e-05, 5.4426441703967e-05, 0.00192429473779745, 
    -0.000308624971445132, 0.000163049750442883, -0.00023832217727297, 
    -0.00126150272833224, -0.000444367604826582, -0.00151011399380711, 
    -4.45294853129563e-06, -0.000288152352340464, -0.000346682139727519, 
    0.0003934384172858, -8.99094118206121e-05, -8.03151641638518e-05, 
    8.1019577105254e-05, -4.40268014612376e-05, 0.00131641409942944, 
    -0.000133170879080035, -0.0005278298207929, 0.000209608916773471, 
    -0.000457595219322344, -0.00123307705442262, -0.00160736655058182, 
    -0.000234313088712183, 4.98186225329623e-06, 0.000222856099538719, 
    0.00125640271776902, -0.000135486919710306, 0.000155349379452675, 
    -5.75979397466167e-05, -0.00042832768006673, -0.000247220094671012, 
    -0.00117776660583705, 0.000128285913639215, -0.000374000888609369, 
    -0.00037693549025975, 0.000539651984414651, -0.000937902158603213, 
    -0.00014215327990069, 1.72960731550337e-05, 0.000143591546111122, 
    0.000868740445045861, -0.000249042280000286, -0.000364644943621258, 
    0.000291145809554553, -0.000127452864037425, -0.00114833835649335, 
    -0.00207477016250947, -3.39792697206131e-05, -0.000273015987074491, 
    5.91106441789002e-05, 0.000435471947305178, 0.000216717424356333, 
    4.75727588976917e-06, 0.000108282094843684, 3.12539028142802e-05, 
    0.000182655984249267, -0.00017026767610786, -0.000779558348053359, 
    0.000247012132058631, -0.000239939765218492, -0.000651692764153429, 
    0.0002977346656854, -0.00180486444429593, -0.00010858768666112, 
    5.82454824143845e-06, 0.000286256477482576, 0.000163942012777616, 
    -0.000330366612129384, -0.000217752042901257, 0.000286581034504439, 
    4.23994446488879e-05, -0.000493921256684938, -0.00172935160202081, 
    0.000101337764488274, -0.000202180843697343, 4.84880358011106e-05, 
    0.000673778920429562, -0.000921985277124473, 8.24964988430425e-06, 
    5.96916771427414e-06, 8.97948070711703e-05, 2.15607946725424e-05, 
    -0.000293099294106168, -0.00049891710550073, 0.000337789600091754, 
    -5.77456693237571e-05, -0.000464512856392673, 0.000171984037741014, 
    -0.00225708407093873, 1.22401370496265e-05, -2.46692397206255e-06, 
    0.000117058671965677, 0.000387868502092219, -0.000355660998268587, 
    -0.000291219660134909, -0.000132003106349912, 0.000228812676956656, 
    2.65552815621496e-05, -2.18268251851994e-05, -0.000985675990767355, 
    0.000215073816042631, -5.46139610045562e-05, 0.000113882257486916, 
    0.000671272763795281, -0.00177960475466506, 8.17335290016828e-06, 
    -4.41820741687307e-05, 5.3522409873305e-05, -0.000433778740825423, 
    -0.000323110635259144, -0.000358828139498152, 0.000371179797215648, 
    0.000183212953641065, 4.78678470328123e-05, 0.00016719843291083, 
    -0.00185794249640949, 6.19470912778628e-05, 6.55959433819677e-05, 
    0.000113127467346485, 0.000525420259772112, -0.000745421484930837, 
    -0.00022649344799385, -0.000109912536636657, 0.000149137963137159, 
    1.69246165222012e-05, 0.000115736650285577, -0.000496255623437239, 
    0.000303849859383049, -3.67621605092095e-05, 0.000177306599518806, 
    0.000469791585054018, -0.0017591953032047, 0.000332073639714685, 
    9.39125961552845e-05, 0.000110109163979514, 8.10673757110394e-06, 
    -0.000569191038907915, -6.98350508898162e-05, -0.000362576022141606, 
    0.000359130691823574, 0.000288341843782514, 0.000206135371972331, 
    9.69181431083235e-05, -0.000941287514015588, 0.00016347365165255, 
    7.2071454928678e-05, 9.667733002932e-05, 0.00041525299293963, 
    -0.000766328318493657, -0.00023247341444877, -0.000152466915708285, 
    9.93448870881008e-05, -9.30982388509259e-05, 0.000188920696908084, 
    -0.000297629041779439, 0.00040248484536409, 0.000202898029935282, 
    0.000306787889052984, 0.000328066824998229, -0.00135856880087984, 
    0.000260974424327929, 0.000166743185464835, 0.000124966287609181, 
    1.7550266062621e-07, -0.000481899757019475, 6.28891146200586e-05, 
    -0.000394512089884264, 0.000369418192359151, 0.000342603354269415, 
    0.000292674825129419, -7.39090876796681e-05, -0.000350256873394908, 
    0.0003112246401162, 1.44033304604742e-05, 0.000115143799039576, 
    9.01345461804437e-05, -0.000494577935771649, 0.000524710970793227, 
    -9.56241476160125e-05, -8.54547663717062e-05, 0.000174869104813476, 
    -0.00030722769905867, 3.7003254053492e-05, -0.000261997263324716, 
    0.000451280084424532, 0.000484255638085862, 0.000154947282222592, 
    0.000139885237836458, -0.000653788399731912, 0.000266666046108737, 
    5.73598691595882e-05, 4.92089030431012e-05, -0.000190312603469618, 
    -0.000471632305532191, -0.000113157566047482, -0.000413321159460174, 
    0.000425234098505356, 0.000150777041295738, 0.000486437599352336, 
    0.000165137321493376, -0.000128848447238142, 0.000442596739918202, 
    0.000153188399976692, 0.000147706721199219, 8.32255702638799e-06, 
    -0.000452606406310536, 0.000381179665584231, -9.15659780758695e-05, 
    6.36881081571877e-05, 0.00020054825170533, -0.000465163827088107, 
    -3.186521586834e-05, -0.000293606584530397, 0.000478409687260251, 
    0.00074096038287104, 0.000165815443616457, -0.00018611737755225, 
    -0.000174381678977293, 0.00036556683729694, -1.84073091213403e-05, 
    5.26358463759431e-05, -0.000263320938163548, -0.000384603598597906, 
    0.000525045058802383, -0.000197103060441771, -0.000418820850547809, 
    0.000502809702940223, -0.00034497041322589, 0.00041021580208238, 
    0.000406650061275136, -8.92774474392952e-05, 0.000523947907828451, 
    0.000512934994298476, 1.32745428648902e-05, 1.59861961667409e-05, 
    -0.000106174814667987, 0.000259298420139797, -0.000211212931278834, 
    -3.5382144141157e-05, 0.000167563927273786, -0.000589548192771605, 
    -0.000220668655235634, -0.000291193363047509, 0.000557276459213137, 
    0.000617611529118825, 0.000320249721353779, -1.98162840059439e-05, 
    2.92096406146529e-05, 0.00043018771752252, 0.000223116161304309, 
    2.59692532491187e-05, -8.66028118076579e-05, -0.000411414707425478, 
    0.000379571106495716, -0.000190321627325302, -0.000320565603823427, 
    0.000548706202213214, -0.000920763652423947, 0.000317023150751006, 
    0.000410963624633006, -8.11563906158144e-05, 0.000584315894037459, 
    0.00101051047663651, 2.33529112204919e-05, -5.16245937586004e-05, 
    5.19469778952724e-06, 0.000294593181358881, -2.60496564749274e-05, 
    -8.5327375135555e-05, 0.000161636661639801, -0.000586559859534313, 
    -0.000253145402951266, 0.000567101097292463, -0.000356179680101326, 
    0.000731138582208563, -0.000101814860114667, 0.000484685581021662, 
    0.000436575833873176, 8.99364659391334e-05, 0.000495072905122386, 
    0.000541766993639994, -1.491714123604e-05, -2.19678161226893e-05, 
    -0.000161964744312025, 0.000225264176653338, -0.000239836202308008, 
    -0.000383177707114384, 0.000496981642269179, -0.00124878745988538, 
    1.28194860406161e-05, 0.00050991849037981, -3.77466740903259e-05, 
    0.000695094869731354, 0.00103136798403005, 0.000168923321054791, 
    5.56437160112923e-05, 1.35050056794233e-05, 0.000293514133480324, 
    0.000151863781367794, 0.000160378019409594, -0.000420535327116901, 
    -0.000254974683431784, 0.000434508075371815, -0.00041627726722552, 
    0.00085587202467409, -0.00077561767033732, 0.000533126920068828, 
    0.000664129181010175, 9.63194629093137e-05, 0.000627365968591507, 
    0.00102347237288297, -1.01909617030042e-05, -4.32269259966541e-05, 
    1.24027834204624e-05, 0.000202506607575757, 4.77321571642139e-05, 
    -0.000403829113999351, 0.00048697782194207, -0.00119586505182141, 
    -5.44786214656757e-05, 0.000715754911952176, 0.000485340176430383, 
    -0.000210331443500792, 0.000891262843367476, 0.000313126898732738, 
    0.000412779644103673, 0.000485860269947445, 0.000197320672035503, 
    0.000341693205886328, 0.000505625138339241, 7.9822237099401e-05, 
    -0.000410466508032527, -8.00703429799363e-05, 0.000310591198682318, 
    -0.000613201511340803, 0.000767805014682038, -0.00114208839504109, 
    0.000388844596007189, 0.000831419466027265, 0.000128757345039508, 
    0.00075720777440131, 0.000986127230681646, 0.00021088780459018, 
    6.74997520980963e-05, 0.000131640962564634, 0.000174365961502334, 
    -9.48173068760582e-05, 0.000457014899314255, -0.000971187502072678, 
    -3.23383665996286e-05, 0.000560630149602416, 0.000249662311634101, 
    -0.000375778147926996, 0.000955530459159738, -0.000401940317558521, 
    0.000619234744222963, 0.00100273625613185, 0.000296259276572943, 
    0.000512241144014304, 0.000815915556303058, 0.000158336994157265, 
    -0.000216648695357669, 0.000113925737930567, 0.000211962073287939, 
    -0.000549496003168637, 0.000615430662356647, -0.000896247757149848, 
    0.000277487513683863, 0.000922225330951612, 0.000669400343820527, 
    -8.45437231109275e-05, 0.000877092502598944, 0.000476308311863991, 
    0.000451397731437031, 0.000462783681270422, 0.000334563520369132, 
    0.000189860469198274, 0.000345971823893342, 0.000380555406771389, 
    -0.000748163637832354, 1.60671701662347e-05, 0.000493808315452535, 
    0.000226680871002787, -0.000526824883489361, 0.000769410087097099, 
    -0.000658602616963788, 0.000605025633842588, 0.000993822050138135, 
    0.000214841824203311, 0.000636690949880008, 0.000800374748528832, 
    0.000324436336402931, -0.000149735698134867, 0.000275240233651088, 
    0.000148347710431608, -0.000354548550191167, 0.000401012136098728, 
    -0.00070285163813684, 0.000272431926351771, 0.000783832151973126, 
    0.000185189861993427, -0.000227952482563812, 0.000904396098792529, 
    -0.000229351411950988, 0.00067708504901354, 0.00086115486624956, 
    0.000336998310445578, 0.000307276799959399, 0.000644798466586771, 
    0.000409481123066414, -0.000608462253423135, 0.000151512323717312, 
    0.000291946675206413, -0.000680373797998691, 0.000432194914892467, 
    -0.000563870466922583, 0.000490033769237356, 0.000991513698792009, 
    0.000729175968549767, 3.07775411179955e-05, 0.000810152538931422, 
    0.000399129534336385, 0.000506538813965475, 0.000218333697568049, 
    0.000478257403086397, 0.000118710326238173, 0.000284802510382128, 
    0.000329992227975802, -0.000437666012897042, 0.000233280687249201, 
    0.000592202545680895, -0.000332614018034438, 0.000720217659819692, 
    -0.00045385828592639, 0.000690381505354311, 0.000229807711064725, 
    0.00043976735219915, 0.000571377143765124, 0.000376307448439786, 
    -0.000481899105039348, 0.000296695184195618, 0.000222870776894716, 
    -0.000637597587927344, 0.000109299286662628, -0.000224275152365604, 
    0.000424418603375799, 0.000948763268797809, 0.000104019979762366, 
    -0.000310682998252799, 0.000841752841766286, -0.000170109013236982, 
    0.000648845279561803, 0.000668674922082216, 0.00052395561155556, 
    0.000134489870292596, 0.000664231826001969, 0.000324818887677245, 
    0.0003544780834723, 0.00035973031202665, -0.000678480664987319, 
    0.000309832726504321, 0.000553057166716574, 0.000997576111871999, 
    3.80474394973293e-05, 0.00060857947760821, 0.000368053928798115, 
    0.00046380220856007, 3.1136640310547e-05, 0.000587073956906775, 
    0.000168372149752757, -0.000130898526011307, -1.4092003394113e-05, 
    -6.68682546024837e-05, 0.00037234702273614, 0.000606624380624622, 
    -0.000395639578027796, 0.000761357225606485, -0.000232971010057795, 
    0.000662598344619289, 0.00045519148919061, 0.000165347802155942, 
    0.000656250841509793, 0.000250203142998751, 0.000372929117201213, 
    0.000234041772967851, -0.000661802819427147, -8.6345442805272e-05, 
    0.000449688729590134, 0.000868431827428596, -0.000339384426021132, 
    0.000700462728503566, 0.000158936787519171, 0.000600701071581606, 
    0.00067195113816214, 0.000819748963581568, 0.00016747060221365, 
    0.000422451426718597, -3.82478690827045e-05, 0.000450934238184408, 
    0.000430427897038566, -0.000316956605960207, 0.000415660427549382, 
    0.000547969374070976, 0.000947827935417791, 0.000403989685547108, 
    0.000256027809749765, 0.000550160913472869, 0.000436557796505563, 
    0.000757475016927632, 0.000188674841739157, -0.000336698096312157, 
    -0.00035734790327982, 0.000432774645221182, 0.000572111860667055, 
    -0.000473947392795736, 0.000658476667789606, 0.000568906934205776, 
    0.000999205869663289, 0.000124599625864034, 0.000705440971430966, 
    3.79115670785814e-06, 0.000507773110124996, 0.000320294231914454, 
    -0.000133323145228873, 3.66676874106025e-05, 0.000320714707520928, 
    0.000866889079951729, 0.000264179304392677, 0.000375140453410763, 
    0.000745248065521917, 0.00121320730833576, 0.000105353129067701, 
    0.000281022954799044, -0.000475416946778396, 0.000426281363163919, 
    0.000469553154939583, -0.00021154407598714, 0.00036976565283125, 
    0.000425817589748755, 0.000801039236671804, 0.00103223998144521, 
    0.000104385334082489, 0.000352224693158267, 0.00099145206168598, 
    0.000231248772127336, -0.000226805881594962, -0.000277515154436438, 
    0.000290119908287384, 0.000657956962959916, -0.00017979497788744, 
    0.00026606681898852, 0.000634936924291807, 0.00179790196194219, 
    -6.81831085146225e-05, -0.000519098533530934, 0.000588469800374401, 
    0.000425125726574287, 0.000207545819873733, -5.64938733270408e-06, 
    0.000389657704056931, 0.000835570607823208, 0.00100386915109327, 
    0.000101254101099269, 0.000767519755622442, 0.00132274322387325, 
    5.1250748592039e-06, 0.000279937853973497, -0.000433294643049992, 
    0.000414204935430101, 0.000579409073487074, -0.000187950890333785, 
    7.51968565379323e-05, 0.000521024247679032, 0.000713631808574345, 
    0.00189281211265548, -0.000181583775453982, -0.000143764475934374, 
    0.000864022984850608, 0.000330460920427563, 3.1005216070631e-05, 
    -0.000314225408195631, 0.000490006105758443, 0.000820803522925132, 
    0.000475313595909279, -3.49038410409918e-05, 0.000788689956546346, 
    0.00188625945282606, -0.000367626253955864, -0.000486755005189833, 
    0.000485308809248405, 0.000495152774793922, 0.000451002152626994, 
    -4.59090080728202e-06, 0.000659575251552943, 0.00079945707231265, 
    0.00139860252986914, -0.000192251718201107, 0.000358385739280945, 
    0.000969783048569111, 4.19655920186424e-05, -0.00040364536423642, 
    0.00060889841519203, 0.000738266808793972, 3.50642152247526e-05, 
    -7.59644395502111e-05, 0.000715639310044346, 0.000825720341030508, 
    0.00174341914125784, -0.000704264559713556, -0.000307073906407906, 
    0.000308403712040206, 0.000422120046704533, -3.07879814021489e-05, 
    0.000882268479727728, 0.00082423040973135, 0.00082207819279295, 
    -0.000192105120661823, 0.000466629350745031, 0.00133276511009857, 
    -0.000320781675440797, -0.000392026505478004, 0.000478532479362843, 
    0.000627531965515894, 0.000550629222224818, 7.83305110296878e-05, 
    0.000880058981303862, 0.00089054288578523, 0.00112049671784039, 
    -0.000787203188549439, 0.000108137541030408, 0.000336163841107104, 
    0.000190173681190827, -3.28522936013081e-05, 0.000867314243467372, 
    0.000728654148216603, -0.000106380580877712, 0.000337191684269504, 
    0.00103297045798926, 0.00119476648691583, -0.000779852571292062, 
    -0.000267884052074845, -7.80643480250673e-05, 0.000554031100005617, 
    0.000332208188097095, 0.00106896181169821, 0.00082050553545685, 
    -0.000603724588522555, 0.000279778130395881, 0.000471090107783396, 
    -0.000176391088498896, -2.85212170769372e-05, 0.000660636560815626, 
    0.000664381717250215, 0.000214141385010182, 0.000504677405734098, 
    0.00100677967472774, 0.000627068130389577, -0.000920945045513656, 
    5.91552905437785e-06, -0.000173332918974694, 0.00037573106945838, 
    0.000394724577424982, 0.00106307031376098, 0.000734308161917717, 
    -0.000369084989834235, 0.00030530360728848, 0.00108740027508226, 
    0.000951699574126154, -0.000766709946541347, 5.67579699601226e-05, 
    0.00020830611240543, 0.000612406137308364, 0.000688564511441431, 
    0.000977129720777524, 0.000885909097233584, -0.000774999411170951, 
    0.000203064870165996, 0.00011676481987104, -4.07633355366311e-06, 
    0.000394418644097383, 0.000914484237975371, 0.000774119905274635, 
    7.46310816404898e-06, 0.000493534824952378, 0.00108273707031498, 
    -0.0010964160017603, 0.000126050451936222, 8.6413613962619e-05, 
    0.000462114239525444, 0.000770487627783357, 0.00122837843045908, 
    0.000809813118391566, -0.000543370109198942, 0.0001555435051414, 
    0.000760516353233758, 0.000808114243157075, -0.000560357814463395, 
    0.000460182915802093, 0.000564956717690983, 0.000754132948256577, 
    0.000602237194741102, 0.000813155720521957, 0.0010218884573159, 
    -0.00101399292792959, 0.000241936807959558, 0.000257204538692098, 
    9.6238869026757e-05, 0.000612217653715227, 0.00136332582851025, 
    0.000832404700378217, -0.000202990689594632, 0.000168788927604472, 
    0.000905187774266996, -0.00127290346492251, 0.000404924874786948, 
    0.000343970782532722, 0.000608794407292069, 0.000717920490272293, 
    0.000843272948796726, 0.00100132772676268, -0.000753204090219677, 
    9.89910649271063e-05, 0.000509199052376577, 0.000749349794620182, 
    -0.000310917146385012, 0.000607325720223239, 0.00119798670840821, 
    0.000792222444387257, 0.000284073463620404, 0.000321923860408552, 
    0.00103444494057953, -0.00160844775317193, 0.000407230867005947, 
    0.00044327268521191, 0.000376350538035822, 0.000316720739164743, 
    0.00130015919557916, 0.000973644329619413, -0.000556967073839389, 
    -0.000154478058392568, 0.000587089263345079, -0.000998353581938877, 
    0.000552042274227568, 0.000792740299886634, 0.000712931165481764, 
    0.000380445905305635, 0.000352809035492157, 0.00120648337150994, 
    -0.00154706747238663, 0.000213477717565164, -0.000166115993361399, 
    2.29607024743779e-05, 0.000389573952043189, 0.00126353630161963, 
    0.000890588270448529, -0.000214972367001779, -0.000360821454250552, 
    0.000750262436203849, -0.00155152355911797, 0.000481214483991127, 
    0.000531713483331668, 7.95580046480214e-05, 0.000808849999135469, 
    0.00118484982159679, -0.0014556563079386, -7.53570276268595e-05, 
    -0.00024698087734549, -0.000539479092057752, 0.000572670288977311, 
    0.000950070329598141, 0.000817452133970747, -8.55439621298163e-05, 
    -0.00039278616478823, 0.0010925346865292, -0.00156515846902258, 
    0.000258395490534014, -0.000558981741647916, 0.000133859439686975, 
    0.000205739724739955, 0.00109623857103657, 0.00107077285236282, 
    -0.00146096532650535, -0.000336387778574644, 3.49508900596936e-05, 
    -0.00109814168329521, 0.000442866003810815, 0.000637024404011761, 
    0.000597421819946146, -8.196860662649e-05, 0.000126980113800908, 
    0.00114213532561499, -0.0014308658827726, -5.64085410881432e-05, 
    -0.000758433817123074, -0.000397923852144999, 0.000373857973969454, 
    0.00087963105364039, 0.000894634477896156, -0.00116839100285336, 
    -0.000483965329128305, 0.000463675224452042, -0.00106317136831487, 
    0.000209435417774162, -0.00110317197981156, 0.000220234455024556, 
    3.16254708088456e-05, 0.000583794334725702, 0.00104294562814035, 
    -0.00127847357124489, -0.000252634745066303, -0.000380252749390417, 
    -0.000831729614261661, 0.000322038344020384, 0.000690135895248047, 
    0.000545179443857957, -0.000621258877312076, -7.82298422029343e-05, 
    0.000625569144168581, -0.000803739460204207, -3.44851597096979e-05, 
    -0.00155809090945333, -0.000214018654200703, 0.000141943076469502, 
    0.00084408125762125, -0.00109948354277132, -0.000352731256419884, 
    8.46133900781568e-05, -0.000796988872389617, 0.000112924622884212, 
    -0.00152279129661011, 0.000143387794686461, -0.000272963537153954, 
    0.000219842134616977, 0.000609117534374993, -0.000671896912523466, 
    -0.000284309485008946, -0.00136515701741474, -0.000504234542814616, 
    0.000179143029532114, 0.000501849622080289, -0.000746634137041746, 
    3.50179452155294e-05, 0.00027428093730609, -0.000638852411576019, 
    -1.18721121325839e-05, -0.00198174369230991, -0.000209623137869162, 
    -0.000102215352853606, 0.000619775954541878, -0.000610883553686369, 
    -0.000262678000033137, -0.000691575988881665, -0.000504659108978852, 
    7.0900758038213e-05, -0.00146366255768247, 0.000122707132089361, 
    -0.000440594162943518, 0.000201013809502531, 0.000243399037830673, 
    -0.000553158355985138, -0.000286512088164619, -0.00191801930219947, 
    -0.000356348283563665, -0.000205526751160056, 0.000607005449003656, 
    -0.000516680284349989, 4.98256845919699e-05, -0.000285670494304532, 
    -0.000447587372484714, -2.77989807515364e-05, -0.00173351947839555, 
    -0.000168218138757868, -0.000227866899141455, 0.000351671424007748, 
    -0.000514334939208724, -0.000373818689087034, -0.00137824618832343, 
    -0.000426729806629234, -0.000423759733720887, 0.00067527727212142, 
    -0.000464558603521923, 7.43606034670739e-05, -0.000214557603138183, 
    -0.000402720184906867, -0.000134726229988354, -0.0016042233302564, 
    -0.000328123902647743, -0.000254117316920039, 0.00061670873655196, 
    -0.000383950018102533, -0.000179293902281273, -0.00111362701681178, 
    -0.000269605134532252, -0.000372867480586624, 0.000820870731871579, 
    -0.000290918627985741, 0.000108495005779575, -4.47920775256881e-06, 
    -0.000426912451272401, -0.000202272920052403, -0.00142858555846981, 
    -0.000482278517749058, -0.000367236855763464, 0.000988783071820933, 
    -0.000245963775894343, -8.83200882032129e-05, -0.00097748998944387, 
    -3.13177741371431e-05, -0.000149357612293618, 0.000903918819573101, 
    -9.17525395567056e-05, 0.000447711093863692, -0.000220460851342548, 
    -0.000197566220239617, -0.00152343200314197, -0.000321181931254258, 
    -0.000302317971914949, 0.00138630977734056, -0.000133910318121017, 
    -3.12370647461976e-05, -0.000795000828526925, -3.15523761243749e-06, 
    1.67930340700717e-05, 0.000730889149301955, 0.00028762026177106, 
    0.00100002462201806, 4.83810396536115e-06, -0.000177067851353885, 
    -0.00140292918657145, 6.66443537558848e-06, -8.02759163168039e-05, 
    0.00172348880434986, 7.33810312304855e-05, -0.000383711871307906, 
    0.000118733521705932, -0.000120012910536414, 0.000690495343788667, 
    0.000484526825243228, 0.00164948166999489, 5.69192800046196e-05, 
    -0.000173535606325178, -0.0011670619629913, 6.68367329955133e-05, 
    3.46516533947053e-05, 0.00171416945464568, 0.000528052981721358, 
    0.000292708588005104, 0.000257395315960856, -0.000156270546507706, 
    0.000653027592887098, 0.000498665861316174, 0.00215323049982671, 
    0.000305975783014051, -0.000811705288812312, 0.000109805546014849, 
    -1.49506456581898e-05, 0.00155780686064061, 0.000810272881957489, 
    0.0012897348994697, 0.000325094733011545, -0.000329277745358122, 
    0.000317363115162186, 0.00045211633450616, 0.0022255387424685, 
    0.000700329190694571, -0.000143958552171685, 0.000220226400008278, 
    -6.85886042089564e-05, 0.00106382581248092, 0.000723860728311718, 
    0.00183056254481515, 0.000631037302399196, 0.000381383615208068, 
    0.000381537905649647, 0.00199478271704094, 0.000910765347764576, 
    0.000738173772015117, 0.000384306421963909, -0.00027509816409395, 
    0.000556334536366454, 0.000598745117400459, 0.00164760231976311, 
    0.000754918502723607, 0.000378755178525241, 0.000235725933037909, 
    0.00114347809674383, 0.000717601451788277, 0.00131789812957766, 
    0.000652579837504388, -0.000576251215493904, 0.000638102470185832, 
    0.000459527628035085, 0.00120878679690933, 0.000535581467755201, 
    0.000344770462138419, -4.36869259723065e-06, 0.000754827400880894, 
    0.000555907057755358, 0.00130371257571316, 0.00058476126733842, 
    0.000707172512172298, 0.000229284868288534, 0.000586207482518843, 
    0.000337674077060821, 0.000293668546726336, -0.000417619367064559, 
    0.000743541510619722, 0.000237988329765711, 0.000896583231750133, 
    0.000408818147115909, 0.0006416993499168, -1.30985432326921e-05, 
    0.000572387070967309, 7.20223675550957e-05, 0.000566560023667758, 
    0.000731147914228454, 1.8801548782804e-05, 0.000425004391884382, 
    0.000142142807741815, 0.000462179569236139, -0.000414133508093071, 
    0.000846309436745716, -0.000256576512818179, 0.000779366629565725, 
    0.0008376482225959, -0.00015416346439057, 0.000563039173493593, 
    -0.000196553949314749, 0.000771702038654868, 0.000951408174568289, 
    -0.000569477480700698, 0.000303272010021256, 0.00102477990259141, 
    -0.000331636073747797, 0.000904646757645306, -0.00050844963880941, 
    0.000990771670366211, 0.000868675690995447, -0.000532404482625936, 
    -0.000207162602218374, 0.00119661884468002, 0.00123524807956241, 
    -0.000751566338415767, 0.000616025314417345, 0.00111098486692505, 
    -0.000286003695085192, -0.000486444939595841, 0.00121447868622336, 
    0.00127899872899638, -0.00068694275047238, 8.14625518504536e-05, 
    0.00130517876949769, -0.00064615885992459, 0.00104038791659462, 
    0.00130232929081861, -0.000369256520093211, -0.00034052347300459, 
    0.00117115421506578, -0.000667587256171943, 0.000663543461595764, 
    0.00110039568350064, -0.000128247040602001, -0.000512277958952002, 
    0.00105877381663641, -0.000449210037429665, 9.4211473612781e-05, 
    0.00105271358922041, -0.000563429202068344, 0.000858600628559444, 
    -0.000163721683177979, -0.000277321332512263, 0.00100756390137125, 
    -0.000390028812517206, 0.000365014040720687, -0.000354552943210192, 
    0.000689945655946852, -0.00014419843804133, -7.8920493255974e-05, 
    -0.00028025742708076, 0.000356043965488915, -0.000288362327198186, 
    4.79600733294588e-06, -0.000287828750908936, -0.000162419435008889, 
    -0.000283659606977782, -0.000162476264228329 ;

 misfit_initial = -0.287175043125849, -0.500655712857547, -1.188292728781, 
    -1.22008858893034, 0.739995810529539, 0.433400478731816, 
    0.390879661504826, -0.353370903367507, -0.635422137192201, 
    0.155947216855763, 0.217177610644761, 0.0350171434937074, 
    0.222721001072523, 0.0506249018675353, -1.90844817248254, 
    0.0496995292673086, 0.653020639715192, 0.685881324494386, 
    1.42749212047843, -0.124884845580522, 0.0993573971156847, 
    0.217515931173971, -0.173302343270345, -0.843914067799965, 
    -0.203618141994775, 0.161433263824922, 0.10719481286924, 
    1.30779828688122, 0.484078997626729, -0.832224465541, 1.76101618868901, 
    2.89002291992905, 2.0027008185647, 0.2245891574134, 0.378251133511478, 
    0.774460334742391, 0.455675487737177, 0.486266124769172, 
    0.834887247276326, -0.309940963178668, -0.93803481291717, 
    -0.511314222684351, -1.57469188771736, -1.00168860730933, 
    -0.657259944288211, -0.54030927820452, -0.893068233974668, 
    -0.0238211519044729, -0.335669852092093, 0.0782615547374776, 
    -0.407011554073295, -0.437170860617417, -0.161171941408433, 
    -0.469235660666252, -0.327937220716423, 0.33469449788722, 
    0.690608335214309, 0.637106679852346, -0.380756200817629, 
    -0.586264853088156, 0.336332353516218, 0.243495475157376, 
    0.0251642878520553, -0.191613548169585, -0.0958624385270568, 
    -1.40920834558038, -0.52380612202223, 0.2687467794301, 0.499674311657201, 
    0.673850617925651, -0.260613888896839, -0.183106472036889, 
    -0.0475011099961842, -0.763348516938573, -1.4660895066171, 
    -0.423784316914895, 0.0173582951352769, 0.422808895890441, 
    0.56503008534794, -0.112617051387196, 0.463578763795289, 
    0.526341185759858, 1.11282690137725, -0.0225096716108553, 
    -0.761279093125364, -0.0427533286720072, -0.0314140557845688, 
    0.251826053285145, 0.0203620054231912, 0.264380226751388, 
    -0.321061041627635, -0.659319354851231, -0.86910352655138, 
    -1.40826249564828, -1.36613100767985, -0.778149032018924, 
    -0.755357819653848, -0.106271304950427, -0.363663523927089, 
    0.319631134253306, -0.352769459598981, -0.755758130911923, 
    -0.231368377472334, -0.0331786561632974, 0.0938662579033434, 
    -0.660970181296312, -0.518645232812274, 0.478772378785521, 
    0.521989214794409, -0.634379800905798, -0.737720613497146, 
    0.265668183843148, -0.0470014129876439, 0.1854243999784, 
    -0.718135730252722, -0.880466538564284, -0.857034387340643, 
    -0.0716956117374234, 0.355403189672074, 0.312609559170993, 
    -0.993300765413876, -0.425030916460227, -1.23782342132705, 
    -1.25020493110464, -0.8335585657764, -0.981737436752113, 
    -0.0482822317033804, 0.392395924540598, 0.405041711282061, 
    0.46159808971722, -0.339420302778914, -0.5242259992256, 
    -0.113693175404732, 0.240814046695599, -0.479576796811387, 
    -0.708871172588421, -0.0148944135829954, -0.316118075791305, 
    -0.204966442171046, -0.0524375221205586, 0.163779559956536, 
    -1.67599646287627, -1.89382595224206, -1.28126755003725, 
    -1.24063103722185, -2.26318486977712, -1.55173834676967, 
    -0.15614699951966, -0.034887492562401, 0.5293587908923, 
    0.0514598363321417, -0.866302733472994, -1.43459520364004, 
    -0.780676404077614, -0.435633777433004, -0.575247601002218, 
    -1.09794636104106, -0.685349121134351, -0.141223802051496, 
    0.293536524717313, -0.196323773157507, -0.3770157829869, 
    0.0494576216403786, -0.062620118537744, 0.0965007804584683, 
    -0.396784784219095, -0.582444498911232, -0.108242252259232, 
    -0.60807318676027, 0.371107192351356, -0.180204588562018, 
    0.081938782467682, 0.767689573870456, -0.359735292573746, 
    -0.765298240727668, -0.101499120032043, 0.404898157813074, 
    -0.0671404069346515, 0.951037172633922, 1.36416234625869, 
    0.789244756857368, 0.0783274791695021, 0.313328305816469, 
    0.802349144125123, 1.11088150109275, 0.175768924285897, 
    -0.874110091944691, 0.275339121146865, -0.608569711798319, 
    0.299394394222583, -0.110148340685021, -0.121425488731264, 
    -1.12217683217279, -2.25696797993985, -1.63041177279247, 
    -2.69352548522757, -2.7535189987913, -2.06458726171747, 
    -1.14300593038572, -0.111995928134108, -0.135775438790247, 
    -0.292974747482004, -1.51913317537007, -2.74699689055711, 
    -1.10478068998231, -0.724243969563956, -0.367949182440244, 
    0.00162763890656059, 0.348999707437683, -0.203874635163679, 
    0.676500001668652, -0.0365628948851704, -0.197517964040275, 
    -0.425725328111177, -0.277707151352216, 0.0523803576044735, 
    -0.00935928542085129, 0.0572390192928784, -0.0173439309249002, 
    -0.596454246522997, 0.0728920192768445, -0.58588476438326, 
    -0.847400244254941, 0.13802639983775, -0.0835058240146402, 
    -0.471600182691856, -0.23072737884497, 0.294022280794297, 
    0.914903343977622, 1.28228602149755, 1.61404191931057, 
    -0.731711193794209, -0.875827007346874, 0.306338212901207, 
    1.49358969099689, 1.78133440156332, 0.714617789240735, 0.386956314861089, 
    -0.376598009620168, -0.102545315022167, 1.08113117774403, 
    1.03696579882775, 0.800910753187547, -1.17044418056425, 
    -2.18189486939862, -1.82438099071697, -2.46132631456117, 
    -1.49722027265668, -0.712071635948903, -0.358033566023561, 
    0.132414632809557, -0.209240946993807, -0.0287540091742677, 
    -1.29719774565347, -2.66591244364048, -0.204230496752498, 
    -0.198541647099759, 0.305227391689664, 0.350296979771834, 
    0.660839089532272, -0.303068293723934, 0.108926627374331, 
    -0.247836039177241, -0.421123029392723, -0.771509026850845, 
    -0.386865191225221, 0.0240060867606751, 0.324627176851671, 
    0.731437328220461, 0.0606043288034686, -0.259597478391034, 
    -0.328310289266098, -0.34327153258908, -0.849169578391122, 
    0.404657995749758, -0.0152314417853994, 0.0238685601490696, 
    -0.0746754779047443, 0.139198167456018, 0.932271281341248, 
    1.57539174530632, 0.953565097997284, -0.968103868599508, 
    -0.805265045647094, -0.0386432286806793, 0.802805863613023, 
    0.401168277263162, 0.660526431517128, -0.492642339082288, 
    -0.938116270416285, -0.805114949625407, 0.0953364860619432, 
    0.753460355321551, 1.00266745485107, -0.849727594566985, 
    -1.3419796587278, -1.59129851863592, -0.735793290765634, 
    -0.691708709737875, -0.314183230662279, -0.0741332601546363, 
    -0.0583137587963778, -0.229235590926473, -0.577295793490769, 
    -0.676143071373896, -2.20260661300058, 0.38588040567233, 
    -0.381925381115487, -0.24247867451356, 0.434220236195131, 
    0.542181099882635, -0.506274375159723, -0.0536187146928402, 
    0.0147953063844408, -0.199586241030989, -0.380918242650505, 
    -0.121297405501037, -0.0587879306029215, 0.755207975016279, 
    0.562652631964258, -0.90751777417704, -1.96482494305777, 
    -0.355456294118542, -0.606855999793097, -0.485335550970341, 
    -0.449316703010485, -0.28289591491204, 0.263977578640757, 
    -0.299725334677849, 0.409575825096091, 0.908450809013535, 
    0.510648144404962, 0.502381289344531, -0.457388931206846, 
    0.341815609642087, -0.00550599781871774, 0.227000435056715, 
    -0.682323711964923, -0.0838770805689526, -0.569779143146021, 
    -0.646950310637542, -0.129947281412117, 0.154108604659302, 
    0.0855404735367626, 0.646434214528453, -0.585484465651116, 
    -0.889799528560822, -0.881322380297873, -0.337557513803475, 
    -1.09571470368422, -0.507996963078652, -0.47457792433828, 
    -0.554972940207135, -0.619447903340644, -0.759322326408052, 
    0.694307267919933, -0.00715723222446601, -0.238928894693391, 
    -0.0590245535098255, -0.135681961879204, 0.842325087336988, 
    0.198599776116417, -0.107028794548878, -0.0296071398990705, 
    0.2560349256109, 0.403688955291757, -0.0254862016431501, 
    -0.492926061171537, -0.22384943441236, 0.232615292495901, 
    0.26188835106459, -0.252557995201452, -1.43628187158366, 
    -0.10748909395665, -0.300905094801291, -0.963670303152551, 
    -0.857184492991765, -0.279363655411333, 0.564724222745325, 
    0.561772818185933, 1.36627409072356, 0.630719615345794, 
    0.537764496615036, 0.410167567793356, 0.0263797049043735, 
    0.484856309479045, 0.697225619059076, 0.432440057772903, 
    0.174267514412918, -0.341561884205852, -0.602762814817179, 
    -0.311114150223704, 0.139557866771116, 0.0931065100953088, 
    0.410207686324622, 1.08724814004405, -0.290638083097479, 
    -0.856987961721987, -1.28557892706353, -1.14802395469253, 
    -0.629890837907778, -0.761551529749993, -0.347410422189225, 
    -0.506524690057804, -0.236982780423158, 0.511565554429137, 
    0.5430511607499, -0.988621511798491, -0.0820197546313928, 
    -0.360628739390485, -0.15355197982414, 0.161388946274643, 
    0.276551348970031, 0.138730036016064, 0.404464004742984, 
    0.505338211000739, 0.274749570986499, -0.803410240088929, 
    -1.16242185947224, 0.130764826997725, -0.353577449509963, 
    -0.295942149510253, 0.0512204999681831, 0.160456492611896, 
    0.280650436896717, 0.0639210707989113, -1.09584348825507, 
    -0.816880994789284, 0.193663681236074, 0.7919127659276, 
    0.982174612758091, 1.0314830233448, 0.468084048798065, 0.744531829137726, 
    0.461439319767694, 0.7417449256533, 0.413364644848957, 0.492449517117, 
    0.576475866791819, 0.604950281773555, 0.248316037188046, 
    -0.116288116866672, 0.280019177092274, -0.767655203587956, 
    0.0976963695523692, 0.544135936452577, 1.09967487047527, 
    0.44953621439368, -0.722874308486636, -1.86322441252529, 
    -1.16875866952894, -0.574191755854554, -0.701528687269373, 
    -0.24121175665301, -0.557769453814005, 0.489874371066401, 
    1.66609962504093, -0.215229402279464, -1.49114763869746, 
    -0.651222832273275, 0.176488719320824, 0.229674033276757, 
    0.760497714948682, 1.21766394617419, 1.19016909967966, 0.195004691120966, 
    -0.257121460488072, -0.637997443626173, -1.31944629594934, 
    -0.726140383632461, -1.16420056685254, -1.36580864493719, 
    -2.21918505977258, -1.69463939149899, -0.174657680035865, 
    -0.264726695565312, 0.373819514044924, -0.634916894986257, 
    -0.782346273627987, 0.200485217597111, 0.892215985881206, 
    1.14853625839855, 1.15075973739005, 0.203598816197839, 0.768815112262575, 
    0.589166530576306, 0.88028366551026, 0.706781710270867, 
    0.106567757121843, 0.516988036450305, 0.814603731923254, 
    0.332854327738961, 0.750675262472691, 0.769314756329234, 
    -0.138744664261794, 0.246192933314808, 0.67251827281726, 
    -0.517505645665897, -0.292987956944679, -1.51845331872226, 
    -0.86014988179921, -0.540446851891856, -0.835263038282537, 
    -0.00499560414706668, -0.0194188481618474, -0.549598612085931, 
    0.0825304767422841, 0.769679901790305, -1.62902428978168, 
    -1.54700618085116, -0.966353914260916, -0.238069273543893, 
    0.11960675374648, 0.467526128260438, 0.291155904332294, 1.18268350335287, 
    0.0956497443977256, 0.00412070086887262, -0.368922649385111, 
    -0.756279189853704, -0.280137962018703, -1.26243138624853, 
    -1.2577490295389, -1.47068677571438, -2.10521686479917, 
    -0.391913230481795, -0.97344760923407, 0.284072387813792, 
    0.352015614730377, 0.00244584026031447, 0.484255989810758, 
    0.309064147691207, 0.334205139004378, 0.220002715373631, 
    -0.154477165652054, 0.863869909071697, 0.567454364759641, 
    1.05517673424054, 1.47609922067445, 0.0619717868939862, 
    0.0542959490181305, -0.65735906143312, -0.623947821353914, 
    -0.385571952013648, -0.301359332653908, -0.604559028961527, 
    0.892187291972579, 0.987160512045051, -0.365584656098794, 
    -0.430138937580304, -0.577622620967801, -0.280862736587308, 
    -0.874360390067741, -0.869755730244517, -0.689624000165741, 
    -1.23044635173351, -0.238519936455246, -0.300872401040788, 
    -0.405173150565257, -1.85144232354925, -1.38826870219782, 
    -0.532466045981961, -0.163994060374408, 0.312415626961089, 
    0.166770311760445, 0.306387403136492, 0.202937720822156, 
    0.171596495778319, 0.146005166943493, -0.156704930942655, 
    -0.69584272498274, -0.295018918840926, -0.844271597676474, 
    -0.542807374943983, -0.0819556079764716, -0.400556901089577, 
    0.0197171950134978, -0.865571612879177, 0.530891964819311, 
    0.0379169705052762, 0.447281203607472, 0.364240539850837, 
    0.726725618272273, 0.671660618301249, 0.192480530744561, 
    -0.0799054890946094, 0.875431726226235, 0.773735136109823, 
    0.59345215169091, 0.35823284038945, -0.925048073428667, 
    0.240626691017702, -0.145323599360694, -1.13559748351694, 
    -1.50593608686706, -1.16066622512351, -0.330874859249, 0.533067934400355, 
    0.77564236614371, -0.224109349854844, -0.563202211921858, 
    -0.51128958656979, -0.355925686224263, -1.15699583381335, 
    -1.78568956070317, -1.15502730294208, -0.901023156299652, 
    -0.532929647241271, 0.238737223929138, -1.10469217083499, 
    -1.9127716195548, -1.45066278534617, -0.26778507905628, 
    -0.209556593129134, 0.212133446775846, 0.185768493144476, 
    0.368394113822141, 0.520100033282151, 0.251848521440996, 
    0.0686789577337432, -0.660607188618569, -0.498658339611504, 
    -0.464203865934461, -0.995760202588607, -0.236856553628177, 
    -0.365543700655033, -0.526485510853214, 0.306684437834228, 
    -0.300714255118648, 0.606860619654781, -1.17379971887849, 
    -1.08236435135289, -0.505925378748517, 0.297535385000356, 
    0.965782434423121, 0.282260166729533, -0.104625754528573, 
    -1.1671844214551, -1.06108315125132, -0.659607340231068, 
    -0.990302080966887, -1.91138718897067, 0.52083199096177, 
    1.24160367494726, 0.619068934837856, -0.0424798385884495, 
    0.149740039096611, 0.99341342176642, -0.222380648692981, 
    0.0594853092875569, -0.651345766116065, -1.16525434192253, 
    -0.686487390191277, -0.488055018794711, -1.05701680878545, 
    -0.863705137587711, -0.422121300670937, -1.10159310886915, 
    -0.692309107257572, 0.126766460318524, -1.34083100594471, 
    -1.44391798592138, -0.889273497931464, -0.191252010249237, 
    -0.58240368053232, -0.135613101334728, -0.354631029904988, 
    -0.149289639359056, -0.566208164389819, 0.501174441564523, 
    -0.503920390647066, -1.30466675108408, -0.771663311312145, 
    -0.59277962199233, -0.620550842346299, -0.338845437060344, 
    -0.384174305022227, -0.622992855950462, -0.0687689797292812, 
    -0.0702887128180185, 0.761132467473566, -1.78076054358834, 
    -2.13682198407128, -1.19164381887691, -0.00642062259054832, 
    1.47924514848138, 0.391767340131222, -0.462140876936421, 
    -1.68375151088974, -0.760321530211918, -0.0580445989550915, 
    -0.495905172277138, -0.622147499619135, 0.713129760949962, 
    1.43866946368918, 1.60860913636797, 1.27177317532685, 1.73756224404745, 
    0.821961899494945, 1.88277122170907, 1.43095358823623, 1.35895693031412, 
    0.286725891152604, 0.232735954661418, -0.0517290005119975, 
    -2.1038417061551, -0.848445641701017, -0.0790030874128611, 
    -0.0770833529584673, 1.04375866791346, 0.200730157120257, 
    -0.010561893134033, -0.361018494270788, -0.0583269195101188, 
    -0.469316126929806, -0.594141370550476, -0.902649123431756, 
    -0.876743089326499, -0.615906125933403, 0.482393549437719, 
    0.433982127458714, -0.25742890796697, -1.29894114015513, 
    -0.466761740291521, 0.299377728394021, -0.364313744140707, 
    -0.589934782325079, -0.544869929334491, -0.328138695908731, 
    -0.292711736092897, -0.528312773533917, 0.262804486570225, 
    -1.95185212095915, -1.90799958610111, -0.990015954860439, 
    -0.140918679083062, 1.27149865082353, 0.503955692901195, 
    -1.47037501185724, -1.95977935062587, -0.797853597362019, 
    0.0818570667587259, 0.41127496971411, 0.226002161134011, 
    0.505991410228801, 1.02618607832938, 1.1242051240611, 0.751020195228391, 
    1.08431141272843, 0.719628508175325, 0.985727682414943, 
    0.916633198933301, 1.39629981757893, 0.655884908019129, 
    0.581010826866688, 0.292296585877665, 1.11791832017013, 0.89060940525793, 
    0.650005595251448, 1.14064840063756, 0.177065432164545, 1.63648275538664, 
    0.159503153806422, -0.917885828150649, -0.784512456193776, 
    -1.13889385618833, -0.944107264561564, -1.03795977379569, 
    -0.81354218364714, -0.678976497159081, -0.265487585497564, 
    -1.00784051804516, 0.648506647570257, 1.07134923195823, 
    -0.0718876707055616, -0.479231748855162, -1.09277312339151, 
    -0.71223829929008, -0.972507323486624, -0.801094893487888, 
    -1.07869520024354, -1.76297683036285, -1.37311064566343, 
    -0.770105940523389, -1.10529016707697, -0.418066161290991, 
    0.303425028360995, -0.452141896916398, -2.02733159841605, 
    -0.698424273453675, 0.128381382988225, -0.521204477841932, 
    -0.597751949234859, -0.381570474191095, 1.51463822944528, 
    -0.243141500315933, -0.434794364004429, -0.432501928007261, 
    0.10015338878822, 0.822651598360165, 1.88850610790088, 
    -0.654705429832493, 0.732230231800188, 0.22916449846389, 
    1.65238165528909, 0.252703866039266, 1.12460474442399, 0.390670823280903, 
    1.08528199384651, 0.274818413832419, -0.570725874812783, 
    0.0574693567980049, 0.0525736355879403, 0.00939872292971031, 
    -1.45922748406614, -1.48063121766699, -1.26552643601888, 
    -1.38412294454471, -1.67604759595136, -0.595585103823302, 
    0.562584991232997, 0.0909025391580798, -0.73359442596626, 
    1.25270601319167, 2.01970272753492, 0.772695790058626, -1.0579210111224, 
    -1.50747316403637, -1.60727440210767, -1.80689773392758, 
    -1.07232693117175, -1.4166109646794, -1.33726968903946, 
    -0.427369291332109, 0.00089760184840415, -0.894039541348222, 
    -1.17117044568089, -0.59248876276738, -0.415899329960219, 
    -1.21177100444969, 0.137425629664283, 0.154021300633485, 
    -0.850592025570291, -0.899836672376866, -0.161913470323745, 
    -0.735970664352409, -0.415399494868092, -0.906006145827849, 
    -0.436058874180385, 1.59732368455522, 0.617135773037734, 
    0.682060982589503, 0.247144505015076, 0.733815510526821, 
    1.53811170508593, 1.56392539979723, 0.696502137671886, 0.576809470068911, 
    0.881167250070458, 0.210029452242392, -0.546550249619004, 
    -0.05469092774324, -1.23380215986248, -0.248972608325522, 
    -0.488639524014252, -0.682607878852561, -0.959602271581224, 
    -0.393364612331646, 0.4949989752064, 0.731165867736756, 
    -0.218373983605735, 0.833264410889014, 0.20013039046944, 
    0.0171183064019065, -1.30833603828677, -1.44987521771931, 
    -0.961289593507835, -0.935994710358141, -1.41801050730042, 
    -1.72243106813314, -0.844047715445906, -0.471384264824102, 
    0.00519223561240789, -0.173729447261284, -1.03134464256848, 
    -1.37784252376587, -0.909921791768764, -0.940398102012514, 
    -0.117964612784798, 0.13602703346673, -0.176414890051628, 
    0.35008155696313, -1.04937706270889, -0.7101033210233, 
    -0.193303503734459, 0.705463143799679, 1.80709356243802, 
    -0.344646733730559, 0.381370038025559, 1.09319674946498, 
    0.979607118150608, 1.20943913631747, 3.32024302323322, 1.204795916498, 
    0.579425331578021, 1.31305358829087, -0.680815827265322, 
    -0.490506059582989, -0.502870576573047, 0.0505878852122699, 
    -0.0134789429292947, 0.100868299032193, 1.13306376317418, 
    0.505148507581641, 0.901304945022394, 0.334733678132717, 
    -0.732475562492891, -0.98102373223421, -1.35955398169652, 
    -1.17770807780107, -0.896058197781424, -0.696591899784154, 
    -1.31531894838986, -1.09670677861966, 0.162252834041916, 
    0.0273868456475945, -0.419654222570625, -0.418342218296011, 
    -1.34480886065546, -0.9965322212358, 0.109465120723233, 
    0.449447148704758, 0.507643586877955, 0.583600536522977, 
    3.88825748640375, 2.0645739572637, 1.89791551559208, 1.5936831181613, 
    -0.758379123673807, -1.06343125187026, -0.804192125992982, 
    -0.394451093906634, -0.456646867960719, -0.31925156385932, 
    0.0475835655035706, 0.0714544719515864, -0.175105411894045, 
    -0.603407044700597, -0.360716196295119, -1.23400827793703, 
    -1.57500037175352, -1.17609869986102, -1.17691319693994, 
    -0.608708090976018, -0.733308124061103, -1.0989663590691, 
    -0.0700942094479773, -0.234527027746361, 0.0674672909630525, 
    -1.33816619344569, -1.42546879810105, -1.07870789132325, 
    -0.228417660891793, -0.314191269185429, -0.774405914454253, 
    -1.02061679485535, -0.920431304283866, -1.18497037261359, 
    -1.64914258313149, -1.50322445007338, -1.50120913278908, 
    -1.58103924003251, -1.1900932632822, -0.602144436397429, 
    -1.46151964611246, -1.6802252838788, -1.45345316405423, -1.1299917299983, 
    -0.634551451873979, -0.567013437401749, -0.964062146835558, 
    -0.527366309990485, -0.0977143766880761, -0.284056093389027, 
    -0.435734291110643, -0.843444516219263, -0.0243261579311405, 
    -0.325376688826147, -0.864774387021923, -1.03233663609814, 
    -1.58157631764089, -2.14021849153041, -2.51506600751655, 
    -1.60616245906295, -1.93258582400492, -1.87816010904749, 
    -0.76024350536914, -1.15714016245292, -1.60599507680367, 
    -1.33254622208207, -1.54680713801715, -1.1903166376327, 
    -0.841561850331756, -0.390028622550029, -1.16174562015425, 
    -1.15201685395934, -1.55884327425443, -0.864921719862912, 
    0.0107206770456125, -0.83387629485987, -0.995408311814572, 
    -0.659705274914915, -1.83363004217008, -2.2842021527233, 
    -2.86709595449253, -1.23394568206853, -1.77274464371402, 
    -1.45011711490401, -0.661367910456785, -1.46556144688295, 
    -1.10578099128577, -1.75079187746441, -1.8239634120757, 
    -1.04631246069292, -1.09817140903429, -0.781818356848141, 
    -2.14786911096678, -2.62347875473369, -1.12912050212065, 
    -0.650915072796638, 0.936286694745569, -1.24860707006134, 
    -1.05591361368241, -0.387990686879753, -0.569511737598294, 
    -1.49662671300736, -1.52664040919829, -1.30687493164869, 
    -1.74347892706447, -1.4207571784965, -0.696442460995681, 
    -1.47346605628884, -2.36123462013103, -1.76756424287679, 
    -1.23711457209459, -0.92745352498119, -0.890166624974289, 
    -1.13306202234686, -2.49145502802333, -2.63993540119001, 
    -1.05296815748523, -1.15319597397002, -1.12293082769611, 
    -0.774492193866179, -0.299030734429948, -0.397515092028975, 
    -1.12962581203837, -1.61283457019784, -1.62784929784934, 
    -1.34127401091736, -1.13863988666755, -1.66015361197199, 
    -1.75942880112256, -1.56707962663132, -0.989861459708505, 
    -1.17742140522239, -1.24644498539773, -1.16572409127576, 
    -0.793495212896556, -0.90269920937017, -0.790549512571719, 
    -1.07046295863316, -1.37817532288016, -1.11223521288879, 
    -0.923230195477562, -1.68689009758457, -1.77700454453141, 
    -1.44135850606868, -1.16510789722093, -1.09629357763609, 
    -0.754078291810494, -0.927465952943174, -1.81141115957664, 
    -1.40689776715901, -2.00028794955097, -2.03656726901753, 
    -0.8567017271307, -0.97465097793545, -0.854553274730154, 
    -1.36339612219772, -1.39829647634276, -0.689800698771661, 
    -2.45740080551664, -3.31458501640432, -2.21847004561811, 
    -0.202438361696413, 0.0562817353637479, 0.44746123029471, 
    0.593875500153387, 0.436594775248871, -0.124817127578054, 
    -0.507343565962795, -0.869023285322132, -0.964695487022373, 
    -0.845433680154226, -1.37248947929489, -1.63013603395808, 
    -1.05425636111248, -1.99866967381472, -3.63060386359508, 
    -2.29129855835259, 0.367795445502415, -0.311225452153527, 
    0.711346004638505, 1.70019540267168, 0.220321979484037, 
    0.230450909423232, 0.433458315596975, -1.32736580710181, 
    -0.950115060411796, -0.188059351304255, -1.44737941684017, 
    -1.0818188956648, -1.66532387613284, -3.03331475455691, 
    -2.37811775955625, -1.08295143501154, -0.84349629223023, 
    0.445464417554096, 0.575576727563152, 0.583536252549415, 
    0.549854099528653, -0.632675243317236, -0.356788214418584, 
    0.384729586596788, -0.82630428958538, -0.65979699462539, 
    -0.494396996136253, -1.65878898539506, -0.940337955757973, 
    -1.06510200871203, -0.870108152441054, 0.0680813527799051, 
    -0.27691475537726, -0.208146720086155, 0.390027911743012, 
    0.57036213344956, -0.403708798991596, 0.23325630731005, 1.22265905825154, 
    0.897395369107721, 0.773178073511813, -0.591260430055383, 
    -0.233467572975989, 0.0287900316296064, -0.399339804166088, 
    -0.188206051636337, 0.404153493897921, 0.198519175965224, 
    -0.512448110729444, 0.54146828151151, 1.14345805012082, 
    0.281405702977877, 0.67098580309727, 0.0763228666504823, 
    -0.0465951627138139, -0.257794796561623, 0.502285791281403, 
    0.547084395313151, 0.0255811940794359, -0.283605144513519, 
    0.178733468528827, -0.169937459015022, -1.50576877915051, 
    0.0787609030906467, 0.634355057436622, 1.04215051441943, 
    0.435853570564033, -0.4842992657826, 0.244319228256291, 
    -0.401077388159261, -0.348768203088103, 0.659580100941941, 
    0.155009883208148, -1.7542658407424, 0.410300520297713, 
    0.357389431945019, 1.17625249641079, 0.409881175424309, 
    -0.382733236406239, -0.585530631206996, -0.360104965677852, 
    -0.197736486948639, -0.18776313872733, -0.829406563676098, 
    -1.33889786392341, -0.652237792189245, -0.429163660055654, 
    -0.405868390008028, -0.888518646108598, -1.21501092523384, 
    -0.562859398447837, -0.451724356996013, -0.624206247824461, 
    -1.70877972705889, -0.437438474622462, -0.830324022529183, 
    -0.972611856122363, -1.52706821419287, -1.64032648751388, 
    -1.18797141335881, -0.0876551668135894, -0.161685204611191, 
    -0.091332006552971, -0.380435503252046, -0.747343236313704, 
    -0.836501923800403, -0.489747331943873, -1.21272062846144, 
    -1.72974103760674, -0.164450854039511, -0.389721027498244, 
    0.151274323342512, -0.253831154262794, -1.08810931342324, 
    -1.67792576151414, -1.35359100251712, -1.15585945700906, 
    -1.02414330842699, -0.392994694124926, -0.873007741205951, 
    -0.741629198651403, 0.197868395941465, -0.726162403463504, 
    -0.708228188118176, -1.57449194631279, -1.07449663615024, 
    -1.07160143946225, -0.998634664496683, -0.952263097456862, 
    0.142878935680693, 0.732278296413624, -0.287885799890812, 
    -0.667700767091959, -0.761025732203021, 0.190134030511939, 
    -1.23937735434673, -1.01209359752449, -1.6077991520469, 
    -7.45172375188741, 1.1549513262704, -1.56050966376131, -2.31226245106552, 
    -2.98795750199713, -2.81111090763499, -0.466746653569539, 
    -0.511870795065024, -1.87952911879901, -1.92238871234138, 
    -0.825079229874826, -1.09701753747932, -0.2622892710701, 
    0.931889227675931, -0.476452786436483, -0.222723570464965, 
    -18.2237758790698, -18.3599023606526, -17.3642473444502, 
    -10.5752825194152, 0.0505198455966285, -1.04162530832651, 
    -2.04281640407443, -0.675441619762296, 2.85827534724632, 
    1.89618699084946, 0.415325613008122, 0.338249968275761, 
    -0.705057441346923, 1.20680539017926, 0.672549773824471, 
    0.607493441381024, 0.378200714263954, 0.322670338525643, 
    -0.399202907718177, -1.63900152592621, -1.17303291598988, 
    -0.51710048884912, -3.40970830068468, -0.467018583151062, 
    0.3392101309678, 0.934358086526972, -1.72181308727888, 
    -0.585827195744309, -0.317387938694066, 0.518135101874719, 
    1.80551983944772, 2.17562840528973, 0.500390431856892, 0.628584076649106, 
    0.842750897732496, 1.41608540445834, 1.24394704161474, 1.00084594199883, 
    1.71613259625015, -2.85929562008462, -2.71668796350895, -1.2407493468416, 
    4.21733397532975, 3.80021863820017, 1.65412244875495, 0.540354666074186, 
    -0.806590195496106, -2.49762515217853, 2.69476996200524, 
    -0.00454755118468597, 2.080046470995, -0.143791668033089, 
    0.891407444187564, 0.535687167042198, 0.301584279712586, 
    -0.43341343597163, -0.190935219748667, -0.126720949344872, 
    -1.02224302036404, -0.122035056365517, -0.686432637227181, 
    -1.66455208422828, -1.14430692790909, 0.500370563195691, 
    0.0378999480712672, 0.044090598823594, -0.415810930584382, 
    -0.813978427264486, -0.384647701072529, -0.139857488927086, 
    -0.368541112269636, 0.0443580264920485, 0.103669962707014, 
    -1.36747922875166, -0.297435342190382, 0.33199049811607, 
    0.407214105299381, 1.17096046156445, -0.212725377688185, 
    -0.219257333027341, 0.194040462497349, -0.243575952253501, 
    -1.0724149955779, -0.612285906815102, -0.328528435491946, 
    -0.596881489225849, 1.89455837140807, 0.457176749823316, 
    -0.333862065822284, 2.18229233470027, 2.95556564521055, 2.26805739071007, 
    0.307494671300441, 0.331716405795786, 0.736040107782001, 
    0.474192745018849, 0.631177485052801, 1.08085731747047, 
    0.441511526098801, -0.461741329306555, -0.413298631477401, 
    -1.23332753721181, -0.896951653945566, -0.813332167772818, 
    -0.840241443075724, -0.464616976759471, -0.180878003862093, 
    -0.354847633146358, -0.23739897262268, -0.276758647851154, 
    -0.507164662936583, -0.199096754877512, -0.617001367298, 
    -0.626677196804151, 0.0469033632164884, 0.336481838718106, 
    0.171338373549021, -0.628760843910703, -0.881559336892899, 
    -0.166997206561161, -0.288398818726918, -0.372794354580916, 
    -0.40706770671771, -0.334302744297736, -1.79497927029878, 
    -1.01235584058977, -0.043804132264964, 0.258387075970359, 
    0.568569225898474, -0.440127895766427, -0.55276245882697, 
    -0.274814893293844, -0.664423617332695, -1.33720261255344, 
    -0.833713398179148, -0.244488069445463, 0.398540875192674, 
    0.724692439186088, -0.248150008260835, 0.181304268049023, 
    1.12762560536495, 1.28283924635179, 0.205654845975096, 
    -0.915775297297574, -0.161191745282125, 0.0887809670620143, 
    0.225850258977713, 0.112885492472694, 0.580726583770934, 
    0.013648991380828, -0.378431988509953, -0.680608356901993, 
    -1.13697736271297, -1.39191071727719, -1.02836207287667, 
    -0.90125998767479, -0.208798259718783, -0.0966010759877056, 
    0.357878439517672, -0.215967795021919, -0.597025110004461, 
    -0.276692669455532, 0.0914095375165225, 0.117110537518581, 
    -0.896835968095173, -0.832222913528122, 0.166099705841551, 
    0.344498949346796, -0.647756836509412, -0.980839149113315, 
    -0.15542787174037, -0.573352823519198, -0.0588920151543526, 
    -0.89794187181981, -1.23413235788767, -1.39562959485276, 
    -0.470386820709643, 0.0672758789619277, 0.0752222758797583, 
    -1.25453269540299, -0.961796087251936, -1.16619449738739, 
    -1.34985324864286, -1.1640345860795, -1.19747746114812, 
    -0.27708428354746, 0.360152437505672, -0.0147749912578066, 
    0.01705771635697, -0.947379166610363, -0.809251601088112, 
    -0.204757741643187, -0.0408817613068413, -0.759607620674907, 
    -0.878343241708408, -0.272557639582951, -0.518411349132442, 
    -0.692579816182564, -0.407657487505233, -0.111047235369197, 
    -1.66107585630452, -0.572958695103107, -0.784756676406051, 
    -1.34757807923708, -2.3453568123257, -1.68945997419002, 
    -0.42849465687981, -0.260481709594282, 0.81535143421124, 
    0.195198738167499, -0.567123135925729, -1.21915100882337, 
    -1.06396669451078, -0.503290831198822, -0.649568022661011, 
    -1.30908624979284, -0.855837395505921, -0.418730345110276, 
    0.0927736131116408, -0.439722157076101, -0.615935688960523, 
    -0.448072122303662, -0.611857618642966, -0.0535661101310936, 
    -0.693711354535043, -0.968233965749135, -0.524065048560378, 
    -0.967980610614072, -0.0135622321135509, -0.870130791021166, 
    -0.321883838377932, 0.65618160751348, -0.293775051920782, 
    -1.27907702777557, -0.506262369144599, 0.0161447219231148, 
    -0.261132451744772, 0.660746073644152, 0.736499532104449, 
    0.230844281407814, -0.6301065078158, -0.0981264132352022, 
    1.05789722043785, 1.00507496307397, -0.0167186992290924, 
    -1.11287728236033, -0.0342067723577388, -0.793536501512944, 
    -0.166256376936396, -0.587915047769134, -0.482714060683995, 
    -1.43555728898985, -1.9083588742215, -1.35851185378755, -2.1631135455691, 
    -2.62936064593071, -2.02102026606515, -1.06021714909816, 
    0.0383032544393158, 0.0867570754738356, 0.00701303487605998, 
    -1.16546234562553, -2.41621602720318, -1.4815333077696, 
    -0.856168624804443, -0.594974544390441, 0.0140265579626142, 
    0.281904956158296, -0.588883460498035, 0.648220999197893, 
    -0.225691859215207, -0.57039376824398, -0.983067381726559, 
    -0.756377323489006, -0.269408122668331, -0.414376055875207, 
    -0.435028018731121, -0.374816308435784, -0.891288643378978, 
    -0.460476080222776, -1.46048271889587, -0.986376953445784, 
    0.0204079727918005, -0.280239763173391, -0.798277526722693, 
    -0.695458340272244, -0.0600508143526657, 0.590835919591886, 
    1.04327195599358, 1.08226240413248, -0.987325478367671, 
    -1.10134170080387, 0.0315078438391447, 1.58093637308858, 
    1.69186898975502, 0.670477775247851, 0.1249271131103, -0.545078588101551, 
    -0.710187058686538, 0.388495929240671, 0.50234479283513, 
    0.439342041861104, -1.46124840272273, -2.09101726354464, 
    -1.63770153753628, -1.93844854541482, -1.50663951150121, 
    -0.470346821848113, -0.162904011192171, 0.155151800585234, 
    0.132076417431222, -0.439760705782004, -1.30947407398666, 
    -2.14121893597568, -0.542940780140775, -0.286642279239988, 
    0.242644788714745, 0.197520409258125, 0.48820405863653, 
    -0.688983819250302, -0.223319221026861, -0.594608495892803, 
    -0.751331457253666, -1.21673416144065, -0.763925452844645, 
    -0.282083546016998, 0.0635915154594713, 0.370953579498181, 
    -0.141009377254755, -0.284038593728142, -0.0377687013293647, 
    -0.653591903531292, -0.93972087652054, 0.120745597271661, 
    -0.134210952738476, -0.0938910665582426, -0.281608452336899, 
    -0.0681027194511552, 0.605924431926059, 1.33239401025024, 
    0.731055102665508, -1.13251838453318, -0.844957162888118, 
    -0.334488442969074, 0.832576873318103, 0.620588769944224, 
    0.450370625010081, -0.571045622269457, -1.24680365096213, 
    -1.55415726279385, -0.677262200339595, 0.171544694991446, 
    0.622313859980816, -1.17112607857391, -1.84405270671736, 
    -1.48021422930178, -0.821647077315566, -0.828221220043304, 
    -0.170402317965039, -0.102071622433559, -0.0228334176160372, 
    -0.0658411194789688, -0.759976868064558, -1.1744842154514, 
    -1.82943555935563, 0.110541579250896, -0.578996895967645, 
    -0.568222283615434, 0.27310298161213, 0.248437962306403, 
    -0.878987480211428, -0.371843217421137, -0.401097137382349, 
    -0.506271603076529, -0.721577138662277, -0.464995940603257, 
    -0.470118525672163, 0.450886677354303, 0.219130390093687, 
    -1.38265281113069, -2.1320144511214, -0.17579304294573, 
    -0.571095267554576, -0.731371759221173, -0.866959966063305, 
    -0.526771731441471, -0.0188446982674861, -0.516154721894293, 
    0.0471492805734108, 0.607568636954112, 0.359997874081528, 
    0.339857189794026, -0.662047799656031, 0.452009082745337, 
    -0.147361024837851, 0.0124054720107036, -0.430646294628003, 
    -0.307959814936192, -0.381060228747265, -0.596347470778564, 
    -0.367138185391913, -0.112693896956508, -0.1646937395385, 
    0.54365137168682, -0.956536896908986, -1.12774670877263, 
    -0.955543955216704, -0.668382464884911, -1.10471902348187, 
    -0.414369511405548, -0.472851854978549, -0.583793822061418, 
    -0.535916794785014, -0.403327840926133, -0.506759110218122, 
    -0.985499135880752, -0.699989102799048, -0.790072038714369, 
    -0.508823065420581, 0.671406508335375, 0.0460166569248877, 
    -0.441468231570594, -0.30885860776606, -0.301331448365403, 
    0.164394864044755, -0.386977162848674, -0.997659176756169, 
    -0.656010136338661, -0.0511140493261086, -0.0328284385512001, 
    -0.892083737674665, -2.08413043084133, -0.387771108079358, 
    -0.733396645879614, -1.21220642558207, -1.04284479458641, 
    -0.433431146358658, 0.242096062687462, 0.305007898582543, 
    0.992367527000027, 0.281437366877983, -0.0575551803129359, 
    0.277269949181016, 0.171204851326365, 0.391163425281182, 
    0.554729676492536, 0.414304042035867, 0.0545476205401707, 
    -0.59575321517781, -0.739830853799548, -0.292727502143704, 
    -0.0586670028621761, -0.119057047961539, 0.275051493929195, 
    1.08478994079527, -0.618883235311363, -1.04381478770743, 
    -1.38257961395382, -1.01223697290855, -0.71991782599877, 
    -0.509675295113916, -0.267722520444678, -0.747438969554217, 
    -0.669793224861337, 0.221696280096531, -0.436718672372347, 
    -1.60371570016093, -0.648580260128959, -0.460913419307571, 
    -0.638246505796793, 0.113113238825706, -0.0132007329998984, 
    -0.0583924931215574, 0.135855591937855, 0.0244635635977009, 
    -0.0207067898847635, -1.35684030351326, -1.95555371243245, 
    -0.592741876487852, -0.76326090199097, -0.514646848530109, 
    -0.392087146280007, -0.0268566249318392, 0.0311307507441105, 
    -0.237154252899829, -1.31055911265728, -1.07200274544875, 
    -0.0322395046111046, 0.543635845972741, 0.748280384418685, 
    0.702748810097402, 0.0695303682493487, 0.269916629105665, 
    0.313585176361824, 0.585411846704611, 0.24688358452396, 
    0.191672591178347, 0.401132789754568, 0.365673308168413, 
    0.013517208748377, -0.354658951952671, 0.0480989913968077, 
    -0.870546835069486, -0.0311370704805025, 0.619184479204105, 
    1.0272148235789, 0.233729038823882, -0.853394484298104, 
    -1.94212194669309, -0.993057548590217, -0.506783180522272, 
    -0.448253320514191, -0.124644233737548, -0.712393801997271, 
    -0.121243052678865, 0.437228476482714, -0.429293357822645, 
    -1.90957696418527, -1.17483009521631, -0.345117374427568, 
    -0.0237180294066874, 0.415260911907369, 1.26229377232925, 
    1.11550505371848, -0.0163504946404558, -0.718408843780454, 
    -1.0856085986323, -2.01989505056313, -1.57266529929111, 
    -1.78282736469886, -1.65801214902175, -2.48865130779782, 
    -1.90445324032082, -0.216350835289515, -0.471101237150369, 
    0.151706564721579, -0.907720532917051, -1.00814862029559, 
    0.0377999641132565, 0.610784271744551, 0.909543593784723, 
    0.903312568351358, -0.125650110595896, 0.386206459804947, 
    0.418545068093215, 0.527385056231928, 0.78087297567258, 
    0.0198206218318564, 0.358682611848518, 0.521180807688477, 
    0.00262035641790614, 0.446401486600925, 0.505871098551243, 
    -0.394887718508596, 0.233989739708962, 0.367311842687066, 
    -0.636560633949554, -0.487347862175462, -1.57814001695321, 
    -1.04807524592681, -0.745517659216288, -0.716172967342597, 
    -0.0185978182293089, 0.072410517848005, -0.786254770282246, 
    -0.38768470846438, 0.259021702622397, -1.71588728292708, 
    -1.94044015692012, -1.44861954794673, -0.62087235243288, 
    -0.385056468133662, 0.619803824229423, 0.149462188564815, 
    1.00093740193936, 0.178005095519351, -0.285762777780407, 
    -0.761366714626357, -1.28854780402863, -0.813779541549193, 
    -1.69407159452188, -1.50532293852896, -1.78220554647454, 
    -2.42842500985595, -0.682842789554834, -1.20403068417266, 
    0.0378314022676474, 0.0309789458465426, -0.184108745613107, 
    0.0944111114127022, -0.158532874258834, 0.00629633322095202, 
    0.00304459307605587, -0.372137243316355, 0.473110498898963, 
    0.475706134921845, 0.743578524149822, 1.15396159910641, 
    -0.0839714905583813, -0.290943136186645, -1.14320242017928, 
    -1.03905657651451, -0.702666087579629, -0.726608251550256, 
    -1.06797955354735, 0.515923198457622, 0.6503711633147, 
    -0.733240588215782, -0.690679727316503, -0.854748715082283, 
    -0.585983437637383, -1.1409560731024, -1.32261092138816, 
    -0.758625480256216, -1.17697604538372, -0.707568496868518, 
    -0.628234294550092, -0.692160789656318, -2.1555655050674, 
    -1.80987256030743, -0.93522250275675, -0.414014086529368, 
    -0.212920341125864, 0.0147785070993667, 0.146335910819815, 
    0.0933057785824687, -0.245618070789977, 0.0110612005868393, 
    -0.552997701672475, -0.922677559352834, -0.471854178976905, 
    -1.08330573662445, -0.749328868230132, -0.293414678383614, 
    -0.680923466550993, -0.375503288366579, -1.19048773739425, 
    0.224279376882248, -0.285525925384262, 0.149380709232227, 
    -0.0399868645396007, 0.266537807390113, 0.185123498813895, 
    -0.24305525927613, -0.264433060289111, 0.541465514441861, 
    0.696532196178867, 0.190178455553802, -0.194090655288637, 
    -1.77886425792594, -0.107733256618254, -0.426262100553063, 
    -1.55787494347619, -1.9434219843665, -1.70030686881483, 
    -0.829174428303054, 0.021668313435641, 0.385883053487857, 
    -0.616465804434347, -0.889284051884949, -0.819407223344251, 
    -0.757416088290688, -1.3658482993996, -1.84053428149888, 
    -0.9266515135204, -0.86410119704905, -1.18383393919303, 
    -0.0184083636838418, -1.58088504517908, -2.30129061051092, 
    -1.89432488086285, -0.584492684444271, -0.569214406980683, 
    -0.223962767834855, -0.165731385114638, 0.0944800533832169, 
    0.517724316370165, -0.232495607694752, -0.171761971401878, 
    -0.848710731780491, -0.813521521327836, -0.676971257731656, 
    -1.1524783393861, -0.554558754148515, -0.622896800790493, 
    -0.751422538909652, -0.0560810273856172, -0.550942863070261, 
    0.296368643022991, -1.56853641632664, -1.46693778162269, 
    -0.767352775725043, -0.125985105842186, 0.566443367862686, 
    -0.0684406039673213, -0.421468003093164, -0.886860823168814, 
    -1.05238434640474, -1.05906602708475, -1.46916713568187, 
    -2.34578423173616, 0.281586162715959, 0.936085881280446, 
    0.402920436265681, -0.371216416292683, -0.357664331248326, 
    0.530525111921234, -0.585127042854334, -0.24553790760713, 
    -0.897381993933655, -1.3703182663187, -0.979541164135562, 
    -0.853958890429842, -1.36008598092804, -1.01496300549311, 
    -0.676566887221992, -0.886952516208281, -0.309805794004481, 
    -0.114222917264085, -1.78910795038365, -1.83461779611846, 
    -1.34708330733599, -0.57483918826617, -0.999044400488183, 
    -0.764240148698843, -1.11562894873226, -0.343451319372505, 
    -0.759289906383396, 0.112411994963999, -0.840942815431545, 
    -1.80006640656648, -0.992860611656954, -0.882575458418944, 
    -0.894633817835069, -0.59863479794303, -0.687973135307738, 
    -0.884066136882047, -0.252649174801927, -0.256507501683321, 
    0.460427378065402, -2.04275606500964, -2.52133162159865, 
    -1.52126629369095, -0.227035815270216, 1.24462576184849, 
    0.0104264758549322, -1.05947103757742, -2.30836493131618, 
    -1.01109775605904, -0.242710449757761, -0.74448629235182, 
    -0.871212305488632, 0.44504658361562, 1.28568634789544, 1.35400955520225, 
    0.969345848079803, 1.40057157690073, 0.442566202014323, 1.50235163360633, 
    1.078070241411, 0.832695232783189, -0.0189454272741063, 
    -0.146378088032204, -0.410086262625029, -2.189189341371, 
    -1.09735046340608, -0.493577344755201, -0.352199926335001, 
    0.701187041709104, 0.0490887098363279, -1.18468101751835, 
    -0.89271590198702, -0.465479793863262, -0.911238012773294, 
    -1.136113946029, -1.46556956004475, -1.38173676754048, 
    -0.592019684509575, 0.591921007675564, 0.243146045484313, 
    -0.414131897574719, -1.50719774846268, -0.44332698135281, 
    0.235598069555709, -0.54438350516226, -0.832591137780545, 
    -0.858071725263807, -0.589883855367956, -0.447507172117745, 
    -0.769381997823997, -0.0279850652158009, -2.18833701325796, 
    -2.30374787435426, -1.28086806477445, -0.435379812961383, 
    0.834031842720817, 0.028049491995672, -1.73052526935489, 
    -2.35480907646346, -1.00869947620298, -0.221018920664879, 
    0.206504128803218, -0.0625131097836018, 0.196904891943555, 
    0.847916094188972, 0.677011882036158, 0.0453743319796285, 
    0.697882390592843, 0.336427282127367, 0.727960015399685, 
    0.619535901368886, 1.06490371961112, 0.343067038472835, 
    0.222022178153019, -0.0961572239550446, 0.860353045452322, 
    0.569308061164935, 0.245372174027092, 0.516204581061142, 
    -0.383777664810716, -0.0701675052309536, -0.188286580623616, 
    -1.40223051396461, -1.38357845106018, -1.66086687660495, 
    -1.46313364039005, -1.40543865228852, -0.475410570772334, 
    -0.377274934120209, -0.641555633266471, -0.929642053224762, 
    0.636545914034436, 1.19429095812019, -0.107269033798221, 
    -0.843746854867335, -1.44035514073422, -1.10447968722792, 
    -1.23764213019497, -1.12982186469018, -1.33695492852234, 
    -2.10163990975778, -1.58716963792356, -0.965062541201465, 
    -1.44090223895017, -0.535408733342138, -0.00954810427038932, 
    -0.825389019998908, -2.25718380698063, -0.800778624748673, 
    -0.147598156429791, -0.868310671324588, -0.865382232295704, 
    -0.475741002094181, 1.41759245073229, -0.286942752789336, 
    -0.855725452593177, -0.734658180900655, -0.251098871748239, 
    0.612735992135396, 1.52771142559161, -1.05466187810588, 
    0.385220021414852, -0.104307214935075, 1.27539463017973, 
    -0.152704024933499, 0.603654879524607, 0.104490661239214, 
    0.576575324856607, -0.183376167775043, -1.1030918124498, 
    -0.286248134923742, -0.518264121719687, -0.283326674553046, 
    -1.9088026310761, -1.69447065758727, -1.71424527143865, 
    -1.80124202458332, -2.16284403657934, -0.436539529970004, 
    0.905907727256272, 0.00296678505675274, -0.867335680446444, 
    1.14920869976867, 1.91418437956299, 0.742892916838054, -1.42764248123069, 
    -1.76967771395208, -1.98925307980979, -2.10190046466492, 
    -1.54863011701942, -1.804293152669, -1.71400548583373, 
    -0.856636288473349, -0.414447449488571, -1.11839513254329, 
    -1.37486335002578, -1.00063658029231, -0.773255471188041, 
    -1.60143691418931, -0.066871160430213, 0.110734515343647, 
    -1.03326239615232, -1.10813526108437, -0.532527142696919, 
    -1.1175003706309, -0.653391758869495, -1.2370574738289, 
    -0.509206230374026, 1.52760503204854, 0.537970260447276, 
    0.448748948718394, -0.0399610403530293, 0.448473604704072, 
    1.04137376555847, 1.10239165888267, 0.155261351179101, 0.07846649065407, 
    0.593900093579387, -0.304034090322353, -1.17502207746918, 
    -0.642204887970487, -1.58515241529638, -0.57794116907556, 
    -0.799218416531913, -0.927991007809741, -1.02334767293108, 
    -0.420965675105838, 0.40304204730484, 0.106350984375521, 
    -0.775880167458034, 0.898453532928944, 0.23405840303024, 
    -0.131380034297344, -1.63867958873223, -1.72143892032983, 
    -1.24468305541834, -1.33591358347165, -1.74660141492426, 
    -2.09473710708139, -1.34658150914164, -0.906976940234947, 
    -0.443325423062748, -0.586486723870747, -1.4386674882, -1.68892717409849, 
    -1.1519289776915, -1.28372520656943, -0.609161208743836, 
    0.0911641237888761, -0.35380263909182, 0.245300503465592, 
    -1.22489266100796, -0.824471070053226, -0.277322427991291, 
    0.693147457732003, 1.6122547860223, -0.467717176012231, 
    -0.0438192773964996, 0.568488023634219, 0.341962649115305, 
    0.36946706569061, 2.70045356914801, 0.723189303119036, 0.122991702417764, 
    0.586577683017593, -0.929120103223919, -0.764546908662957, 
    -0.836321417351575, -0.134937544456273, -0.00906967187511931, 
    -0.039938426793622, 1.06751381012227, 0.66483950706802, 
    0.821609819157265, 0.314055282505059, -0.975567598223688, 
    -1.25331647714463, -1.56767555762906, -1.43628757695642, 
    -1.25348052730138, -0.978916252469375, -1.67168883520357, 
    -1.58409100535151, -0.482670354911305, -0.540562666241002, 
    -0.592178055159129, -0.63277284061821, -1.59771167314705, 
    -1.28201701350812, -0.144256514587169, -0.0545907423215786, 
    0.390273707446864, 0.376298387829457, 3.61737365149649, 1.59529129892239, 
    1.29188882022688, 0.840006548281096, -0.837591357178074, 
    -1.26767912764337, -1.05123013038254, -0.487960148380262, 
    -0.568644068841833, -0.435639345073642, 0.145429226402287, 
    -0.194252813855216, -0.926835571218803, -1.22812608212722, 
    -0.588749223546232, -1.57092505802562, -1.85880913702747, 
    -1.388789292022, -1.45836913971242, -0.936225646790736, 
    -1.06050360040364, -1.51945155000551, -0.698496794093986, 
    -0.629395419879515, -0.22960862264056, -1.57558800402626, 
    -1.76506663591036, -1.31927009294601, -0.588025922722539, 
    -0.287543926777625, -0.825051597678863, -1.13921054677286, 
    -1.1125167957922, -1.40450770757704, -1.89322822286264, 
    -2.08143000619336, -2.2178062362965, -2.14820358489212, 
    -1.30847732929713, -0.723906840294832, -1.72734733654666, 
    -1.94307606576805, -1.71854685951832, -1.40082041298366, 
    -0.849831453154177, -0.872115631463242, -1.36510799825656, 
    -0.964539710200563, -0.503028556916321, -0.568877255647657, 
    -0.739131493659535, -1.11577103253509, -0.125610920760484, 
    -0.596479218945616, -0.987124507036281, -1.21126169292369, 
    -1.87636717089425, -2.41809620528194, -2.76486525187578, 
    -2.08999185055794, -2.48696759093471, -1.98507699586537, 
    -0.986166117751814, -1.51219488499693, -1.88799971917142, 
    -1.70820696220861, -1.82743547346644, -1.4444824559903, 
    -1.07794010112466, -0.786376603217902, -1.7257992711219, 
    -1.6165661367485, -1.94694088014659, -1.16343238393197, 
    -0.373801897697752, -1.14710811303012, -1.24694532949931, 
    -0.961600503144373, -2.24102714270311, -2.83392568672321, 
    -3.07430892021674, -1.50428353738574, -2.1585403840511, 
    -1.57762382578472, -1.00532214242412, -1.87057868147796, -1.616954233201, 
    -2.15073312476441, -2.16071455643484, -1.31697006315528, 
    -1.30312983843675, -1.29875656970533, -2.88627832966537, 
    -3.0393865337616, -1.48303321029209, -0.756290082890607, 
    0.523864095784692, -1.35173000040942, -1.30574718013144, 
    -0.649713621044787, -0.903054030914148, -1.96315221392115, 
    -1.87034312450369, -1.48948044628171, -2.06671281493046, 
    -1.68540999062783, -1.26694237405361, -2.17792098147897, 
    -2.7516443119134, -2.10115589384665, -1.63947873943284, 
    -1.28339724140757, -1.12150394162363, -1.50663337058815, 
    -2.87776418180981, -2.82632788802036, -1.58766492318627, 
    -1.18058067483397, -1.38393767471119, -1.14876656152392, 
    -0.405781514418084, -0.742518237473382, -1.49845585292069, 
    -1.97913884357224, -2.07935600885988, -1.71364308041032, 
    -1.68596253725113, -1.98545187334658, -2.14752515746061, 
    -1.92988833806852, -1.4236349887093, -1.50933948067887, 
    -1.59606748074641, -1.62060191392117, -1.30224388977426, 
    -0.672714227280773, -1.06443448981394, -1.4512858359558, 
    -1.82135299958445, -1.5667155940976, -1.22563604288557, -2.1635278593911, 
    -2.79365137399998, -2.12367558757631, -1.68998951531789, 
    -1.39432363207209, -1.05582516196181, -1.28024283879674, 
    -1.86707362060903, -1.66976241899638, -2.19292841848624, 
    -2.17803586069674, -1.14562603740819, -1.32507976333252, 
    -1.39037681695437, -1.83225446359723, -1.77489927040784, 
    -1.0385078055251, -2.80043352582448, -3.82731817386116, 
    -3.02742059114323, -0.694949404932284, -0.38732155050262, 
    0.103603805294417, 0.33177636584905, 0.154129824432965, 
    -0.330263666456738, -0.601021851846788, -1.05435744424594, 
    -1.48924849623702, -1.28944345711986, -1.53920283685121, 
    -2.0490401001442, -1.35835996417774, -2.5111086802207, -3.95802353452326, 
    -3.09563478889888, -0.177972802344581, -0.776098858932666, 
    0.112278158836512, 1.42802683841198, -0.0817898216994095, 
    -0.225435109634229, 0.200265589247239, -1.88744592138441, 
    -1.11350143917196, -0.365119087780381, -1.88409557284856, 
    -1.41988185750335, -2.13756400949185, -3.66092295860982, 
    -2.94866291632403, -1.55523030012202, -1.38511672083794, 
    -0.092447795140167, 0.342480568502928, 0.39710811604158, 
    0.249239250667475, -0.999315527435014, -0.519919534400435, 
    0.0437581776131246, -1.55959089023368, -1.18340414283777, 
    -1.055223303438, -1.99954651842192, -1.36153109273313, -1.87045418478942, 
    -1.3867417027381, -0.306496104463916, -0.640767226862722, 
    -0.591383476531355, 0.166825834691009, 0.0692831507388147, 
    -0.831798638452463, -0.0161387256602152, 0.995504341609501, 
    0.329049488406916, -0.0227214483084293, -1.41869050308607, 
    -1.00079450243184, -0.406412157880061, -0.782780872459008, 
    -0.475419559399732, -0.102097189069648, -0.381490279789349, 
    -0.731438908587196, 0.209979808386875, 0.760567567852282, 
    0.00532115475169181, 0.120051728858308, -0.492415283491039, 
    -0.420149770827836, -0.706967376140031, 0.288847361342826, 
    0.208438073386104, -0.428639376514153, -0.605488036313129, 
    0.0508491694251267, -0.495836315811902, -1.82526585014858, 
    -0.175689474837566, -0.0153702948256385, 0.536145519951252, 
    -0.0933139776669023, -1.03194467674425, 0.133713443200776, 
    -0.538082549391721, -0.564996572040708, 0.262134114238801, 
    -0.318795644495147, -2.28326253894544, 0.141269363030259, 
    -0.0203401282751292, 0.619043261429639, -0.206108326728618, 
    -1.21600048832527, -0.660917381531263, -0.40479922057524, 
    -0.526944959451296, -0.81482998146825, -1.38131054108369, 
    -1.87279747941476, -0.990603326631048, -0.977935398730141, 
    -0.889770313556881, -1.54602124030876, -1.71159110989246, 
    -0.930559307506238, -0.855531812771519, -1.02242654446115, 
    -2.12265735491841, -0.74335627304094, -1.14611915819304, 
    -1.27274791567797, -1.75857535191926, -1.95317540469514, 
    -1.44997351576889, -0.53107753016068, -0.528024694776161, 
    -0.36169271077434, -0.838475546811717, -1.05260439624056, 
    -1.23191274588105, -1.06764615785679, -1.40521547120239, 
    -1.92473185605695, -0.366492652613859, -0.724065524584852, 
    -0.194434725193209, -0.306954344573889, -1.27163319485449, 
    -1.91806683438237, -1.85255454299076, -1.55183678587246, 
    -1.27254884646264, -0.621737478942856, -1.12878082093479, 
    -1.25152620466368, -0.137986353847861, -1.05267610290944, 
    -0.902488076208057, -1.5999303207377, -1.11479377693577, 
    -1.39696255809736, -1.3453732274277, -1.40105963923991, 
    -0.193956177249093, 0.463621990588594, -0.709763533946313, 
    -1.11222770071554, -1.66147667616262, -0.229160948882878, 
    -3.77105452402137, -3.64153020088867, -3.30385136315391, 
    -3.41612406009371, -5.61048437472182, 1.6326439187813, 5.24990762355442, 
    9.08734595404086, 1.5601451341483, -2.76482718210268, -2.52643613200492, 
    -4.18180489800997, 0.443576951263243, -2.08184100572137, 
    -1.81257776044387, 0.175950782436765, -0.444994492655608, 
    0.1730318075266, 0.233227934005047, 1.20082398787433, 1.51012543466631, 
    2.42116931300134, 2.62982955144554, 8.25346043597008, 7.97714089270016, 
    7.54914633502395, 8.00652473033736, 12.5574875500504, 14.1220350849387, 
    -1.34040319347193, -2.24851853805887, -10.4710522936223, 
    -8.20528628658934, -0.222783614132993, 0.124987836649382, 
    6.39288125993787, 0.157132586906528, 3.60819693543419, -0.24862729742452, 
    -2.13455865328172, -1.65311076580892, -1.93881150215702, 
    -3.80033000833677, -4.05523232682725, -3.16038659395943, 
    -4.37357450504265, -0.513462456703238, -0.1171367862122, 
    0.23092139468174, 1.41960757190366, 2.52352377820365, 0.81581670816848, 
    1.33328649657611, 1.94467607655501, -2.90265863438158, -3.40186773751047, 
    -3.76980340716541, -6.75731957579704, -3.0832003954084, 
    -1.50985958349493, -2.04446613134764, -2.17378657394058, 
    -1.29751951755857, -1.5146376667222, -1.30224188477014, 
    -0.668896879269871, 0.327344345320455, 0.0748327872829568, 
    0.944000101858309, 4.09893408310893, 4.59595569083433, 5.04417042684437, 
    6.30310182925413, 9.3489769364453, 3.93304405156876, 0.114078261162438, 
    -1.08314194634066, -3.25574067062436, -5.27689986361249, 
    -4.2666823786341, -0.746961787702105, 1.60184302827133, 4.03268417462002, 
    4.20759351986391, 0.892124536425598, 0.777443219682539, 
    0.686714399096644, 0.7942504017727, 0.734055766094599, 0.320638190335387, 
    0.622438365614641, 0.307748214679293, -6.39672578829539, 
    -17.275179202341, -9.85078858485121, -4.73111820031566, 
    -3.99017398837472, -3.47673379403812, -2.22851819428907, 
    0.645922815453888, 8.75434242953336, 7.64775620163926, 
    -0.582422304211203, -12.4398739110898, -15.0181970128226, 
    -8.90418125195007, -7.50286013988583, -6.57498613515374, 
    0.24231431558853, -0.419649069009438, -1.60927930998131, 
    -0.819968549193311, 0.74458919930473, 0.14693230791134, 
    0.108762799688726, -0.490217829720683, -0.599824415196144, 
    -0.26141915315419, -0.219349715449564, -0.364927129546126, 
    0.188159132073573, 0.312750196602227, -1.37795361350634, 
    -0.281479889733083, 0.539203526185612, 0.694139151095508, 
    0.858776423124672, -0.0217564112775381, -0.592916151893341, 
    0.384374207517428, 0.0666831546252089, -0.465227420616312, 
    -0.607257392323155, -0.551665873858522, 0.175274486144059, 
    0.818414055478338, 1.21296474545987, 1.11876383160737, 2.03569743215456, 
    2.77664650007598, 2.31190599590151, 0.0704227663922419, 
    0.0514024783286704, 0.322002745625807, 0.329008520158252, 
    0.149961699740753, 0.470928039162835, 0.251834173942669, 
    0.679269201308244, 0.789589562347026, -0.309924305850671, 
    0.0870610580277109, 0.0261152667172571, -0.0299929047123371, 
    0.134196343195052, -0.134409936805877, 0.199553726924147, 
    0.408176215905267, 0.278159965775115, -0.260580804405448, 
    0.076383663241435, -0.995683226346875, -0.583282293829308, 
    0.0624748344150117, 0.329485141349295, 0.309015158348904, 
    -0.577938994992273, -0.781172901668761, -0.154714714077819, 
    -0.514855169613675, -0.569682073798869, -0.204912365595771, 
    -0.0171049896914566, -1.7806150553196, -0.900536381638362, 
    0.115364582967099, 0.286244899466279, 1.05415882820394, 
    -0.0872994855196652, -0.776324347111035, -0.260236958936484, 
    -0.00569666941212077, -0.896217085571696, -0.8418731760811, 
    -0.126010782023678, 0.412299476831719, -0.293422194536626, 
    -0.150950335306925, 0.662544058284431, 1.68228147604919, 1.6427309539672, 
    0.610973260346639, -0.822179601816329, -0.367267189907499, 
    0.182510021646753, 0.0672982463326743, -0.288877073198197, 
    -0.135867649364014, -0.385791552604964, -0.264202699424541, 
    0.36931509618126, -0.191199433480636, -0.722368811487013, 
    -0.514979824491357, -0.155693452892858, 0.45473566790831, 
    0.363500356465161, 0.749979919066481, 0.201434394102988, 
    0.0511782097402547, -0.173174050244942, 0.623894463414052, 
    -0.0981782511307561, -1.16109885823311, -0.966098243908506, 
    0.112841042752869, 0.305963670179343, -0.68387309728303, 
    -0.926906206670179, -0.153999034791212, -0.701544835546901, 
    -0.140947713540314, -0.0381005091685394, -0.906940227467081, 
    -1.57058307152644, -0.808524317433252, 0.250713328160979, 
    0.383609940791079, -0.581136423304245, -0.847933932794906, 
    -1.09445903883343, -1.29717486047927, -0.860025339437605, 
    -1.00657843714004, -0.538718874516779, 0.402464629364272, 
    -0.279069983402431, -1.17080143336334, -0.471553720289473, 
    0.413895420238748, 0.445041868416975, 0.0995295176420097, 
    -0.897090527836668, -0.750518896509842, -0.634928283861322, 
    -0.519697114150404, -0.486967476493732, -0.674175588824344, 
    0.0162894722456475, -1.22411983536568, -1.12212120944443, 
    -0.911394505757075, -1.01814029155264, -1.64578945930263, 
    -1.1887008396051, -0.00852181302720467, 0.399732973820286, 
    1.20564611818794, 0.678288076715927, -0.162434290794233, 
    -0.762099487098782, -0.605202197417594, -0.184248979090968, 
    -0.757658590835844, -1.49496645529706, -1.02474856659109, 
    -0.466434528652373, -0.223245482930574, -0.501757496575204, 
    -0.340722628898917, -0.286469644562555, -0.866311176619523, 
    -0.201714296015174, -0.369895371501059, -1.20921148186547, 
    -1.03463284399846, -0.801280916530129, 0.174514087192708, 
    -0.98976055801514, -0.61954600376389, 0.482624063146626, 
    -0.290830465543976, -1.58306617225458, -1.10487790610911, 
    -0.413370666082882, -0.451456611583425, 0.481857994458545, 
    0.0183339985131159, -0.643520722642075, 0.0176997641634902, 
    0.435673653068411, 0.747712451199138, 0.224125355589484, 
    -0.419148039974182, -1.07337541701432, -0.449035395205386, 
    -0.809964592775558, -0.305546369666869, 0.23195735651298, 
    0.450014493921191, -1.30181855580911, -1.99332452107719, 
    -1.67963960208391, -1.50853176518941, -1.52931408389318, 
    -1.5359428112036, -0.567420711478128, 0.53909278732053, 
    0.344176506612799, 0.799192990416282, -0.807572934275065, 
    -1.22553070822255, -1.22933944031239, -0.96356439697268, 
    -0.475022673722432, -0.207971446027084, -0.0257894766294342, 
    -0.850127708706383, -0.16478136093049, -0.547591124041924, 
    -0.662310527996977, -0.85802746532909, -0.976413071970175, 
    -0.229120123632733, -0.334817770287454, -0.736199885525513, 
    -0.657708815991613, -0.95603015185048, -0.675965579914299, 
    -1.79981155281177, -0.852994641828824, -0.00526353934283463, 
    -0.323753973295218, -0.699857543952871, -0.847654883358389, 
    -0.252957824711157, 0.271147706620694, 0.758786052713791, 
    0.429980277282285, -1.25668004032177, -1.09964148009033, 
    -0.160141026502503, 1.48095713672304, 1.30501972014583, 
    0.218782414558194, -0.471601916857853, -0.625725287613248, 
    -0.615258535405783, 0.355717861463973, 0.800473211074895, 
    0.935515990711959, -1.27575910061116, -1.48973129204706, 
    -1.98562292218642, -1.34764611795554, -1.11981457956363, 
    -0.0197022724876694, 0.195861595186124, 0.177197541218423, 
    0.244010776760226, -0.112536110496104, -0.952137366757304, 
    -1.27931833031887, 0.0497472530465703, 0.0244060883323893, 
    0.295159969184828, 0.0377197990483502, 0.129256950369134, 
    -0.900976237265363, -0.895351975768577, -0.684493934429939, 
    -0.424621108373029, -1.01395227765853, -0.539876007811078, 
    -0.141049758213447, 0.433722142201032, 0.187323794994367, 
    -0.303147469487532, -0.156957683584098, 0.0684816039066893, 
    -0.90740159643206, -0.793332072142876, -0.151257887004097, 
    -0.29399109310404, -0.172226170110537, -0.369516751852768, 
    -0.0210472789602933, 0.605038023566022, 1.11605357935406, 
    0.576170741445847, -1.03345383230641, -1.0618940561678, 
    -0.492170934469112, 0.602538061286149, 0.634414196548279, 
    0.231306579382164, -1.01816960768405, -1.03176210928414, 
    -0.901290532414576, -0.119423187760646, 0.157831451317194, 
    0.778873089267988, -0.399785055784561, -1.20681476251668, 
    -1.0776700066971, -0.620184665252363, -0.340751699390656, 
    0.0452131701052272, 0.49446419922206, 0.153895944117544, 
    -0.115548964096295, -0.200424022163901, -0.26045242660754, 
    -1.30566355277927, 0.45275737987386, 0.23438606345092, 0.375299760443113, 
    0.0162419185779772, -0.10432845200727, -1.22768761416134, 
    -0.757639450421745, -0.703208071151673, -0.470986577792631, 
    -0.52640416107169, -0.42115275260409, -0.227717857836125, 
    0.656281463761728, 0.0344005407779013, -1.60104850344971, 
    -1.75505040207723, 0.0751461290971639, -0.514239084293804, 
    -0.756828865518928, -1.11097383806121, -0.840292058786569, 
    -0.156962800786649, -0.307962770010137, -0.0965530467744458, 
    0.807348434540271, 0.682292347509654, 0.322274923257466, 
    -0.891368331332227, 0.445932123882247, -0.149135092187249, 
    -0.0510917838392588, -0.203353934133554, -0.245174154591736, 
    -0.35714527277491, -0.362221587918334, 0.329101780303698, 
    0.0686550842139644, 0.120907432105035, 1.25975568540608, 
    -0.69277898805737, -0.862818841156376, -1.13100353339225, 
    -0.401491379040806, -1.00939114529177, -0.260251455541716, 
    -0.207951833112117, -0.213013311168919, -0.0869860584148618, 
    0.0928872312390272, 0.612393250017793, -0.742544267944845, 
    -0.387784493819368, 0.548516477128933, 0.590359074490312, 
    0.643909275536227, -0.225621026725475, -0.925425147674321, 
    -0.590258992683972, -0.667231772837886, -0.164289537491316, 
    -0.551622123422937, -0.724381075728058, -0.31895850960491, 
    0.267884407888292, -0.0305410911115445, -1.79393221733574, 
    -2.28708442248147, -0.241978178153626, -0.762573689820329, 
    -1.35233362088191, -1.23854556400912, -0.638973382585717, 
    -0.0909237645289496, 0.0306869455207037, 0.34744383356113, 
    0.552705243506924, -0.0417166399392244, 0.267842194033023, 
    0.125668620760009, 0.30489082015714, 0.443829134030476, 
    0.513376809693828, -0.0756163133027821, -0.324434442387633, 
    -0.557123169717282, 0.00413793178578814, 0.162852884867117, 
    0.134977272033723, 0.642867683691586, 1.25341770027775, 
    -0.427651947378043, -0.778827927955166, -1.00435984550685, 
    -0.416225176360833, -0.465277422803663, -0.19701922912573, 
    0.352376895513524, -0.356404359325184, -0.200044579512744, 
    -0.0151505388464912, -0.211317896844568, -1.73005708048632, 
    0.465229229017847, 0.849123794135647, 0.382952326241943, 
    0.294087551410085, 0.076548879839109, -0.0336092654249676, 
    -0.0948743971044586, -0.227580563287848, 0.235519596371949, 
    -1.44343509926526, -1.37361308178515, -0.506704922285603, 
    -0.920079739768793, -0.287460220079505, -0.852015798268693, 
    -0.191546807066329, 0.0894208762519799, -0.271754988807729, 
    -1.46866500116437, -1.16370386039682, -0.237947329697752, 
    0.378698029373212, 0.414326209486369, 0.705226788652333, 
    0.245701675573122, 0.0199886089428691, 0.458048887385929, 
    0.530497696233407, 0.511222602009087, 0.223255450464386, 
    0.828474311055056, 0.449726391574443, -0.0367700344659827, 
    -0.15009550943164, 0.471036032907479, 0.316667745400507, 
    -0.0199730066661141, 0.63235170112641, 1.17129706183464, 
    0.290617561934039, -0.568169111673633, -1.64296358342745, 
    -0.877180749230941, -0.096128991845208, -0.269125701100772, 
    0.284033124203118, -0.291644810001097, 0.126390508845855, 
    -0.155476536778685, -0.844688290487362, -2.03377814441576, 
    -0.393865604828063, 0.553958091276492, 0.770890455840298, 
    0.601915674482347, 1.63404953659299, 0.982408220655957, 
    -0.25421088488879, -0.91939961845299, -0.851299909669043, 
    -2.23120501739507, -1.95238608366608, -1.58727454181976, 
    -1.63099917965162, -2.35637150735302, -1.74003126361174, 
    -0.227349424432207, -0.30027147897151, 0.172787928977001, 
    -0.984149362036333, -1.02498244324422, -0.129488398129554, 
    0.373793269430105, 0.841325902269232, 0.551928557254029, 
    0.0502156850786006, 0.125154558441953, 0.603843568162645, 
    0.486696243633169, 1.15258214782752, 0.667758149952293, 0.47842081339887, 
    0.180924786642609, -0.0136995239220106, 0.382702043891436, 
    1.07410663389442, 0.370989206957861, 0.349522923277723, 
    0.374982449285408, -0.333907685503845, -0.154710642546845, 
    -0.494748156721103, -0.870717240365151, -0.780176777245156, 
    -0.179149985905549, 0.269152878683552, 0.136515977760179, 
    -0.297005758271758, 0.358795131793621, 1.296582478347, -1.55497285989826, 
    -2.10486755375098, -1.51118677716774, -0.20044537040909, 
    -0.0710292105573482, 0.507421578899709, 0.520634929258472, 
    0.7910251911761, 0.195461556345338, -0.447379896548332, 
    -0.838242834610639, -1.53841146727069, -1.24536293687359, 
    -1.71373862886061, -1.5317933822609, -1.75277986647193, 
    -2.73961179540246, -0.71300183585291, -0.985499860549055, 
    -0.0406774797158915, -0.107591297256397, -0.331347410062408, 
    -0.138507364314013, -0.227723687897079, -0.00446108028891334, 
    -0.0659203077026271, -0.398234826501729, 0.201824159231263, 
    0.531956893282466, 0.796284481907334, 1.19425728806836, 0.6202524389697, 
    -0.0445916519976652, -0.540791367394728, -0.813717330143753, 
    -0.702882185498042, -0.490372841290672, -1.00175569303159, 
    0.443248406729255, 0.815908395423368, -0.532188028230514, 
    -0.578298373153125, -1.00036451126321, -1.15355016919053, 
    -1.07911138138553, -1.27508529975694, -0.74152558692874, 
    -0.56463948322969, -0.334282200748315, 0.13664782352, -0.674377540879831, 
    -2.28881023973121, -2.00235133769641, -0.791394258600269, 
    -0.28479044163543, -0.480548715845366, 0.0475689931832068, 
    0.147664813600006, 0.0725140624067855, -0.466478350725126, 
    -0.212300070235942, -0.697071176776332, -1.10966000533127, 
    -0.442051448984793, -1.30564951363593, -0.810342494800178, 
    -0.395623614778176, -0.955393597681411, -0.643097520035831, 
    -1.31428921496701, 0.0834917724655337, -0.539766424986765, 
    0.0671511664453517, -0.265485762407329, -0.0697326287320532, 
    -0.0838035223783429, -0.464531422408556, -0.437704618369201, 
    0.0727507024491603, 0.710605577698726, 0.331301139003086, 
    0.32591974423783, -1.12097586029707, -0.273053202463811, 
    -0.0551655616109281, -0.982236954850757, -1.84541858623184, 
    -1.96576198087816, -0.831795363845953, -0.174114655410516, 
    0.00122415117677743, -0.614440714590581, -0.812259923615719, 
    -1.13725329030011, -1.41715737783805, -0.986003526629031, 
    -1.76739909535536, -0.768878133682684, -0.509066258941058, 
    -0.577029594202489, 0.299834561238977, -1.65977969929281, 
    -2.45517668912723, -2.0157478664397, -0.334965689861173, 
    0.32976501851901, -0.303378419346432, -0.374179764663625, 
    0.593057625932767, 0.552676330687172, -0.308192016429762, 
    -0.451063953180104, -1.12885063424817, -1.08290886616261, 
    -0.307829187919144, -1.41192745682116, -0.667710337221084, 
    -0.815301531369061, -0.618358044855412, -0.226663067094681, 
    -0.686822336705046, 0.136701044663345, -1.7878386637407, 
    -1.65418655107551, -1.00400864182574, -0.327364136375063, 
    0.458662066243845, -0.247513027943973, -0.502133590594829, 
    -0.615174186833842, -0.949821049194517, -0.619988790096109, 
    -0.793232701676732, -1.94162565676436, -0.455053925757829, 
    0.623531360071392, 0.280184346503982, -0.793082214010017, 
    -0.31269306503602, 0.394381274136002, -0.513147012471986, 
    -0.403656536888297, -1.27047214671052, -1.56175765390534, 
    -1.25913504501945, -1.75162881289612, -1.63810468624617, 
    -1.18541562914903, -0.949043932405602, -0.276002201630967, 
    0.437153139343605, 0.132097720756454, -1.94798205933302, 
    -2.0238916164205, -1.5934002684704, 0.120225462909271, 
    -0.0926917241149727, -0.144156066235954, -1.6127737520074, 
    0.294141849167957, -0.607788080679592, -0.27436553238104, 
    -1.06193475433627, -2.22445796302337, -1.39622249246134, 
    -1.0569541014378, -1.11459374293055, -0.528540447718551, 
    -0.793819614112286, -1.00392379397267, -0.343708452694864, 
    -0.21954216106268, 0.406872134152239, -1.64820986070221, 
    -2.64971646410827, -1.48390398558302, 0.0493944037541816, 
    1.40536744586554, 0.0120220326441389, -1.12138722552106, 
    -1.60643780447799, -1.19814036429432, -0.702034644299174, 
    -0.857942179265305, -1.32365231888561, -0.387122121136474, 
    1.08587557495039, 1.00606494359279, 1.06148102052154, 1.0981760068802, 
    0.365826306737302, 0.750942671993537, 0.575129667445635, 
    0.324708068932482, -0.325016134134013, -0.714717415831099, 
    -1.82127484184102, -1.0929362102851, -0.308531091837354, 
    -0.0660006352529097, 0.474931606038722, 0.0540180041177092, 
    -1.50704850282159, -1.08777715291388, -0.645088906420637, 
    -0.197184817298277, -0.360315713510042, -1.02556598770852, 
    -0.960173820963215, -0.448731758342165, 0.408197591619404, 
    -0.109378805546942, -0.805126650851395, -1.88788268142142, 
    -0.51989380788219, 0.177287279078926, -0.681781332382725, 
    -0.758521297208472, -0.966972481605932, -0.747513782127744, 
    -0.542942117556815, -0.755153075361217, -0.116691308187584, 
    -1.9873591363626, -2.59570651698335, -1.31024657142745, 
    -0.446249331677371, 0.986424606778273, 0.266660459513965, 
    -1.91460416555672, -2.59465197194773, -1.45731116455938, 
    -0.326729897087521, -0.272719647572299, -0.47850698907892, 
    0.389771969753783, 0.957164391812046, 0.39440094618314, 
    0.127084642169396, 0.156382072222918, 0.36637270549098, 0.54562782804783, 
    0.470398759600967, 0.865748320165451, 0.719647218690653, 
    -0.360764745869426, -0.380631783935117, 0.437079099426769, 
    0.654722052856561, -0.0603052558609729, 0.104547018605499, 
    -0.954553724615614, -0.456829989771306, -0.52031616679542, 
    -0.567111772211319, -0.76908919626459, -1.43475948284621, 
    -1.57167651050809, -0.823814812976575, -0.342697266385938, 
    -0.321172539677557, -0.925368068931069, -1.21109584558349, 
    0.442115618449574, 1.21535606461445, -0.163428161160626, 
    -1.00172830005033, -1.59483388618748, -1.21229640316271, 
    -1.52961743539819, -1.40143794378382, -1.49306323922048, 
    -2.00415384979074, -1.71811991511673, -1.0149880395904, 
    -1.29761315891057, -0.65377475751327, 0.0116118557487832, 
    -1.22194368782089, -3.24319056252059, -1.37271994564143, 
    -0.352873696707716, -0.972034322541866, -0.778028619372471, 
    -0.651736994697858, 2.01349837092393, 0.270449142873832, 
    1.42489702088529, -0.343331471269053, -1.5161127123518, 
    0.351114803435255, 1.36696787875276, -1.22873984780368, 
    0.0179764344156164, -0.412843815205135, 0.948927154708255, 
    -0.552856676872056, 0.563921251209787, -0.214433848736522, 
    0.149965389836799, -0.4810379008777, -1.59851484726036, 
    -0.443477430473658, -0.840648502499191, -0.355342737464809, 
    -1.02842947306478, -1.13754634069445, -1.02438254396912, 
    -1.64406135727506, -2.05549467500318, -0.573705100921229, 
    0.590596085958444, -0.220242305916285, -0.859148580638331, 
    0.799046926586571, 1.92903261228524, 0.72709170475084, -1.64464275661061, 
    -1.85707394210546, -2.23121092076915, -2.42696846593858, 
    -1.89250562604946, -2.05409428639169, -1.93529022267043, 
    -1.26594426419037, -0.514185754559162, -1.07344447264203, 
    -1.34841402471089, -1.31642097860388, -0.983203796522134, 
    -2.63870346735233, -0.810724897621881, 0.205607946724249, 
    -1.46010890027113, -0.850601760509763, -0.532903348119742, 
    -1.33945420919872, -2.86283122279451, -0.430938160407893, 
    0.317126454502619, 0.372027937851009, 0.359619991224882, 
    -0.308816914421426, -0.378794306892081, 0.540520524012917, 
    0.630569842954767, -0.422615075008559, -0.540188382560935, 
    0.325128546711176, -0.648870135169058, -1.56043073620898, 
    -1.08161428485501, -1.04191335563153, -0.629495106142635, 
    -0.577995447731325, -0.572495810508613, -0.696377967582262, 
    0.401916524157016, 0.231100857941886, -0.217120617775635, 
    -0.970993447866562, 0.705817673750753, 0.248162700918595, 
    -0.101413209280716, -1.81847127247529, -1.92610129099395, 
    -1.47342150421831, -1.70296691194386, -1.95808840758225, 
    -2.24574486228896, -1.65956059612232, -1.22789929168188, 
    -0.735889642982888, -0.707669619337166, -1.49581809762758, 
    -1.83365218126821, -1.41703202580998, -1.96686313679479, 
    -1.25172889099271, 0.106683592882821, -0.606464278816237, 
    0.231635947483768, -1.28376764837448, -1.4575105729704, 3.41473567507468, 
    -0.915936846790537, -0.48987515743006, 0.0399532492281418, 
    -0.244822511742797, -0.473394569341798, 2.14504405552535, 
    0.351316477126722, -0.232607288807187, 0.0930717857436527, 
    -0.588031364393604, -0.0236030513315377, -0.270729019136509, 
    -0.0268279350117417, -0.233965825852147, -0.0471809511843713, 
    0.658344782034677, 0.591016191315283, 0.777212865156578, 
    0.191487453821813, -1.1020910329381, -1.33420871973061, 
    -1.68056830817566, -1.45695670886262, -1.44851254876085, 
    -1.20375134666808, -1.76255896237713, -1.73323589192042, 
    -0.712079134676902, -0.882773505051433, -0.755266552602665, 
    -0.996429316288108, -1.88288864739772, -1.61872754372967, 
    -0.581785334168985, -0.233955867995834, 0.172603786547736, 
    0.44558307441946, 3.28976817135586, 1.24040095060379, 0.747451172819877, 
    0.295941110297546, -0.115309760526783, -0.131910117158176, 
    -0.458161909776535, -0.280632025399354, -0.460419943947974, 
    -0.205777461065306, 0.607019533666193, -0.314145725406161, 
    -1.3359927899275, -1.50444841969686, -0.776670707343432, 
    -1.77688862721831, -1.88888635065291, -1.41184701298521, 
    -1.5133451911544, -0.999166519908181, -1.22834461460649, 
    -1.6520903295985, -1.13557536061659, -1.05351741952074, 
    -0.488404843666297, -1.95062524989605, -2.07629002942856, 
    -1.54752730010108, -0.912192485396597, -0.200398897832104, 
    -0.491660551444504, -0.743860924890436, -0.743604668531983, 
    -0.808431418315521, -1.00088696901063, -1.89708753445718, 
    -2.59727027600959, -2.51096830896734, -1.44493357052367, 
    -0.866015496554779, -1.99811010717811, -2.0737467965526, 
    -1.89585453355699, -1.40679328793849, -1.24961321228135, 
    -1.01609739020069, -1.57938110664614, -1.52065500473067, 
    -0.811050613733495, -0.943159319350642, -1.04292440041319, 
    -1.51782112693093, -0.599637756181646, -0.561015997753707, 
    -1.03430420974173, -1.02871286417155, -1.51748448535881, 
    -1.72419859403014, -1.78650231728589, -1.54516301465612, 
    -2.36916962081839, -1.98849513704281, -1.18237184183756, 
    -1.6693746807523, -2.10249278597598, -1.91682213717213, -2.4627247592307, 
    -2.10570789970409, -1.31058729421026, -1.13611874269591, 
    -2.13899674669493, -2.26564923267109, -2.46564722943778, 
    -1.5259169045347, -0.768766317831897, -1.15237336200743, 
    -1.02722666535747, -1.282866472915, -2.30197393636899, -2.5639258986977, 
    -2.26551848261996, -1.08750907766259, -1.88692446229994, 
    -1.69407534797953, -1.10028434947748, -1.91947992823451, 
    -1.74049146817937, -2.70000059924847, -2.80394603044097, 
    -2.19005805691309, -1.48166893425608, -1.68578084478392, 
    -3.35552367958769, -3.58054451218028, -1.80418736926629, 
    -1.28999797203892, 0.337117599228485, -1.47219094834589, 
    -1.49273684690984, -0.87201557666738, -1.39302341644171, 
    -1.94469951319996, -2.11110057763049, -1.10610299700185, 
    -2.07186819239669, -1.76762804366188, -1.09128751068386, 
    -1.82813219470503, -2.22260712030433, -2.50325185224821, 
    -2.21503265506188, -1.91075402854103, -1.3338225244795, 
    -1.66772616269111, -3.07372488241988, -3.00921620923429, 
    -1.73823319573171, -1.25246899269776, -1.66080546550705, 
    -1.47300934328585, -0.81324809215257, -0.974482327945707, 
    -1.82851908064295, -1.57953781057436, -2.10536642968555, 
    -1.81046046481607, -1.40874028116846, -1.44912575759291, 
    -1.62351593478821, -2.48691853664435, -1.74507951280064, 
    -1.86934205617338, -2.21802851257663, -1.99469068283509, 
    -1.69298535708071, -0.747039894324608, -1.48403173842486, 
    -1.95606331075702, -2.28292750385635, -1.96797850045157, 
    -1.45422254485592, -2.46147871581049, -2.84833531523333, 
    -2.28933519132816, -1.86683122885542, -0.959693005916646, 
    -0.640446433837463, -0.92255085541157, -1.39370807628318, 
    -1.8058665714545, -2.04793161347421, -2.35367362191315, 
    -1.49617514467542, -1.4799836422095, -1.48281255205096, -1.8987654333238, 
    -2.33539215254463, -1.5952851205334, -3.13803164781149, 
    -4.07452026317494, -3.37679062763589, -1.02410828673196, 
    -0.40259325760144, 0.133153168237254, 0.59200312130363, 0.48576683690543, 
    -0.336766295047082, -0.517869930280574, -0.97123942056534, 
    -2.01093479355794, -1.45916652281733, -1.60737241091225, 
    -2.60196201150611, -1.55525442991625, -2.73064730063953, 
    -4.12046044337119, -3.33917179059943, -0.598265784828991, 
    -0.968140829486175, -0.266196276276931, 1.33489835622521, 
    -0.0231832922357178, -0.549622912968748, -0.211096177543899, 
    -2.25612764562725, -1.27926586889627, -0.493262216377794, 
    -2.35434265043228, -1.70241710059465, -2.36835873179472, 
    -3.88063916621177, -3.16796454369366, -1.92969787176665, 
    -1.68176822081317, -0.475086252368531, -0.0251903460658642, 
    0.41071930910173, 0.406632178586057, -1.37878967149967, 
    -0.581081169880235, -0.207449639171537, -1.77064750154888, 
    -1.55746702230976, -1.34916708256761, -2.32573777257786, 
    -1.70920396854349, -2.22681906027562, -1.62946235944332, 
    -0.490468220990388, -0.848841645680509, -1.03497163525802, 
    -0.0947969946391236, -0.297333976049852, -0.917861407115184, 
    -0.223440010816347, 0.733828272968537, 0.0679532470836364, 
    -0.169848383364268, -1.66929968349819, -1.10109221172294, 
    -0.558472879814498, -0.684702149500191, -0.946291719283847, 
    -0.620686378277195, -1.10147886920784, -0.907951838936083, 
    -0.0344649033335465, 0.643345131024526, -0.10973721371673, 
    -0.0206730833982416, -0.81324873787636, -0.581451365893551, 
    -0.890719418307477, 0.124234916425898, -0.298961354766893, 
    -1.08095958082685, -1.12877231354608, -0.251064769955032, 
    -0.93050792561018, -2.03604410568241, -0.349175032972067, 
    -0.370928541083835, 0.147587524796573, -0.237910167427322, 
    -1.22974977668099, -0.170826594729556, -0.878599379600424, 
    -0.916865994286771, -0.141037549393559, -0.96322311958827, 
    -2.69684762570519, -0.248950657719225, -0.452997103311761, 
    0.140867660628463, -0.410540083684694, -1.50599191395918, 
    -0.753457807994513, -0.885371895988558, -0.972678479810938, 
    -1.59317737813879, -2.13192541891404, -2.34294564625719, 
    -1.41326809868243, -1.52326995266649, -1.30362850276872, 
    -1.8019459062032, -2.01229438750314, -1.43956542396831, 
    -1.40751910100447, -1.50018427331941, -2.53181634259433, 
    -1.30887002380091, -1.59014246350432, -1.83570012715168, 
    -2.26731457995824, -2.24794749079547, -1.889361213558, 
    -0.318305227100706, -0.867097274422259, -0.432986971239346, 
    -1.23065605217402, -1.58009056929358, -1.74582508401137, 
    -1.63667231139216, -1.88498535621851, -2.27799570275991, 
    -0.253568495781824, -0.940916959001132, -0.289987643039482, 
    -0.230585382850723, -1.40434759588836, -2.30589844808472, 
    -2.24401975315022, -1.88288853966603, -1.68045199862216, 
    -0.691066493951968, -1.10391459693917, -1.85962390230955, 
    -0.812771588669094, -1.15976072325973, -1.2508865857981, 
    -1.85574648672434, -1.62662386661052, -1.58157052988631, 
    -1.7957846751738, -2.25226256075055, -0.840922993348601, 
    0.253857236984749, -0.930798813549143, -0.595654117905768, 
    -2.38951378328321, -0.0698255831869416, -2.46414006831358, 
    -5.91606840357928, -5.84135782038949, -5.24770246668172, -3.182288814572, 
    -2.04153396888525, -5.34278807943021, -1.35864296685977, 
    -8.08299460839507, -5.85960977303057, -4.42300047106117, 
    -9.4718766035028, -4.32973224234006, -0.317449997178728, 
    -3.32012332497331, -1.06866599687174, 0.920341717054125, 
    -2.79172025940768, -1.78829701917629, 1.37915953033347, 
    -6.85917661054006, -6.77767142840285, -6.27347296728553, 
    -4.56371207041299, -2.30402475707065, -0.63213485726984, 
    -2.14686678014273, -0.121393955335645, 1.16396039794594, 
    3.11880384654703, 18.8447289524061, 22.8377617668197, 25.964468031424, 
    23.5033845081495, 7.34263177040759, 7.5514219076986, 7.88592195962323, 
    11.8563840073456, 7.22052691173189, 2.42726427848297, -6.50073229714039, 
    -3.24279740026398, -2.42847896605257, -1.94449725369504, 
    -1.56898676335976, 4.26641745029215, 20.3375644295255, 8.35161650393662, 
    7.78073072614335, 5.71601207517345, 5.18986188552617, 4.79299439150367, 
    4.51863479140471, 4.86385602135329, 9.36662533492836, 7.67109175648031, 
    -0.324814220443918, -2.80763701704153, -5.36030320334026, 
    0.133202335536433, -0.495528498100741, -1.57148691109581, 
    -0.844696218019205, 0.745595429067167, 0.231121234801277, 
    0.187480467601828, -0.320313785400232, -0.319760914328029, 
    -0.117538090311884, -0.0563892812667444, -0.220706575443028, 
    0.454305730440847, 0.504641342044705, -1.29744673782288, 
    -0.309890105303472, 0.659687243900318, 0.728146863268511, 
    0.295172979283893, -0.263785374682932, -0.730565373494825, 
    0.39296661077143, 0.0913121595574973, -0.450348513085661, 
    -0.772644104530449, -0.751067606212414, 0.00689198791177681, 
    0.767853128764133, 1.55516563157792, 1.41085546152128, 2.4424623357238, 
    3.22045222689229, 2.62834546234848, 0.275591950552059, 0.679038778276646, 
    0.669240164150477, 0.552971599346415, 0.453170719945799, 
    0.540199279970972, 0.445194732395842, 0.548952033260344, 
    0.555816683935935, -0.432383627718362, -0.287842028226972, 
    -0.380823324522575, -1.39710636982374, -0.532047818039856, 
    -0.465479039110495, -0.271990075819031, 0.338302447411474, 
    -0.19401582978432, -0.182777878587732, -0.0251564929366754, 
    -1.09939333805414, -0.697534060006735, 0.0862336429264499, 
    0.581205078136326, 0.379551559886719, -0.347075565899688, 
    -0.462120100552488, -0.0467021383855748, -0.394026701282106, 
    -0.424259178408084, 0.0846985743862128, 0.224988245974829, 
    -1.65161539385713, -0.831974858825202, 0.21468346944201, 
    0.400633914818029, 1.00256526212868, -0.230319645328994, 
    -0.962465606820602, -0.154136874369244, 0.294318411529768, 
    -0.660091740161985, -0.951293093497618, -0.243603902385598, 
    0.428106782718141, -0.210703641078118, 0.406948283990292, 
    1.06926953065532, 2.00116269127751, 2.02233249092552, 1.07958619132628, 
    -0.479350066891513, 0.137736803079451, 0.683171033848318, 
    0.413206861337621, -0.122019373044928, -0.0294446849932939, 
    -0.0680228867976496, 0.0704093006170003, 0.268614346163609, 
    -0.276968253386922, -0.797464977634443, -1.32492021554297, 
    -0.938109232278763, -0.133916377283936, -0.476277605289948, 
    0.151389969056166, -1.00937337775433, -0.602915347757862, 
    0.191987250879277, 0.714640707624055, -0.220133944393437, 
    -1.19837933775985, -1.01489661472845, 0.21222290936163, 
    0.354796001566324, -0.442665649397203, -0.521283089661981, 
    -0.00215212093147343, -0.426910978528605, 0.0743344650176958, 
    0.154037963369098, -0.445365192440739, -1.58244491156144, 
    -0.797775881274365, 0.177018849646338, 0.353776645621067, 
    -0.390217529307466, -0.906135394243508, -1.13729261617287, 
    -1.15001809571237, -0.773370454934801, -0.841159671315346, 
    -0.453813642789163, 0.364906466074011, -0.318961770219746, 
    -1.24960079584205, -0.0587222580470703, 0.854638112940527, 
    0.499026330479801, 0.363090132473629, -0.679234339754795, 
    -0.330433200352012, -0.32883935206486, -0.0274661528369213, 
    -0.0964799805771621, -0.552147286236804, -0.0237154483914193, 
    -0.993608205173864, -0.911287742264397, -0.60735277198432, 
    -0.832078422847515, -1.59553441066299, -1.7170075612292, 
    -0.519945340426751, 0.109731063918241, 0.455104424481676, 
    -0.704801172137066, -1.17238750659978, -1.69102145411548, 
    -0.10661984784428, -0.0556394868516374, -0.850764279306917, 
    -1.51651819792525, -1.08392408042958, -0.410605686755039, 
    -0.14677967827434, -0.283946038613525, -0.00165112677112056, 
    -0.212777131928794, -0.606505650892002, 0.0242159278805598, 
    -0.234778199098344, -1.02411298596333, -1.08215235077265, 
    -0.707182964981463, 0.0842458290965986, -1.18933192027706, 
    -0.558177442495527, 0.582018637718429, -0.0174401182609918, 
    -1.30374891118058, -1.14175510968936, -0.502221934317659, 
    -0.269327924258151, 0.434209779395176, -0.34248153490108, 
    -0.931148163585593, 0.0265278645357947, 0.557416235642032, 
    0.945120036986178, 0.239525908884493, -0.312637796951947, 
    -0.790254657841407, -0.24048287268895, -0.530185114593458, 
    -0.363625511882018, 0.0724537513056855, 0.225315835130346, 
    -1.43376280187701, -1.7729458574801, -1.06931485534849, 
    -1.54436935136208, -2.13750541122125, -1.54442283003997, 
    -0.938109278464156, 0.332395580747922, 0.0329286172520149, 
    -0.0957473963801577, -1.82257545575254, -1.19178962727389, 
    -0.843528952355985, -0.714300771980945, -0.561510802516558, 
    -0.339864751169277, -0.0538097268112026, -0.852460055690383, 
    -0.15172849185765, -0.344056913773505, -0.409107265936424, 
    -0.783578160198388, -0.812077251608367, -0.0632467041668594, 
    -0.273720632893015, -0.83275934131839, -0.701603241629862, 
    -0.726740623501763, -0.877871937246968, -1.82592057617359, 
    -0.635321913452986, 0.069934411477468, -0.234750720446675, 
    -0.656151196607762, -0.875967370462085, -0.260211589337489, 
    0.339035814781461, 0.867353353280604, 0.0513826520993721, 
    -1.32675993783612, -1.01662731480936, -0.133391660131301, 
    1.5924819959368, 1.35963028270017, 0.329245512971603, -0.643287674347781, 
    -0.676682983774515, -0.583123914064756, 0.390083961274921, 
    0.869258193860984, 0.746976955412362, -1.58401182893479, 
    -1.61945516945413, -1.53212519561576, -1.56079959415058, 
    -1.25315422357803, -0.140648039204563, -0.101081561976035, 
    0.357199136068296, -0.155932101145071, -0.525057223444865, 
    -2.20234409814074, -1.28383423934564, 0.610719604781433, 
    0.922357879431724, 0.583274609516886, 0.533454842670258, 
    -0.0541113760541378, -0.997677028686415, -0.916133943571653, 
    -0.617586053169306, -0.306050071198691, -0.894524223322741, 
    -0.440820742307744, -0.0292312778468151, 0.511705317997357, 
    0.165214221240206, -0.0746674493356014, 0.259481789900384, 
    0.466953083199977, -0.845239939230376, -0.744154859557882, 
    -0.380697427722461, -0.404886681718688, -0.223829406979261, 
    -0.36772167898969, 0.144306441818598, 0.959411295993902, 
    1.32030406965734, 0.577561327294389, -1.01189734512574, 
    -0.849010957836964, -0.484758951339135, 0.710226529321574, 
    0.879063348759348, 0.333870323655896, -1.01661479923107, 
    -1.00344049760148, -0.839969575469555, 0.0462323608595261, 
    0.36589558807659, 0.917250700664769, -0.837685564347619, 
    -1.31108245317479, -1.18833704820668, -0.817681149923244, 
    -0.249884973573278, -0.01675505448123, -0.127476194748386, 
    0.117731820797369, -0.0427864345124496, -0.47522364039732, 
    -0.865038719769832, -1.40716065405702, 0.765562486012499, 
    0.543119969100099, 0.871859425800015, 0.00637314626272811, 
    -0.254108397399531, -1.52999748784323, -0.83467349552262, 
    -0.655703510868912, -0.4722895355789, -0.485531213221675, 
    -0.465249098075553, -0.149406527645306, 0.849394419994085, 
    0.200941762418489, -1.06770078125094, -0.82626664658533, 
    0.665655650977354, -0.389630884247238, -0.875790174944466, 
    -1.26978740143778, -1.04474205537773, -0.179968678753091, 
    -0.219262538481502, 0.0338493723674071, 1.2781679957994, 
    1.23188895189526, 0.528548543296514, -0.995575178188433, 
    0.40055027080832, -0.479312231318856, -0.0231886897715139, 
    -0.144517722865349, -0.140058597779404, -0.358985249986561, 
    -0.209012616297213, 0.409318664359257, -0.101990049624381, 
    0.116700498661171, 0.841715520185478, -0.406166002552344, 
    -0.752698476101505, -0.980244997922579, -0.708533820867792, 
    -0.844446166336734, -0.367265811840998, -0.641264423046279, 
    -0.178691257013552, 0.156970692997671, -0.233256324390974, 
    0.429597401143815, -0.458485810407536, -0.204423337148922, 
    0.379468176262785, 0.478645320874707, 0.648020536759919, 
    -0.238440278031069, -1.21749363506495, -0.746733915451072, 
    -0.787377178160895, -0.234414142750268, -0.672037634305216, 
    -0.770643315660613, -0.172428799745479, 0.436751942949196, 
    -0.184857280538666, -1.98710112774686, -1.76188880866209, 
    0.375804064477969, -0.620962638248215, -1.36909894335931, 
    -1.32932797855275, -0.623244690823332, 0.102373950374415, 
    0.0424678772887166, 0.182581234688719, 0.964537815497093, 
    0.511741137514772, 0.458987535996784, 0.13721813068813, 
    0.255063471281325, 0.347802208440102, 0.688178752437651, 
    -0.0941926950766137, -0.316317088563718, -0.359659464047648, 
    -0.00466161853335478, 0.191971527333408, 0.306309695468543, 
    0.700393079158341, 1.06836608735802, -0.341088824979243, 
    -0.645183177180177, -0.532437527545353, -0.603113597032854, 
    -0.917263269700532, -0.463465998937314, -0.258093587546915, 
    -0.37664153260049, 0.156376454723128, 0.212951201883516, 
    -0.318880662292576, -1.56138223446657, 0.399252349002772, 
    -0.103542494074604, -0.15269094516392, 0.705565353723845, 
    0.173348502564004, 0.0132915611348444, -0.293968241085105, 
    -0.370430338943355, 0.0333641659465167, -1.71846189741171, 
    -1.71180615505427, -0.603569268371555, -0.801692134411813, 
    -0.333957922632955, -1.40939766939487, -0.247436430406119, 
    0.331154385073855, -0.206213777289213, -1.53712480173621, 
    -1.27483091812265, -0.222781099778868, 0.423898714218023, 
    0.445570113379574, 0.70994840134857, 0.683452727242124, 
    0.296668018789878, 0.585090683707858, 0.713579893075353, 
    0.611953205503477, 0.314482179277698, 1.35848740791832, 0.48585453790305, 
    0.15144731179225, 0.0915311509547445, 0.319163055202938, 
    0.588715481251278, 0.585829589672207, 0.685052917489477, 
    1.24484444143674, -0.00140955183409286, -0.401248866170825, 
    -1.13000895929331, -0.96973690143578, -0.997181541583032, 
    -1.05068791469864, -0.482938089107083, -0.29467118605853, 
    0.669975994654131, 0.228303019839746, -0.808941530573755, 
    -1.55600976503519, -0.508587528439266, -0.0916759037615034, 
    0.0229792634561932, 0.821448233146018, 1.82515565252794, 
    0.78785874984594, -0.552718774810659, -1.12419830056107, 
    -0.936915785526309, -2.1777039747365, -2.35372876425957, 
    -1.76368701006298, -1.62793685165639, -2.11131098065867, 
    -1.6246902486626, -0.134331969757085, -0.123456639920825, 
    0.232757338168579, -0.947024907784675, -1.03574235264615, 
    -0.131561365799358, 0.488394861209684, 1.08711719760788, 
    0.708191916957168, 0.181029757063267, 0.262711856339011, 
    0.752434231447636, 0.6765610564528, 1.41082461638519, 1.05007024874407, 
    1.0139827824075, 0.562605524446953, 0.155545784404003, 0.740797784520666, 
    0.749984646391773, 0.705420067887159, 0.492547453375054, 
    0.0832827770968469, -0.5178325086891, -0.333463808266932, 
    -0.404474543641782, -0.375918744921373, -0.504692687409785, 
    -0.655385620317417, -0.192795767142111, -0.213480035897606, 
    0.240475839313983, 0.669469441749149, 1.85638866872471, 
    -0.769485682247577, -1.39202822280148, -0.932427191132872, 
    -0.671486575736546, -0.170805785343333, 0.208007159416104, 
    0.660645564575022, 0.715989215487456, 0.164738699820344, 
    -0.732696871553031, -1.12604688897718, -1.64864078337512, 
    -1.68537819453284, -1.97451397993767, -1.79543024487874, 
    -1.91745825449521, -2.75819610164409, -0.675446958610768, 
    -0.895876426147706, -0.098704231819422, -0.133929887450681, 
    -0.307677965506663, -0.256645288384054, -0.148820355322838, 
    0.133606183296702, 0.219291949258551, -0.0198951430876981, 
    0.43211034507737, 0.739073197058877, 0.733578584278769, 1.3727345945046, 
    0.711843338536067, 0.158901345996183, -0.510221574791334, 
    -0.571596090119115, -0.690431866551363, -0.655194923932811, 
    -0.836670398702468, 0.578777691548096, 0.907436167054647, 
    -0.536200370931672, -0.274548436527082, -0.676922049510038, 
    -0.481313948597153, -1.05324243896133, -1.26804181331256, 
    -0.372417846052024, -0.685071896923315, -0.0895289648036401, 
    0.519344399395383, -0.178539671915629, -1.45096157979293, 
    -1.65018312708257, -1.10372224315801, -0.234586604832794, 
    -0.426517124224617, -0.289668323874421, 0.166065243893705, 
    0.581212382566489, -0.789971687902851, -0.423004847279227, 
    -0.282674946206232, -1.35043820138967, -0.582446507041494, 
    -1.64066903155151, -1.06786727525668, -0.662838030135973, 
    -1.24476699645908, -0.853840330882534, -1.45857868849481, 
    -0.0234269810930687, -0.668444278901936, 0.138020527600542, 
    -0.505081582372333, -0.206394134236318, -0.228068761115714, 
    -0.470097725293095, -0.144739659837594, 0.13369417013263, 
    0.991994680938597, 0.861072355439552, 0.934542713487638, 
    -0.431584354174239, -0.40035396433181, -0.450308401303836, 
    -1.0208479932096, -1.64794922150064, -2.09843713927047, 
    -0.828317626735027, -0.101793995010571, 0.287827699438234, 
    -0.325452472596699, -0.385501815226679, -0.82302064369502, 
    -0.49998923793348, -1.14569176015471, -1.30426540421206, 
    -0.628767763747189, -0.713578813676334, -0.395612016432825, 
    0.768727581010231, -1.42683913128048, -2.02107920337747, 
    -1.53434124199889, -0.544497778925921, 0.203335652308372, 
    -0.34703450403903, -0.560291638707904, 0.293471789151987, 
    0.79258774862045, -0.335147237949363, -0.7159191234547, 
    -0.794499181862536, -1.32378590394511, -0.400990232520257, 
    -1.68528138231506, -0.963571903317431, -1.12159105287278, 
    -0.934500994503455, -0.411966928158161, -0.86057373766133, 
    -0.0142491705081227, -1.98666345064078, -1.72484575228208, 
    -1.12285580239601, -0.635708513319653, 0.117285781896479, 
    -0.600497022090107, -0.465208034960729, -0.12691452278685, 
    -0.557332566692454, 0.292229111002538, 0.366262636001546, 
    -1.02965259398681, -0.397650105597123, 0.401033651123548, 
    0.0787773658770297, -1.25088655681006, -0.708295673590018, 
    0.22684062319374, -0.0598821316122722, 0.00844435715937397, 
    -0.605599421539367, -0.97191227997329, -0.976582281266229, 
    -1.67807801400767, -0.76207232150713, -0.954057105758133, 
    -0.504706023294248, -0.0207494403395225, 0.272812590153193, 
    0.0779922204305983, -1.05363126682897, -1.54191348735525, 
    -1.24773357924449, 0.0158099949486346, -0.028082576256665, 
    -0.120020827167249, -1.00059065582821, -0.0404429820534702, 
    -0.467213779798445, -0.867336346003356, -1.33688583043225, 
    -2.25187836451129, -1.70708896299917, -1.1353632666924, 
    -1.46259539834359, -0.748250291463251, -1.17766096232192, 
    -1.32863556490701, -0.389356375081689, -0.317246158467706, 
    0.28316170204949, -1.66322762400713, -2.65907328714552, -1.555142500756, 
    -0.101887509367273, 1.2838170931196, -0.259069765926885, 
    -1.22391782667284, -1.2496937958573, -1.36548442921173, 
    -0.151329099656148, -0.38645368661459, -0.352379552405303, 
    0.607923731815622, 0.994921098824415, 1.07599576145236, 1.0137721905234, 
    0.918678078767671, 0.984603800475714, 0.309093171388617, 
    -1.49450172728686, -0.426722964978135, -0.271368446558728, 
    0.40464481501382, 0.0569855431295085, 0.208425460380459, 
    -0.0295492595264735, -0.927747305439497, -0.582573185119615, 
    -0.534933237588948, -0.532061076509009, -0.598084540312849, 
    -1.41897319967386, -1.3467895136657, -0.566408156509235, 
    0.173038953091922, -0.158777814115858, -1.78028273721559, 
    -1.93118951350606, -0.0578407364332278, 0.172048881701992, 
    -0.779569080902816, -1.07066577843268, -1.41827708002508, 
    -1.07622311003563, -0.673970645410926, -0.900886996822505, 
    -0.137998577651652, -1.94215767170869, -2.73310937552084, 
    -1.4362004941834, -0.657573056113527, 0.753714172590851, 
    0.0136135808356252, -1.96375273437889, -2.59864654057477, 
    -2.37330531395831, -0.368846413104653, -0.297363643069124, 
    -0.0439042984321736, 0.673464178235825, 0.710668260053846, 
    -0.0137337940599142, 1.34348638226708, 1.60000222531914, 
    0.639935048580953, 0.345620503765374, -0.0691726552290373, 
    0.238820272892494, 1.21682950806643, 0.317758210548016, 
    0.244204141432953, -0.736367054721239, -0.666973912649418, 
    -0.534915966287874, -0.072137757272297, -0.747526619723082, 
    -0.988788858658429, -1.81479281586296, -1.88387646401172, 
    -1.0303624650665, 0.102983429363279, 0.163609429030336, -1.0246609789174, 
    -1.6182038707868, 0.44486222937361, 1.3614755416013, -0.196498331394031, 
    -1.29371304394684, -1.9643664749681, -1.53086103281026, -1.5856097244051, 
    -1.39383562534223, -1.49287539877, -1.94668969651831, -1.70466487019758, 
    -0.952833675705484, -1.37774446573224, -1.19810808432247, 
    -0.339537117141178, -1.50022998005058, -3.98570040969422, 
    -2.02615210855947, -0.313445777057519, -1.23304310284752, 
    -0.942223099121891, 0.707024897654556, 0.955310308666988, 
    0.326562613237744, 0.506379471310492, 0.700624562031193, 
    0.246111182937527, -0.179082315254774, -1.71104242557189, 
    -0.958932070743315, -0.909969416508472, -0.0848159019987623, 
    -1.23265477083108, -1.33553944686815, -1.31294392223115, 
    -1.78727566857407, -2.0695745901367, -0.796761054665724, 
    0.405781445591495, -0.310530245117926, -1.29059576188857, 
    0.607693030620657, 1.94508072719137, 0.756924821088062, 
    -1.96709065485105, -2.21422527996013, -2.58878366869562, 
    -2.81854760050002, -2.09023148753078, -2.21277595835258, 
    -2.17204201403478, -1.34960557289351, -0.549646860241841, 
    -1.12076095469053, -1.55035367144293, -1.57423497042719, 
    -1.72088053994532, -2.79177424525774, -1.08876937212633, 
    0.496126643547985, -0.949766016854644, -0.616780182395649, 
    -1.6035910291161, -2.81182319753896, 0.442532905476503, 
    0.784169554557264, 0.670265461486803, -0.317250765466248, 
    -0.372253866383283, 0.349063011655949, -0.532358160348712, 
    -1.20700078812852, -0.647300924400185, -1.22510083828018, 
    -0.800653337529438, -0.719213824499221, -0.777629066838146, 
    -0.81332245005227, 0.354237518045672, -0.056210105274177, 
    0.081442952377806, -1.34241389616253, 0.223564274397692, 
    0.453201057019399, 0.136457434077784, -2.21108997945598, 
    -2.14412668460033, -1.70613751624495, -1.73535006235481, 
    -2.08710679479424, -2.43950619897781, -1.74491688675516, 
    -1.41833123427713, -0.674406305025204, -0.852782119494186, 
    -1.81027105485136, -2.12731876897664, -1.73813482349357, 
    -2.20238143068291, -1.62337659407937, 0.637620992473331, 
    -0.039644859908492, -0.572199189447267, -2.37790943481158, 
    -2.81182319753896, -0.401903222378488, 0.0974623937030072, 
    -0.0235697562838915, -0.193480103913179, 2.37115328362846, 
    0.657957399356358, 0.0876855060577542, 0.42667126988835, 
    -0.862623805544791, -0.171790095244111, -0.29989152080554, 
    -0.269216282697355, -0.495323190071284, -0.158717880627739, 
    0.336773918045585, 0.388721479716887, 0.483811045517832, 
    0.144223216065016, -1.0632338738337, -1.36611816933292, 
    -1.95406030299144, -1.77972952432939, -1.74472018421894, 
    -1.35342859420474, -1.84560191438384, -2.01864267525874, 
    -0.933349736580116, -1.30462229955308, -1.41089226457458, 
    -1.3950776954827, -2.13015385834338, -1.89133412483956, 
    -1.00393361632392, -0.377427757893285, -0.138207712191987, 
    1.13430801272911, 3.48291140334569, 1.64922042829879, 0.85945868539896, 
    0.6204869995817, -0.39834271570248, -0.259948762078315, 
    -0.659829867280806, -0.484896197107085, -0.509893285570895, 
    -0.126295266427143, 0.401417962818238, -0.645767614339214, 
    -1.58782504545711, -1.54106503716332, -0.634473782277749, 
    -1.85333896349936, -2.06404909236626, -1.57336581795906, 
    -1.71900038621922, -1.31359421452126, -1.4371102370221, -1.8866881892367, 
    -1.5854433752311, -1.73053214335144, -1.27124743572588, 
    -2.18741846218628, -2.26381040781408, -1.77064670704575, 
    -1.27074522507655, -0.456056938004741, -0.681903057522879, 
    -0.987141923429635, -1.01805063999948, -0.914375324753398, 
    -1.11361572456811, -1.98852901073264, -2.88548254103326, 
    -2.79803871642783, -1.30815935351848, -0.655651734909921, 
    -2.22393248954482, -2.21576356753126, -2.00603596069404, 
    -1.55916520726584, -1.57469727337083, -1.43063482675536, 
    -1.95662437883612, -2.00060356907455, -1.301374579724, -1.60743669891426, 
    -1.24219975798173, -1.46123455472555, -0.382721726665687, 
    -0.772723891138547, -1.23417468281245, -1.26485188462124, 
    -1.80497058865047, -1.85260546804516, -1.94614508889895, 
    -1.66211425668816, -2.60647025930977, -2.03523011442694, 
    -1.20856759993247, -1.56698050342455, -2.26229574649354, 
    -1.92934850166492, -2.10642732840944, -2.17357705545436, 
    -1.62935798521441, -1.38893148964018, -2.57031089092172, 
    -2.87482598978551, -2.96493539368584, -1.345238703834, 
    -0.0552846629085561, -1.1401558242136, -1.17155488973373, 
    -1.1398180771225, -2.61643568060482, -2.61028246899446, 
    -2.21904765336033, -1.23227275841661, -2.09871282272862, 
    -1.82810816501639, -1.33290160001381, -2.07514076346023, 
    -1.97839996784741, -2.79283613377381, -2.56012353813919, 
    -2.13000740973912, -1.34663390431551, -1.72595384429288, 
    -3.85219897451621, -3.94437676622354, -2.02379614663522, 
    -1.45873433758203, 1.14072156853383, -1.48501507482526, 
    -1.59331305595761, -0.77296057981056, -1.55295827163307, 
    -2.43394754891766, -2.2145441092048, -1.20815846811783, 
    -2.18940256181997, -1.8836942103774, -1.31163781235402, 
    -1.95972375534204, -2.28226517832931, -2.46110122972337, 
    -2.51115889303419, -2.29213223572479, -1.9638863136929, 
    -2.15061816785158, -3.39952914612048, -3.40721866595097, 
    -2.00037086790434, -1.3163008494008, -1.6582458341908, -1.25171633775299, 
    -0.62354038503956, -0.951545120889499, -2.15202086190749, 
    -1.6011198931202, -2.28829890383134, -1.87808552366312, 
    -1.24737254372548, -1.33207872350554, -1.59248117852993, 
    -2.24543911681728, -1.78784938838476, -1.98932085565063, 
    -2.73697835519558, -2.20710045178775, -1.97572436804933, 
    -0.939326843078887, -1.62429321415128, -1.81649514662447, 
    -2.19174905185118, -1.78299657346815, -1.48368117466235, 
    -2.78352081448571, -2.83214317730117, -2.15921568103156, 
    -1.60767086833455, -0.627141643439528, -0.413073898472156, 
    -0.764540630530632, -1.1107865803967, -1.72879790767197, 
    -2.03414003621306, -2.56397026929008, -1.60332376318985, 
    -1.36906191709682, -1.4320273951301, -1.948424109327, -2.50989780152714, 
    -1.8393667717786, -3.50785153257994, -4.03956027078782, 
    -3.28222758962689, -1.24254679919174, -0.301546841759208, 
    -0.0335379123606128, 0.504961808288886, 0.678451033397569, 
    -0.0758480678600293, -0.117110613594158, -0.615943441863708, 
    -2.12664685094849, -1.29597061261951, -1.30521405533839, 
    -2.69035053272471, -1.47810056071674, -2.95570975575402, 
    -4.23903240739921, -2.9676976538665, -0.751733888731625, 
    -1.01619373442495, -0.540428291750632, 1.26794623545892, 
    0.386154393464766, -0.184088769279915, 0.0918859234308167, 
    -1.98204926132131, -1.01194469367262, -0.343398285467105, 
    -2.42515151680553, -1.70242289160372, -2.27182879329269, 
    -3.84716440367228, -3.076821335228, -2.13091418521124, -1.80504101385962, 
    -0.530890781771385, 0.120793650214992, 0.553234689191715, 
    0.513312810468571, -1.25059770025099, -0.350415686786922, 
    -0.335342160803545, -1.7690031751241, -1.42856413492443, 
    -1.13897537638922, -2.13638850151523, -2.34424111316993, 
    -2.40436898030356, -1.68750722422415, -0.63296642892265, 
    -0.797900286614914, -0.723552533185989, 0.0231730076067382, 
    -0.489794779839405, -0.607884271190273, -0.0806680603998977, 
    1.49930846365409, 0.750356945712363, 0.0830242484437485, 
    -1.49177506097839, -0.632506150502699, -0.0933038441344314, 
    -0.434280600679888, -0.717656025857702, -0.712712752035003, 
    -1.3787187437013, -0.819686473248815, 0.158071592980948, 
    1.05231144230694, 0.350124664538463, 0.534428054909686, 
    -0.207323162977984, 0.244307268389035, -0.370135662639153, 
    0.119168612995981, -0.508715509722331, -1.09682726924244, 
    -1.40127512814321, -0.132218940995381, -0.702872899451115, 
    -1.44241239304574, -0.323726588498103, 0.220140737963539, 
    0.77552806223391, 0.560362463145943, -1.01811404327641, 
    -0.416399083752941, -0.934282326009588, -1.13250353307257, 
    -0.288644118137937, -0.778599612557787, -2.46590632731679, 
    -0.280970083489103, -0.367592400809915, 0.0970179547239525, 
    -0.218017858569723, -1.54228579201507, -0.736581624645387, 
    -0.99117279087217, -1.05558123713094, -1.74709072061395, 
    -2.05640148667163, -2.51788353032701, -1.66901379478296, 
    -1.52183086221691, -1.31477331860058, -1.93836100915279, 
    -2.09161191036371, -1.28598618250203, -1.84552749997561, 
    -1.8826821245933, -2.59604862472014, -1.77588788537894, 
    -1.88160545928802, -2.05570961548389, -2.60052073457212, 
    -2.30097568750238, -1.71539459551683, -0.880611761369847, 
    -1.71269897178979, -1.54851969071024, -1.4343087694599, 
    -2.04793657184811, -2.39783486499, -2.17622255589883, -2.17287612557712, 
    -2.35304635954199, -0.740576389450207, -2.21323187502485, 
    -2.30903888939586, -0.999553042930952, -2.24200326332847, 
    -2.96825399725926, -2.4331969272268, -2.0966703239479, -1.69259054336587, 
    -1.90659990881458, -2.45193702372426, -3.47175226673742, 
    -2.23942223217374, -1.60507945275446, -1.23518262553889, 
    -1.72325892177482, -1.4369889951343, -2.54271359433808, 
    -2.96147147613101, -3.28297170190339, -1.3653610870045, 
    0.0816145625067044, -2.19470036272942, -1.63801730459876, 
    -2.62326426703748, -0.201924417731298, -5.81242609591001, 
    -4.02157229791401, -3.32341523609815, -3.09213971470065, 
    -5.59089083570127, -0.448545724739821, -0.793030323019632, 
    -0.414668451145392, -0.435439976451916, 5.04731541430132, 
    4.8235817337364, 4.56132238870595, 4.73663595257108, 5.57738428804697, 
    3.36561073829228, 19.4449554844084, -0.187002193625411, 
    -2.04161896780595, -1.85205506023488, -0.982102427529803, 
    -0.349994125336757, 0.451998431456371, 1.10076013790817, 
    1.33279474632114, 9.0057056355819, -2.61639237349242, -3.13444542616892, 
    -8.9189467893886, -8.44857696393164, -5.01806325111794, 
    -1.19997236019487, 0.662045758608736, 3.33486417126799, 
    -11.0366152447575, -11.1626945438658, -11.8621381583019, 
    -12.1078372158841, -10.9996814728277, -0.828823234592517, 
    -1.20773416250039, -1.84681150342119, -4.80504294600139, 
    -21.8139000821211, -14.8040495607695, -9.17511320698878, 
    -4.36112777496263, -4.02554046491517, -0.801441055812546, 
    -1.41980716137903, -0.945347198533593, -0.630786781707181, 
    0.0718167023083555, -0.53345478375523, 0.503445288184047, 
    0.398592217331217, -0.235119556801038, 0.872453599609292, 
    -2.15960078025205, -1.20336247731611, -0.268529825582066, 
    -0.872014819371469, -0.982275117220301, -3.35068542478096, 
    -1.44612716537114, 0.55871129901878, 0.145062566914762, 
    -1.52797061116967, -1.34582788033664, 0.591677482662437, 
    -3.30974623090603, 1.11664594783874, 0.158522198694742, 
    -0.574705108583876, -0.369671510814658, -1.61906763748206, 
    0.705230187898934, -0.111598439583827, -1.69812577792521, 
    0.0128563349579391, -1.00512365037197, -0.967165617424863, 
    -0.404194317574386, -0.854945292001664, -1.10635543119082, 
    -0.148956160516349, -1.52438657775102, -1.43421004803318, 
    -0.829718843425795, 0.0179400340865263, -1.05958566312239, 
    -2.03927659055139, -0.602210910611307, -1.93462649085661, 
    -1.23061159978322, -0.518549247596724, -0.545232047180383, 
    -1.09931648027544, -2.68257834485517, -0.496042804261627, 
    2.07751107947197, -1.33287225428627, -0.433995245231366, 
    -0.517310484880765, -2.30247228651369, -1.39354235997349, 
    -1.28823672824546, -0.151457486134418, 1.39554128217568, 
    0.0313661573045479, -0.205127450059631, -0.470694414425595, 
    -3.08373423428528, 1.19705570824633, -1.01499362023814, 
    0.804834975232859, -0.517552184430607, 0.574736024497588, 
    1.22602906175329, -0.840419524634792, 0.245505422184612, 
    -1.2677931069135, 0.710516193379931, 0.155817123408476, 1.15055109411787, 
    -0.873617639159556, -0.145270185019963, 2.06978956218542, 
    -0.019124475410192, -0.903701369751821, 0.615869019464338, 
    1.48989882021212, 0.950302545128613, 1.32178866552688, 
    -0.144175046479919, -0.370067729951513, 0.0710945184936043, 
    2.37381859902792, -0.756213311603862, 0.17418122983263, 
    0.309429541092217, 1.84966732116429, 1.0525689869113, 1.94947327753612, 
    -1.94915741849222, -0.846708716989854, 0.0455535916987701, 
    0.595754228793915, 2.0828903648882, -0.583704125484855, 1.30328899246574, 
    0.0299158670543323, -0.0326634181114963, 0.707331909004227, 
    2.54986381538891, -2.11725342812485, -0.0393913327636289, 
    -0.0483661109750178, 0.387734186192173, 1.4564320164458, 
    -0.262619644367142, 1.84599075548674, 0.0214399211960939, 
    -3.57975142652727, -1.23737866897257, 0.0249304950804358, 
    2.37777028950745, -2.1374611391392, 1.28166502601877, 
    -0.0149737612833697, -0.270142855866366, 0.840487564151, 
    -0.267151647718916, 2.10171149902047, -0.383272368610989, 
    -2.94503519864215, -0.89317335574423, -0.557180236243496, 
    1.40201919422657, -1.9871143246418, 1.91416636298107, -0.428269572027941, 
    -2.43127800996426, -0.765933946716266, 0.141786081265304, 
    -0.874352699919472, 1.86248575228524, -1.11383592606764, 
    -2.67345411106953, 0.381489428876503, -0.444936376355186, 
    0.433565100575985, -1.09085517868008, 1.82451818033284, 
    -1.40223407038688, -1.33806871505031, -1.22319804521434, 
    -0.352510041427016, -1.65316688557887, 0.80622692519898, 
    -0.660112388010552, -2.13396874390777, 1.37274802423669, 
    0.000512843896697396, 0.177595164352071, -0.398190373279492, 
    -0.734708470582987, 1.10918050682736, -2.05481655859399, 
    -0.716118354920332, -1.20091278867453, -0.322070830872671, 
    -1.64624738964693, -0.190671784697929, 0.476495597626712, 
    -0.77777878465987, 1.41968625759284, 0.525817793096728, 
    0.0210517558459078, -0.747407193133334, -1.48947831155387, 
    -0.000526385864965673, -1.21542115805009, 0.266802756229283, 
    -0.781192725313287, -0.187507059020582, 0.565762995528478, 
    -0.307129005957357, -1.06392916801169, 1.14379889326943, 
    -0.164228228955032, 0.546172846180978, 0.282632160616684, 
    -0.854752994133866, -0.558610950516986, -2.04582795001633, 
    -0.725072377942261, 0.0279932057597548, 1.44105211598808, 
    -0.189926282402052, -0.592250605375011, 1.17476174405408, 
    0.634897339338561, -1.09169677387277, 0.978590817824296, 
    -0.837806268261344, -0.461888454550412, 0.698158654555083, 
    -1.21538691373958, -0.0418838704661376, -0.670150674532069, 
    -1.04238827662333, -1.20605724321911, 0.382070215758015, 
    1.31633936397384, 0.0904991424647894, -1.15772553683386, 
    0.661341430615518, 0.131879934093003, -0.676690174479427, 
    0.413177733561362, -1.46956391895344, -1.03688203825409, 
    1.87820373887361, -0.905355387866646, -0.0129179260081311, 
    0.529737322273157, 0.44714007697524, -1.1028831978398, 
    -0.211888145974513, 0.278767847971947, -0.151963640613674, 
    -1.31256090525994, 0.74921218555478, -0.437032293334659, 
    -0.252296997402192, -1.36685244328342, -0.251915855779656, 
    -0.78550439233836, -1.12082765172015, 1.62932880437024, 
    -0.203190613880301, -0.276963939843693, 0.51111801370222, 
    0.655220648017654, -0.981212941755437, -0.913692977135674, 
    -0.179785934764953, -1.07880266566753, -1.24709596960253, 
    1.73924140965262, -0.489885020971625, -0.0267981282384228, 
    -0.032885938244058, -0.543052904748403, 0.567105614119541, 
    -0.920718698200523, 0.024812724448417, 0.0419707907520314, 
    -0.853333827404019, 0.234843003906009, -0.0528426692438466, 
    -0.992380398310858, -0.63722044107027, -1.67542082124696, 
    -0.0354977693590053, -1.88017689219569, -0.947456851176004, 
    1.37951252557445, 0.020809522661662, -0.224872290651412, 
    -0.721660766245181, -0.835166174855578, 0.975033830035552, 
    -1.11589169375621, -0.898066707875462, -0.514134415468587, 
    -1.33274797718406, 0.357510728877734, -0.532268113384858, 
    -0.972469985765568, -0.157406382663455, -1.96922360718204, 
    -0.0514798440574241, -1.73815204918791, -0.583316023550001, 
    -0.504882424882463, 0.433809383624052, -1.06073825943713, 
    -1.88906011701424, -1.44812318730069, 0.209709815202865, 
    -1.51784842201058, 0.334993862724211, -0.643443255603553, 
    -1.27517290460286, -0.807583209610549, 0.2169542094607, 
    -0.204263567067146, -1.2008399936169, -1.86048727193592, 
    -1.92280436866797, -0.466553301445848, -1.33640803741125, 
    -0.626456694562098, -1.55726135668502, 0.429178623685002, 
    -1.92032951751821, -1.98754587798403, -2.05437611027217, 
    -0.547520116587234, -1.52400569552052, -0.191003642592391, 
    -0.45959997282925, -1.39947149471144, 0.431219919063978, 
    -0.704197619359222, 0.485531863265058, -2.21093739091942, 
    -3.11155603244859, -1.92027529079187, -0.828532663371816, 
    -0.89770848850868, 1.20812573660057, -1.02335174196512, -1.105403882886, 
    0.174223294550846, -1.28261534294428, -0.996355066318499, 
    -2.00200086292136, -0.435724669842649, -1.63540318021864, 
    -2.06603232121819, -1.04672382479447, -1.14378023028444, 
    0.814732507051625, -1.30196341846767, 0.658155529659638, 
    -3.30450993419358, -2.58949708092517, -2.06567760002695, 
    -0.838816747585158, -0.258078118325055, 0.229825982246078, 
    -1.01802119443571, -0.6024780437065, 0.16007872457211, 0.654303468956027, 
    -0.364910798263184, -1.68480544034266, 0.267672038628067, 
    -2.66419491088499, -2.91016435349258, -1.46511762010956, 
    -0.747799589089873, 1.78080558288307, 0.0158921108144749, 
    -1.01928570219051, 0.598274831314932, -2.81943523216899, 
    -0.773846343516325, -2.12753166276758, -0.81785892026896, 
    0.0220302980309102, -1.19416761436718, -0.809920448834315, 
    -0.986538961846675, -0.0185948759441698, 1.48975818225486, 
    -0.430573165579, -1.02231180761064, 0.363245540060508, -4.06394738287696, 
    -2.21947690314366, -1.27720093645711, -0.15877043519009, 
    0.273851180810694, -0.837750385023289, -0.569873831139969, 
    1.02350983319692, -0.569558809533111, 0.139882915392344, 
    -2.45131982225313, -0.671373997399502, -0.963792121262409, 
    -1.72653643238774, -0.222359034051491, -1.35017006191908, 
    -0.590978061501097, 0.877694911741468, 0.547295853693961, 
    -0.75053080950726, 0.00689568015230565, -0.0682071655128444, 
    -4.06277102383625, -0.101124145702933, -1.31381929281156, 
    0.353415022875863, -1.00104131408734, -1.00263882548033, 
    -0.51142179469729, 1.01978222105681, 0.922677325723147, 
    -0.102225351095069, -2.48941365057671, -0.830531326604544, 
    -2.91160134647101, -1.34365023525724, 0.31045362095886, 
    -1.46712562703325, -0.749543586899589, -0.573879632278296, 
    -1.51967922240334, -1.22485682419456, 1.19344081519398, 
    0.293280043254115, -2.12219437826501, 0.995992433728947, 
    -1.12610479917733, 0.107710445677628, -1.33087623703137, 
    0.177711429598137, -0.452959701792864, -0.120087543869342, 
    -1.11043099317105, 0.220109193108971, -0.809075863875942, 
    -2.03791324043762, -1.98528757127455, -3.78364331221066, 
    0.30967411609015, 0.145535245268257, -1.80792549026768, 
    -0.218285418519279, -1.8810167021965, -2.90803189356513, 
    -0.903197214607098, 1.74407615573104, 0.663256238116985, 
    -0.347814817753487, 0.60092710361612, -1.20341919291632, 
    -1.19375201326753, -1.05422442062959, 1.6117599322182, 
    -0.984737436065741, -1.01192020827814, -1.75594919823163, 
    -2.22280346251803, -1.95815045614043, -1.5008424629349, 
    -2.09748354355156, -2.24489319413995, 1.74571207256683, 
    -0.0149899108935762, -1.57884370200756, 0.162338286580193, 
    -1.58528048401281, -1.38078901560408, -0.220940403855798, 
    1.71645236346865, -0.399933120710486, -3.38560735347821, 
    -0.0928441653172594, -0.443110682608605, -1.86035105400781, 
    -1.80066393258019, -0.113848486029616, 1.88270339280773, 
    -1.89451590275858, -0.951720397759301, -2.30105625604912, 
    -4.15874009987425, -2.35377627125043, -0.845623194945514, 
    -1.5882055474208, -0.075276002681636, 2.36327826100872, 
    -0.685669836664766, -1.15981356351, -0.371414198451364, 
    -0.558107393467758, 1.214689701182, -0.827136766352988, 1.19554832755781, 
    -1.5316558231184, -2.42253412364202, -1.50661249052669, 
    -2.31688964872631, -0.655816652925934, -0.439801776036869, 
    1.36341157674059, 1.34392906737813, -1.66764393884607, 
    -0.885945511790439, -1.47617643779079, -2.79319737143996, 
    -1.90443431665642, -0.0078250998005177, -2.41483613391753, 
    -3.58628763305101, 0.906868829153129, 2.29353421521109, 
    -1.90832146003406, -0.602273368722921, -0.526777633102408, 
    0.278057717393006, 2.39296174822626, -2.45440842905026, 
    0.0548810500882475, -1.73567332098834, -1.49383828996671, 
    -2.66394996443957, -3.94386373457755, 0.669972303011798, 
    1.28222364775462, 2.69865487547224, -0.500963080496257, 
    -0.648542800223783, -1.26768946653384, -0.104386534704403, 
    0.256235866951811, -1.94733569068448, 0.388926212608167, 
    -2.93138238687613, -2.60618664028895, 1.21751515835453, 
    0.0683746901468094, -2.94340348172779, 1.52280071249564, 
    0.402883215948449, 1.00175675490719, 1.79284158858852, -3.03451623430015, 
    -1.03045164696505, -2.37003496850454, -0.716392124514495, 
    -1.864310922507, -4.1483867411901, -0.370490126568424, -3.02676074435718, 
    1.37370138116231, 3.36959472986127, -2.83290321876037, 0.362342167843682, 
    -1.34581243857171, 0.179379383573167, 1.87615727211375, 
    -2.74654723647668, -0.339405492742491, -2.45932538673513, 
    -1.33967434070716, 1.79008413565255, -3.0305571322609, -2.53507044917318, 
    3.17832045069604, 1.15699548100957, 1.16837450414743, -0.524967267714781, 
    -1.6407313164196, -1.91605621521781, -3.10638874649026, 
    -0.481863305123839, -0.0719425941264382, -3.56920836499679, 
    -1.39166619315188, -2.68113411307792, 1.07681759884039, 2.56076102406469, 
    -4.02262915308334, 2.05960483245008, -1.01975106691561, 
    0.0986153121668368, 1.47522599826979, -3.21582613685109, 
    -1.60247725646461, -2.71109636193214, -0.571810617210836, 
    1.81429816098352, -4.30256984580051, -0.37104496032622, 2.07025922522325, 
    -2.36111468140239, 0.612660206795792, 0.648586563973103, 
    -3.3009451638052, -0.288286296961572, -2.34852734504719, 
    -3.27310013281294, -1.66868071438478, 1.0463336957011, -3.15036129236602, 
    -0.724591353844108, -2.17522543641361, 0.943262761639789, 
    0.244378680788191, -3.30308117149574, 3.48512400812733, 
    -0.466334160384932, -0.178722437026558, -0.194947901037941, 
    -1.83021060264658, -2.877131380304, -3.54208313844469, 
    -0.888800295896039, 1.0204033958201, -4.00292642810441, 2.04795867344475, 
    0.400475270890688, -2.31253216403532, -0.315772845812757, 
    0.711935930186276, -5.0671822169556, -0.029452733468853, 
    -2.10121170782533, -3.1471916070393, -1.85633000523601, 
    0.931385210717704, -2.98935145199532, -0.0408122291283401, 
    -1.44872527903559, 0.61318810163586, -1.76267368175157, 
    -0.819431018960779, 2.97518906606179, -0.96696792014821, 
    -0.440998534899772, -1.17268180690788, -2.31179872076318, 
    -0.278503445004128, -3.65588807178943, -4.25884761262462, 
    -2.82751651055169, 0.104649676141818, -3.47875468630108, 
    2.09284834778357, 0.980180619344909, -1.99948252675746, 
    -1.01140038320352, -0.099029144737969, -5.22869003991181, 
    0.273629426901892, -1.37939215130911, -2.17402069842908, 
    -1.22853009065231, -0.0249708316627406, -1.82008016561436, 
    -0.572020842850768, -1.34323459065225, 0.011229752786851, 
    -2.33252883230332, 1.84851452923055, 1.594532452466, -1.06433072427135, 
    -0.959454884367075, -1.03462429043842, -4.30898533394693, 
    -0.0395015068721002, -3.67694032290719, -4.47496308332037, 
    -4.33746327067385, -0.179737337704994, -3.22082412357909, 
    0.134111458171161, 2.33345039085126, -1.52093204722126, 
    -1.39457183756232, -1.47421915813159, -3.33838116514373, 
    0.638409361014559, -0.937034898008889, -0.247873350259074, 
    -0.975810395411118, -1.48485325565325, -1.02862042586814, 
    -0.632763795025383, -2.20052054809305, -2.70287971689601, 
    -0.721833886867389, -1.93247275766847, 2.36016955486672, 
    1.74786739477825, -1.0954083072824, -1.1305659692716, -0.863392254057475, 
    -5.46526966881754, -0.0524111137058945, -2.75233640187939, 
    -3.14313204642587, -4.07120380833398, -0.235094205973205, 
    -2.45879294362638, -1.39660841092989, 2.2377820504366, -1.35579731938344, 
    -1.41978466828432, -1.83877310244299, -0.893194748823275, 
    0.402902709386991, -0.994174780442899, -0.135376135910418, 
    -0.389920617412581, -1.52633198494628, -2.26372973044992, 
    -0.324410511501224, -3.83541366364809, -3.92448236918169, 
    -0.747722857002293, -1.55692805317392, 0.816938202423978, 
    2.98859251493497, -1.08965917414887, -1.11374416415522, 
    -1.88391220909416, -4.79892103224257, 0.293200817742195, 
    -1.53963996259505, -1.55971677258997, -0.985506387972017, 
    -3.8165535118596, 0.088026012020017, -1.7516093828195, -1.65948381035935, 
    0.220603275257363, -1.94418168472423, -1.83341721308829, 
    -1.26197216895333, 0.228183229791111, -0.202349648714897, 
    -1.67555439882074, -0.634655384999889, 0.00150742737968015, 
    -1.2429612599528, -3.90568376162425, -0.193040390598888, 
    -3.46982292980818, -3.41900771446052, -0.288184633442529, 
    -1.43615077614008, -0.278050345874872, 3.19774262950611, 
    -0.957952802116005, -1.47064094482012, -2.27988727522624, 
    -3.4618066437528, 0.365428929742138, -1.64140517331228, 
    -1.65698159854086, 0.229619254230114, -3.72768622252553, 
    0.465556731724421, -1.3572319774801, -1.68156427378949, 
    -2.54897741221771, -2.50638952488308, -1.98777630954787, 
    -1.14848500124008, -0.341532224809673, -0.159107543136221, 
    -2.02626219960606, -0.146424098633628, 0.295221139305867, 
    -1.4523611001054, -4.64889297508078, 0.31718395105207, -1.6975295680229, 
    -1.32585062363817, -2.25607288035677, 0.147446794532767, 
    -1.56970407569682, -0.130374171395098, 1.35703928044355, 
    -1.27654859504967, -2.65037351231771, -1.56896130863451, 
    -2.34992310995135, -0.615248259208313, -2.70471213702398, 
    -1.68887416997713, 0.45587884155654, -2.36326834693595, 
    -0.17594659601945, -0.903941165254755, -1.49262891962239, 
    -3.53243465343236, -1.97171984954866, -1.22817404120573, 
    -1.46516322093179, 0.0175580931644529, -0.021144139039371, 
    -1.70788170800668, -0.296327312150021, -1.90330212436572, 
    -4.23070430380171, 0.787425130448065, -1.27150870374872, 
    -0.299442694793606, -2.23235745715393, 0.518118709767187, 
    -0.976049124873728, -0.379550072707656, -1.42724150441851, 
    -2.25066445728618, -3.17419420210508, -1.23781537585881, 
    -1.82248747455431, -1.50832178059297, -3.29431019114212, 
    -1.64697348133128, -0.320703308583195, -1.51243381569545, 
    -1.93002542661699, -0.429228497954687, -1.72759265410537, 
    -0.925832655764159, -2.30954589692761, -0.927096384141193, 
    0.0603038744159547, -1.5952437706385, 0.29454860026129, 
    -1.11709848451752, -1.90512123930674, -1.56833728055142, 
    -1.80138373324685, -3.39574075683388, -0.0720936166779595, 
    -1.77899054919314, -0.566582635256805, -1.87499210100554, 
    -0.417963088826002, -0.385370251390438, -0.687444389420552, 
    -2.80745992299032, -2.93907146965919, -2.31625998968159, 
    -1.29399003896478, -0.860065841337666, -1.25686653335313, 
    -2.92411152095216, -1.22921266878121, -1.92966670313868, 
    -2.30943992966817, -0.0620137076610051, -1.37303112642212, 
    -0.6798696360332, -1.59238735170356, -0.680126846287107, 
    -0.0428383613355475, -0.852179014725437, -0.435550083992736, 
    -1.93173509859587, -3.13510000342351, -2.3032548365984, 
    -1.34436047365337, -2.68318490292914, -1.42183488639112, 
    -2.75781875018791, -1.20315600951501, -1.70254568990851, 
    -1.95776083171899, -0.455443896474001, -1.89991443697047, 
    -0.818614170851758, -2.38008490399725, -2.58364482358603, 
    -1.13621949466292, -1.15356075008426, -0.246317082523297, 
    -1.56214178241268, -2.77189026871712, -1.07989630456348, 
    -2.71576017303369, -2.37784740390093, -0.529536138170007, 
    -1.54935334029391, 0.579661162087237, -1.71604299338729, 
    -0.941785134496493, -0.663851852117858, -0.203931792063594, 
    -1.43343772360831, -1.65061750160009, -4.22586924434808, 
    -2.36419261532508, -0.313181564301971, -1.59091099571082, 
    -1.28512487312241, -3.22078985278726, -1.82801321476327, 
    -2.57147990201807, -2.05126375413034, -1.12209216319555, 
    -1.99851298316591, -0.930497171447278, -2.22556856664154, 
    -1.32589397995117, -0.628643371526058, -0.546996100362935, 
    -1.02875195481132, -1.78193765071123, -3.55881862674223, 
    -0.46970745194083, -2.18435616508889, -3.04700611729286, 
    -1.35844590182899, -2.29927610375816, -1.42910335615007, 
    -1.69534700713667, -1.75855160121818, 0.0701497451770103, 
    -1.5769282611271, -2.19471424627873, -1.06002863247531, 
    -3.75746936402222, -1.63372859938459, -0.0886651551370173, 
    -0.866559188999251, -0.643548092065505, -3.16866399819029, 
    -2.10789923042536, -3.46857602851781, -1.92349849637429, 
    -1.50030414105054, -1.89435649254601, -2.4337844631159, 
    -0.807673419984188, -0.618206884900853, -0.136035700900575, 
    -1.54733784732968, -4.35043427302761, -0.0546679246369544, 
    -0.465063378879042, -3.2243149470919, -1.45740659202469, 
    -2.80004486539315, -1.19359897359074, -2.9683512213834, -1.8821263310106, 
    0.0497182602424704, -1.82525631358528, -1.93528900535685, 
    -1.48420561688013, -1.79087597245483, -0.641169400824774, 
    -0.186367195325107, -1.97801280722148, -0.309359692482308, 
    -2.86021475451915, -0.626145711717421, -2.21183638919487, 
    -1.31741021880761, -2.31667260548622, -1.23358502690408, 
    -1.70578358730481, 0.336064836454936, -1.40448301071627, 
    -1.20215907089718, -3.86072738449997, 0.042591785426864, 
    -0.19225203870461, -3.097609412425, -0.46703224966641, -2.76668135984053, 
    -1.42959307924764, -3.43642800179354, -1.72703806621333, 
    -0.113259942264376, -2.10532648718068, -2.07549154546084, 
    -0.675371780018518, 0.112174434142156, -0.301608726839331, 
    -0.352707183084378, -2.26156237734913, 0.443408238245796, 
    0.311785466379595, -1.33178222709391, -2.64757319169367, 
    -0.627604421240157, -2.3861509803935, 0.949519802153586, 
    -0.917609862412149, -1.57201156253756, -2.11236655309854, 
    0.73143566206654, -1.72308005113855, -2.96712450912602, 
    0.698744222487523, -2.26608095577694, 0.0453951499972904, 
    -1.08723563740776, -0.616951928777546, -2.86865555954285, 
    -1.9871758212649, -1.23198987170216, -0.0426979638678941, 
    -1.59202951025395, -0.849179020799107, -2.0384241442223, 
    1.35383476331414, 0.372532802759021, -1.16485405234294, 
    -2.42026163989037, -0.713284752030874, -1.7881688205009, 
    1.02251552935365, -1.4305253032263, -2.12159705923559, -1.18821324555837, 
    -2.05274171608966, 0.957240643744637, -1.62439323844321, 
    1.66272922656205, 1.95271441784862, -1.02590444735246, -3.29209453235342, 
    -2.02809798994846, -1.35349600310736, 0.431854181449996, 
    -0.275325157420876, -1.73425623474151, -2.35407170303324, 
    -1.36206734946192, 0.340953383701019, -1.85868007607853, 
    0.659163773434046, -0.374326417986438, 0.119780906088988, 
    -2.50141802942273, -2.08489966172792, -1.48328678692248, 
    -0.438327064871238, -1.45503015818914, -0.091965435967338, 
    -1.54301652396925, 1.72315182914627, -0.948150166254774, 
    -2.33511301344465, -0.858183379894096, -0.59167827946886, 
    0.639406499110166, -0.535426889334825, -2.84239041371001, 
    -2.77442787464832, -1.44033004326228, 1.56214296805605, 
    -1.46172403284955, 0.109216017126446, -0.611435670348453, 
    -3.11481044426849, -2.10929301623842, -1.26932473521283, 
    0.553866416313525, 0.788454051601646, -1.81123063647397, 
    -1.71875844771804, 0.00342401653588981, -0.167050601663248, 
    -0.649677279245477, 0.881233559658374, -0.531340795432135, 
    -0.497736681335252, -1.72002703992886, -2.81645308757261, 
    -2.61481287188871, 0.00297520170277343, -0.557899634727981, 
    0.987290653809811, -1.41204637090047, -0.642709722557737, 
    -0.584716778985874, -2.05508993669022, -0.435840204017464, 
    -0.690672405603151, -0.644094931133207, 0.819319449167319, 
    -3.29488962094813, -1.77379174603864, 0.00997477576819977, 
    0.273086337101371, 0.0666730238904678, -1.71079059720761, 
    -0.936403752586216, -2.34531616755034, -2.255088724057, 
    -1.73637946614907, 0.400657567587841, 1.08985889692963, 
    -0.581153426547974, -0.960249414179951, -1.61909776581355, 
    -0.38786762448987, -0.0036604532544688, -1.2002009881696, 
    -2.59847018058199, -0.456471533790478, -2.81820090646589, 
    -1.89716551818248, 1.00815873215992, 0.352999923130497, 
    0.210036726253163, -0.531363947221796, -2.2909672517635, 
    -0.201221377452437, -1.41828146871538, -1.24868532207409, 
    -1.20013577758447, 0.663222361533345, -2.57028728770503, 
    -0.295178598791597, -1.23529441131386, -0.493581576688421, 
    0.950687690412935, -2.87947848883768, -3.18029894475052, 
    -0.804987406643984, -1.39943328447394, -1.9690180292748, 
    0.554459615187476, 1.40896942516329, -0.653401688967193, 
    -0.994449606649431, -2.13684209985172, -0.162603415920604, 
    0.593108257590389, -1.86802128952968, -3.18550076614505, 
    -0.561387411381405, -0.614555340934274, -0.572018529897254, 
    0.43780951889237, -1.14546903692243, 0.255297004738648, 
    -3.66420935818551, -2.07472790904336, 0.142241525104263, 
    -1.89082831379771, -1.50443700551746, 1.24857564387656, 
    -0.649314542101295, -1.88905230336708, -0.750176868029419, 
    1.62564841354706, -2.8871116284994, -3.72149680234679, -0.55266508692889, 
    -1.65682615888965, -1.41478875864303, 1.58956985522924, 
    -1.71695255957415, -0.769163461347169, -3.13501665075, 
    -0.637926933721236, 1.35017513433292, -2.02180845833786, 
    -3.37528146016308, 1.20276566381504, -0.184241387072181, 
    -2.07776203283231, 1.22892846960699, -0.883496248608212, 
    1.22068284558463, -3.15739726637691, -2.67252184879103, 
    0.385152689518612, -2.16779803620272, -2.36215126498514, 
    1.75773910108254, -0.951817538315203, -2.58416622541754, 
    -0.471323050789599, 1.63679508184445, -2.40759010597062, 
    -3.32247245395689, 1.24332655159031, -0.154175773382644, 
    -2.47086110251706, 2.48573666132463, 0.494732368389039, 
    -1.71727192134767, -0.977956894243632, 1.21883690088376, 
    -1.77223477781338, -2.25947204152711, 1.99022382673892, 
    -0.578678004303332, -3.04650478703427, 2.43378634698859, 
    0.49475988076535, 0.549027340687213, -2.33745800463993, 
    -2.75239647109822, 1.09956874112329, -0.301575932956257, 
    -1.88191082737041, 2.60530466010373, -0.0934679912443365, 
    -0.163759293312933, 0.938305526220872, 1.20083298015654, 
    -1.45201317223908, -0.836328951922322, 1.98745341284692, 
    -0.376039329233328, -3.18210556324884, 3.83455261552685, 
    -0.662767443150541, -0.550143401484422, -0.569414942986262, 
    0.695896394111791, 0.235727644134314, -0.315101508017163, 
    2.20845311918272, -0.490373558439094, -0.680095158485436, 
    1.46443058681273, 2.2891377814732, -0.257574229727237, -1.39758201886746, 
    0.0373013398320292, 1.57552090030681, -0.255513142073945, 
    -1.51834404564575, 3.3476631760529, -1.27820205947662, 1.50763576175298, 
    1.85284886943441, -0.227533524015618, 0.58125708073991, 
    0.884741181619653, 1.79826743019442, -0.88079728188792, 
    -1.76511268464911, 2.56090464094426, -1.72907266698972, 
    -0.199367987642445, 1.49658997596335, 0.66881360232432, 
    0.408211090475478, 0.724793284022543, 1.39347988255543, 
    -1.45221307648387, 0.868803456120699, -0.292731382573886, 
    -1.76359166713985, -0.393844613680686, 1.0673950267927, 1.41214770135698, 
    -1.02579159095923, -1.41683995588829, 2.38544222170949, 
    -2.04391197697848, 1.70732939500965, -0.739944264114876, 
    0.558376386787012, 1.19009716045323, 0.0212189511806675, 
    -1.58391401612172, -0.978810350109602, 0.493497150070361, 
    -3.13942678246991, -1.50478956310847, 1.26681162992852, 
    0.494164097316788, -0.434428165468179, -0.666993610908852, 
    0.662134506584577, -1.76105348423301, 1.07840734149033, 
    -0.37331683862713, -1.97092826966133, -0.870125382108963, 
    0.561269145902549, 0.0929048397063668, -1.67991507399174, 
    -1.53302723179882, 1.31366392998666, -2.95952228021802, 
    -1.40480124190567, 2.21660788145358, -0.760625460577309, 
    -0.153971572323054, -1.65260717540469, -0.613133161188473, 
    -1.54190879946835, -0.801734197197082, 0.025962870440209, 
    -2.64523544233777, -2.73932935270671, 0.0244779495493085, 
    0.306073684753963, -1.65981025942748, -1.12910335399114, 
    0.924417550317727, -1.58277924664632, -1.63682658170037, 
    -0.788472464784942, -1.41055234511493, -1.23726191719084, 
    -2.06868878054208, -0.234179281892047, -1.56775751714423, 
    -1.71725790482918, 0.907491157734924, -2.08418477502286, 
    -3.51393334294018, 0.698549818428812, 0.0347166073839363, 
    -1.29333288753725, -1.96778295806951, 0.288211824093769, 
    -0.438120408452766, -1.27400998531436, -1.80615811647785, 
    -1.34779279374366, -2.88798374306438, 0.177052738771001, 
    -1.76031760632701, -0.928879292745158, 0.558509343145766, 
    -0.692842764077243, -3.43654804894354, -1.09911036806597, 
    -0.142700527702185, -1.21063124040312, -2.37655033602907, 
    0.0834852708786683, -0.0144463225490256, -0.71170518237537, 
    -1.03426755624074, -0.864410087888937, -3.73131020788826, 
    -0.122809874569367, -1.69891735328859, -1.11724202607488, 
    -0.318519514136813, 0.221555120107621, -2.22911744824676, 
    -3.50225108811066, -0.0912606086567732, -1.30785907994815, 
    -0.133208697247832, 0.0328774364880095, 0.15244113675258, 
    -0.983538257443754, -0.366221737636531, -3.35537520309196, 
    -0.802771505468937, -0.641770237473907, -1.61874922247829, 
    -0.772899842258547, -0.994046153020075, 0.630555236869474, 
    -0.799849075561002, -4.06000122474407, -0.197454632675751, 
    -1.62963444426059, -0.844626249527069, -0.119037264869097, 
    -0.280232238016344, -2.27913976792685, -0.45911152099909, 
    -2.02617449308026, -3.2663547782836, -1.00879831161863, 
    -1.28463974732797, -0.982493115448323, 0.803953716696724, 
    -0.0923521197144658, -3.80976475557336, -0.764124457347805, 
    -1.26073931982987, -1.85017135505824, -0.46939709355491, 
    -0.576092067780094, -3.23052437048626, -0.422529673953997, 
    -0.774779056851271, -4.40958103878749, -0.999348322769603, 
    -1.24079833069049, -1.05208542795737, 0.611151742473706, 
    -0.976271428547868, -4.2209886753261, -1.33827187220091, 
    -0.310838826989308, -2.29575403175575, -1.25638876091122, 
    0.262664538195653, -2.83223601024313, 0.0815211629307193, 
    -0.824730297415988, -4.10610612042259, -0.835471973008012, 
    -1.32274426639594, -1.55468289978024, 0.0967950037933596, 
    -2.52229029526472, -4.36689493117315, -1.12108976936922, 
    0.563062082918762, -1.82319625540722, -1.46300349353349, 
    -1.95277801685504, 0.435282210779296, -2.33151136866143, 
    -4.14397617129742, -0.755852270807461, -0.882291079330925, 
    -1.74632565162032, -1.06172696831473, -1.05710659340471, 
    -3.63393422833901, -0.447816199583408, 0.619161323399845, 
    -0.827473829600196, -1.16820587147802, -1.54123989927974, 
    0.130092105669952, -4.73895204908567, -4.16111795791626, 
    -0.478214722004571, -0.200092011941105, -1.51512894247762, 
    -1.12044733901215, -2.7398251921718, -0.183485888708196, 
    -0.734612294868432, 0.0756112658430022, -1.48565479756675, 
    -1.38456548121185, -0.765156538772585, -3.2744456171915, 
    -3.58409850318321, -0.137284273427858, 0.718260648914269, 
    -0.949986318642091, -0.50349848369448, -2.37350075578534, 
    -0.471779262754501, -3.00473390838594, 0.619822773694442, 
    -1.67255877068658, -1.61283175808833, -0.571571815173279, 
    -2.84002269904879, -0.422724680045568, 0.691019325755137, 
    -0.251533192997648, -1.06236837579148, -2.16221665292154, 
    -1.05999060824075, -1.93965019391714, 0.242985330580277, 
    -1.2297285106527, -2.01320899861121, 0.0552815967616513, 
    -2.4694087539085, -1.00643418511793, -0.272946135707283, 
    0.198870803232864, -1.61655052458545, -2.34495239360569, 
    -0.795298039569408, -0.828063758708958, -0.467926618403714, 
    -2.02247373360032, -0.765110738935971, -2.38943909373079, 
    -1.69330154739948, 0.753865160515552, -0.305381045662987, 
    -1.38690068067415, -3.01305496589518, -0.634339179707914, 
    -1.74540654846969, -0.235147092063801, -2.07066341338562, 
    -1.29740713833216, -1.77598403459927, -1.36437313561761, 
    4.04356809131269, -1.08426546942589, -0.551929416156758, 
    -3.29758419106273, -1.49266458499764, -2.31831863982754, 
    0.150364249786481, -2.6129540063417, -0.862328808776344, 
    -1.8387631419389, -1.18524234655374, -1.46461072964831, 
    -0.177435366264608, -4.00566074805969, -2.29513521863333, 
    -2.02187204756914, 2.57709905615756, -2.20768393892932, 
    0.172856535374781, -2.88622973744221, -1.75469436922222, 
    -1.58979546787126, -0.223863531399489, -4.37126955555025, 
    -2.41077073535027, -1.7466086150253, -1.26438803777872, 
    0.762214796353854, -4.42535703622188, -2.52585823353635, 
    -1.30373547307519, 1.7735469125505, -3.39587669807236, -1.59429291383045, 
    -1.1798886199303, -0.866981450563242, 0.408904458611145, 
    -4.50616755901967, -2.89452937727045, -1.16642543244946, 
    -1.95613101421256, -0.402944265977139, -0.532891934720996, 
    -0.658924956916966, 1.85190092041122, -2.89183081767836, 
    -2.50752418783209, -0.503332346320161, -1.18110588575401, 
    0.68702045749357, -0.21946453638018, -0.817842904101733, 
    -1.61731264345078, -1.55571701980413, 0.527204845810478, 
    -0.83145212437772, 2.96753157524781, 0.383509632422001, 
    -0.55429844751492, -1.48041849327292, 0.150018404492575, 
    0.703338657259517, -0.711502412667067, 0.876442825885933, 
    0.206710752768062, -1.45295455040465, 2.96762948738678, 1.23569777365766, 
    -1.09004161361968, 1.48167267560471, 0.140502613746042, 
    -1.21373001420339, 5.20025866121111, 1.89958891053138, -1.29746019081608, 
    2.98479194124444, 0.766646272267045, -1.61455509671514, 2.46066515023738, 
    -0.611907166994381, 5.78723540153079, 1.20163741486258, 
    -1.88271848389783, 3.95919160098665, 0.364595316894506, 1.94597121675894, 
    -0.446485755776342, 6.60187978198992, 0.646769077620851, 
    4.18025753856767, 1.05559972829607, 0.775599385912471, 1.48286935463306, 
    2.99947753091509, 0.895203854974942, 5.95472633368029, 2.48348275187945 ;

 misfit_final = -0.287175043125849, -0.500655712857547, -1.188292728781, 
    -1.22008858893034, 0.739995810529539, 0.433400478731816, 
    0.390879661504826, -0.353370903367507, -0.635422137192201, 
    0.155947216855763, 0.217177610644761, 0.0350171434937074, 
    0.222721001072523, 0.0506249018675353, -1.90844817248254, 
    0.0496995292673086, 0.653020639715192, 0.685881324494386, 
    1.42749212047843, -0.124884845580522, 0.0993573971156847, 
    0.217515931173971, -0.173302343270345, -0.843914067799965, 
    -0.203618141994775, 0.161433263824922, 0.10719481286924, 
    1.30779828688122, 0.484078997626729, -0.832224465541, 1.76101618868901, 
    2.89002291992905, 2.0027008185647, 0.2245891574134, 0.378251133511478, 
    0.774460334742391, 0.455675487737177, 0.486266124769172, 
    0.834887247276326, -0.309940963178668, -0.93803481291717, 
    -0.511314222684351, -1.57469188771736, -1.00168860730933, 
    -0.657259944288211, -0.54030927820452, -0.893068233974668, 
    -0.0238211519044729, -0.335669852092093, 0.0782615547374776, 
    -0.407011554073295, -0.437170860617417, -0.161171941408433, 
    -0.469235660666252, -0.327937220716423, 0.33469449788722, 
    0.690608335214309, 0.637106679852346, -0.380756200817629, 
    -0.586264853088156, 0.336332353516218, 0.243495475157376, 
    0.0251642878520553, -0.191613548169585, -0.0958624385270568, 
    -1.40920834558038, -0.52380612202223, 0.2687467794301, 0.499674311657201, 
    0.673850617925651, -0.260613888896839, -0.183106472036889, 
    -0.0475011099961842, -0.763348516938573, -1.4660895066171, 
    -0.423784316914895, 0.0173582951352769, 0.422808895890441, 
    0.56503008534794, -0.112617051387196, 0.463578763795289, 
    0.526341185759858, 1.11282690137725, -0.0225096716108553, 
    -0.761279093125364, -0.0427533286720072, -0.0314140557845688, 
    0.251826053285145, 0.0203620054231912, 0.264380226751388, 
    -0.321061041627635, -0.659319354851231, -0.86910352655138, 
    -1.40826249564828, -1.36613100767985, -0.778149032018924, 
    -0.755357819653848, -0.106271304950427, -0.363663523927089, 
    0.319631134253306, -0.352769459598981, -0.755758130911923, 
    -0.231368377472334, -0.0331786561632974, 0.0938662579033434, 
    -0.660970181296312, -0.518645232812274, 0.478772378785521, 
    0.521989214794409, -0.634379800905798, -0.737720613497146, 
    0.265668183843148, -0.0470014129876439, 0.1854243999784, 
    -0.718135730252722, -0.880466538564284, -0.857034387340643, 
    -0.0716956117374234, 0.355403189672074, 0.312609559170993, 
    -0.993300765413876, -0.425030916460227, -1.23782342132705, 
    -1.25020493110464, -0.8335585657764, -0.981737436752113, 
    -0.0482822317033804, 0.392395924540598, 0.405041711282061, 
    0.46159808971722, -0.339420302778914, -0.5242259992256, 
    -0.113693175404732, 0.240814046695599, -0.479576796811387, 
    -0.708871172588421, -0.0148944135829954, -0.316118075791305, 
    -0.204966442171046, -0.0524375221205586, 0.163779559956536, 
    -1.67599646287627, -1.89382595224206, -1.28126755003725, 
    -1.24063103722185, -2.26318486977712, -1.55173834676967, 
    -0.15614699951966, -0.034887492562401, 0.5293587908923, 
    0.0514598363321417, -0.866302733472994, -1.43459520364004, 
    -0.780676404077614, -0.435633777433004, -0.575247601002218, 
    -1.09794636104106, -0.685349121134351, -0.141223802051496, 
    0.293536524717313, -0.196323773157507, -0.3770157829869, 
    0.0494576216403786, -0.062620118537744, 0.0965007804584683, 
    -0.396784784219095, -0.582444498911232, -0.108242252259232, 
    -0.60807318676027, 0.371107192351356, -0.180204588562018, 
    0.081938782467682, 0.767689573870456, -0.359735292573746, 
    -0.765298240727668, -0.101499120032043, 0.404898157813074, 
    -0.0671404069346515, 0.951037172633922, 1.36416234625869, 
    0.789244756857368, 0.0783274791695021, 0.313328305816469, 
    0.802349144125123, 1.11088150109275, 0.175768924285897, 
    -0.874110091944691, 0.275339121146865, -0.608569711798319, 
    0.299394394222583, -0.110148340685021, -0.121425488731264, 
    -1.12217683217279, -2.25696797993985, -1.63041177279247, 
    -2.69352548522757, -2.7535189987913, -2.06458726171747, 
    -1.14300593038572, -0.111995928134108, -0.135775438790247, 
    -0.292974747482004, -1.51913317537007, -2.74699689055711, 
    -1.10478068998231, -0.724243969563956, -0.367949182440244, 
    0.00162763890656059, 0.348999707437683, -0.203874635163679, 
    0.676500001668652, -0.0365628948851704, -0.197517964040275, 
    -0.425725328111177, -0.277707151352216, 0.0523803576044735, 
    -0.00935928542085129, 0.0572390192928784, -0.0173439309249002, 
    -0.596454246522997, 0.0728920192768445, -0.58588476438326, 
    -0.847400244254941, 0.13802639983775, -0.0835058240146402, 
    -0.471600182691856, -0.23072737884497, 0.294022280794297, 
    0.914903343977622, 1.28228602149755, 1.61404191931057, 
    -0.731711193794209, -0.875827007346874, 0.306338212901207, 
    1.49358969099689, 1.78133440156332, 0.714617789240735, 0.386956314861089, 
    -0.376598009620168, -0.102545315022167, 1.08113117774403, 
    1.03696579882775, 0.800910753187547, -1.17044418056425, 
    -2.18189486939862, -1.82438099071697, -2.46132631456117, 
    -1.49722027265668, -0.712071635948903, -0.358033566023561, 
    0.132414632809557, -0.209240946993807, -0.0287540091742677, 
    -1.29719774565347, -2.66591244364048, -0.204230496752498, 
    -0.198541647099759, 0.305227391689664, 0.350296979771834, 
    0.660839089532272, -0.303068293723934, 0.108926627374331, 
    -0.247836039177241, -0.421123029392723, -0.771509026850845, 
    -0.386865191225221, 0.0240060867606751, 0.324627176851671, 
    0.731437328220461, 0.0606043288034686, -0.259597478391034, 
    -0.328310289266098, -0.34327153258908, -0.849169578391122, 
    0.404657995749758, -0.0152314417853994, 0.0238685601490696, 
    -0.0746754779047443, 0.139198167456018, 0.932271281341248, 
    1.57539174530632, 0.953565097997284, -0.968103868599508, 
    -0.805265045647094, -0.0386432286806793, 0.802805863613023, 
    0.401168277263162, 0.660526431517128, -0.492642339082288, 
    -0.938116270416285, -0.805114949625407, 0.0953364860619432, 
    0.753460355321551, 1.00266745485107, -0.849727594566985, 
    -1.3419796587278, -1.59129851863592, -0.735793290765634, 
    -0.691708709737875, -0.314183230662279, -0.0741332601546363, 
    -0.0583137587963778, -0.229235590926473, -0.577295793490769, 
    -0.676143071373896, -2.20260661300058, 0.38588040567233, 
    -0.381925381115487, -0.24247867451356, 0.434220236195131, 
    0.542181099882635, -0.506274375159723, -0.0536187146928402, 
    0.0147953063844408, -0.199586241030989, -0.380918242650505, 
    -0.121297405501037, -0.0587879306029215, 0.755207975016279, 
    0.562652631964258, -0.90751777417704, -1.96482494305777, 
    -0.355456294118542, -0.606855999793097, -0.485335550970341, 
    -0.449316703010485, -0.28289591491204, 0.263977578640757, 
    -0.299725334677849, 0.409575825096091, 0.908450809013535, 
    0.510648144404962, 0.502381289344531, -0.457388931206846, 
    0.341815609642087, -0.00550599781871774, 0.227000435056715, 
    -0.682323711964923, -0.0838770805689526, -0.569779143146021, 
    -0.646950310637542, -0.129947281412117, 0.154108604659302, 
    0.0855404735367626, 0.646434214528453, -0.585484465651116, 
    -0.889799528560822, -0.881322380297873, -0.337557513803475, 
    -1.09571470368422, -0.507996963078652, -0.47457792433828, 
    -0.554972940207135, -0.619447903340644, -0.759322326408052, 
    0.694307267919933, -0.00715723222446601, -0.238928894693391, 
    -0.0590245535098255, -0.135681961879204, 0.842325087336988, 
    0.198599776116417, -0.107028794548878, -0.0296071398990705, 
    0.2560349256109, 0.403688955291757, -0.0254862016431501, 
    -0.492926061171537, -0.22384943441236, 0.232615292495901, 
    0.26188835106459, -0.252557995201452, -1.43628187158366, 
    -0.10748909395665, -0.300905094801291, -0.963670303152551, 
    -0.857184492991765, -0.279363655411333, 0.564724222745325, 
    0.561772818185933, 1.36627409072356, 0.630719615345794, 
    0.537764496615036, 0.410167567793356, 0.0263797049043735, 
    0.484856309479045, 0.697225619059076, 0.432440057772903, 
    0.174267514412918, -0.341561884205852, -0.602762814817179, 
    -0.311114150223704, 0.139557866771116, 0.0931065100953088, 
    0.410207686324622, 1.08724814004405, -0.290638083097479, 
    -0.856987961721987, -1.28557892706353, -1.14802395469253, 
    -0.629890837907778, -0.761551529749993, -0.347410422189225, 
    -0.506524690057804, -0.236982780423158, 0.511565554429137, 
    0.5430511607499, -0.988621511798491, -0.0820197546313928, 
    -0.360628739390485, -0.15355197982414, 0.161388946274643, 
    0.276551348970031, 0.138730036016064, 0.404464004742984, 
    0.505338211000739, 0.274749570986499, -0.803410240088929, 
    -1.16242185947224, 0.130764826997725, -0.353577449509963, 
    -0.295942149510253, 0.0512204999681831, 0.160456492611896, 
    0.280650436896717, 0.0639210707989113, -1.09584348825507, 
    -0.816880994789284, 0.193663681236074, 0.7919127659276, 
    0.982174612758091, 1.0314830233448, 0.468084048798065, 0.744531829137726, 
    0.461439319767694, 0.7417449256533, 0.413364644848957, 0.492449517117, 
    0.576475866791819, 0.604950281773555, 0.248316037188046, 
    -0.116288116866672, 0.280019177092274, -0.767655203587956, 
    0.0976963695523692, 0.544135936452577, 1.09967487047527, 
    0.44953621439368, -0.722874308486636, -1.86322441252529, 
    -1.16875866952894, -0.574191755854554, -0.701528687269373, 
    -0.24121175665301, -0.557769453814005, 0.489874371066401, 
    1.66609962504093, -0.215229402279464, -1.49114763869746, 
    -0.651222832273275, 0.176488719320824, 0.229674033276757, 
    0.760497714948682, 1.21766394617419, 1.19016909967966, 0.195004691120966, 
    -0.257121460488072, -0.637997443626173, -1.31944629594934, 
    -0.726140383632461, -1.16420056685254, -1.36580864493719, 
    -2.21918505977258, -1.69463939149899, -0.174657680035865, 
    -0.264726695565312, 0.373819514044924, -0.634916894986257, 
    -0.782346273627987, 0.200485217597111, 0.892215985881206, 
    1.14853625839855, 1.15075973739005, 0.203598816197839, 0.768815112262575, 
    0.589166530576306, 0.88028366551026, 0.706781710270867, 
    0.106567757121843, 0.516988036450305, 0.814603731923254, 
    0.332854327738961, 0.750675262472691, 0.769314756329234, 
    -0.138744664261794, 0.246192933314808, 0.67251827281726, 
    -0.517505645665897, -0.292987956944679, -1.51845331872226, 
    -0.86014988179921, -0.540446851891856, -0.835263038282537, 
    -0.00499560414706668, -0.0194188481618474, -0.549598612085931, 
    0.0825304767422841, 0.769679901790305, -1.62902428978168, 
    -1.54700618085116, -0.966353914260916, -0.238069273543893, 
    0.11960675374648, 0.467526128260438, 0.291155904332294, 1.18268350335287, 
    0.0956497443977256, 0.00412070086887262, -0.368922649385111, 
    -0.756279189853704, -0.280137962018703, -1.26243138624853, 
    -1.2577490295389, -1.47068677571438, -2.10521686479917, 
    -0.391913230481795, -0.97344760923407, 0.284072387813792, 
    0.352015614730377, 0.00244584026031447, 0.484255989810758, 
    0.309064147691207, 0.334205139004378, 0.220002715373631, 
    -0.154477165652054, 0.863869909071697, 0.567454364759641, 
    1.05517673424054, 1.47609922067445, 0.0619717868939862, 
    0.0542959490181305, -0.65735906143312, -0.623947821353914, 
    -0.385571952013648, -0.301359332653908, -0.604559028961527, 
    0.892187291972579, 0.987160512045051, -0.365584656098794, 
    -0.430138937580304, -0.577622620967801, -0.280862736587308, 
    -0.874360390067741, -0.869755730244517, -0.689624000165741, 
    -1.23044635173351, -0.238519936455246, -0.300872401040788, 
    -0.405173150565257, -1.85144232354925, -1.38826870219782, 
    -0.532466045981961, -0.163994060374408, 0.312415626961089, 
    0.166770311760445, 0.306387403136492, 0.202937720822156, 
    0.171596495778319, 0.146005166943493, -0.156704930942655, 
    -0.69584272498274, -0.295018918840926, -0.844271597676474, 
    -0.542807374943983, -0.0819556079764716, -0.400556901089577, 
    0.0197171950134978, -0.865571612879177, 0.530891964819311, 
    0.0379169705052762, 0.447281203607472, 0.364240539850837, 
    0.726725618272273, 0.671660618301249, 0.192480530744561, 
    -0.0799054890946094, 0.875431726226235, 0.773735136109823, 
    0.59345215169091, 0.35823284038945, -0.925048073428667, 
    0.240626691017702, -0.145323599360694, -1.13559748351694, 
    -1.50593608686706, -1.16066622512351, -0.330874859249, 0.533067934400355, 
    0.77564236614371, -0.224109349854844, -0.563202211921858, 
    -0.51128958656979, -0.355925686224263, -1.15699583381335, 
    -1.78568956070317, -1.15502730294208, -0.901023156299652, 
    -0.532929647241271, 0.238737223929138, -1.10469217083499, 
    -1.9127716195548, -1.45066278534617, -0.26778507905628, 
    -0.209556593129134, 0.212133446775846, 0.185768493144476, 
    0.368394113822141, 0.520100033282151, 0.251848521440996, 
    0.0686789577337432, -0.660607188618569, -0.498658339611504, 
    -0.464203865934461, -0.995760202588607, -0.236856553628177, 
    -0.365543700655033, -0.526485510853214, 0.306684437834228, 
    -0.300714255118648, 0.606860619654781, -1.17379971887849, 
    -1.08236435135289, -0.505925378748517, 0.297535385000356, 
    0.965782434423121, 0.282260166729533, -0.104625754528573, 
    -1.1671844214551, -1.06108315125132, -0.659607340231068, 
    -0.990302080966887, -1.91138718897067, 0.52083199096177, 
    1.24160367494726, 0.619068934837856, -0.0424798385884495, 
    0.149740039096611, 0.99341342176642, -0.222380648692981, 
    0.0594853092875569, -0.651345766116065, -1.16525434192253, 
    -0.686487390191277, -0.488055018794711, -1.05701680878545, 
    -0.863705137587711, -0.422121300670937, -1.10159310886915, 
    -0.692309107257572, 0.126766460318524, -1.34083100594471, 
    -1.44391798592138, -0.889273497931464, -0.191252010249237, 
    -0.58240368053232, -0.135613101334728, -0.354631029904988, 
    -0.149289639359056, -0.566208164389819, 0.501174441564523, 
    -0.503920390647066, -1.30466675108408, -0.771663311312145, 
    -0.59277962199233, -0.620550842346299, -0.338845437060344, 
    -0.384174305022227, -0.622992855950462, -0.0687689797292812, 
    -0.0702887128180185, 0.761132467473566, -1.78076054358834, 
    -2.13682198407128, -1.19164381887691, -0.00642062259054832, 
    1.47924514848138, 0.391767340131222, -0.462140876936421, 
    -1.68375151088974, -0.760321530211918, -0.0580445989550915, 
    -0.495905172277138, -0.622147499619135, 0.713129760949962, 
    1.43866946368918, 1.60860913636797, 1.27177317532685, 1.73756224404745, 
    0.821961899494945, 1.88277122170907, 1.43095358823623, 1.35895693031412, 
    0.286725891152604, 0.232735954661418, -0.0517290005119975, 
    -2.1038417061551, -0.848445641701017, -0.0790030874128611, 
    -0.0770833529584673, 1.04375866791346, 0.200730157120257, 
    -0.010561893134033, -0.361018494270788, -0.0583269195101188, 
    -0.469316126929806, -0.594141370550476, -0.902649123431756, 
    -0.876743089326499, -0.615906125933403, 0.482393549437719, 
    0.433982127458714, -0.25742890796697, -1.29894114015513, 
    -0.466761740291521, 0.299377728394021, -0.364313744140707, 
    -0.589934782325079, -0.544869929334491, -0.328138695908731, 
    -0.292711736092897, -0.528312773533917, 0.262804486570225, 
    -1.95185212095915, -1.90799958610111, -0.990015954860439, 
    -0.140918679083062, 1.27149865082353, 0.503955692901195, 
    -1.47037501185724, -1.95977935062587, -0.797853597362019, 
    0.0818570667587259, 0.41127496971411, 0.226002161134011, 
    0.505991410228801, 1.02618607832938, 1.1242051240611, 0.751020195228391, 
    1.08431141272843, 0.719628508175325, 0.985727682414943, 
    0.916633198933301, 1.39629981757893, 0.655884908019129, 
    0.581010826866688, 0.292296585877665, 1.11791832017013, 0.89060940525793, 
    0.650005595251448, 1.14064840063756, 0.177065432164545, 1.63648275538664, 
    0.159503153806422, -0.917885828150649, -0.784512456193776, 
    -1.13889385618833, -0.944107264561564, -1.03795977379569, 
    -0.81354218364714, -0.678976497159081, -0.265487585497564, 
    -1.00784051804516, 0.648506647570257, 1.07134923195823, 
    -0.0718876707055616, -0.479231748855162, -1.09277312339151, 
    -0.71223829929008, -0.972507323486624, -0.801094893487888, 
    -1.07869520024354, -1.76297683036285, -1.37311064566343, 
    -0.770105940523389, -1.10529016707697, -0.418066161290991, 
    0.303425028360995, -0.452141896916398, -2.02733159841605, 
    -0.698424273453675, 0.128381382988225, -0.521204477841932, 
    -0.597751949234859, -0.381570474191095, 1.51463822944528, 
    -0.243141500315933, -0.434794364004429, -0.432501928007261, 
    0.10015338878822, 0.822651598360165, 1.88850610790088, 
    -0.654705429832493, 0.732230231800188, 0.22916449846389, 
    1.65238165528909, 0.252703866039266, 1.12460474442399, 0.390670823280903, 
    1.08528199384651, 0.274818413832419, -0.570725874812783, 
    0.0574693567980049, 0.0525736355879403, 0.00939872292971031, 
    -1.45922748406614, -1.48063121766699, -1.26552643601888, 
    -1.38412294454471, -1.67604759595136, -0.595585103823302, 
    0.562584991232997, 0.0909025391580798, -0.73359442596626, 
    1.25270601319167, 2.01970272753492, 0.772695790058626, -1.0579210111224, 
    -1.50747316403637, -1.60727440210767, -1.80689773392758, 
    -1.07232693117175, -1.4166109646794, -1.33726968903946, 
    -0.427369291332109, 0.00089760184840415, -0.894039541348222, 
    -1.17117044568089, -0.59248876276738, -0.415899329960219, 
    -1.21177100444969, 0.137425629664283, 0.154021300633485, 
    -0.850592025570291, -0.899836672376866, -0.161913470323745, 
    -0.735970664352409, -0.415399494868092, -0.906006145827849, 
    -0.436058874180385, 1.59732368455522, 0.617135773037734, 
    0.682060982589503, 0.247144505015076, 0.733815510526821, 
    1.53811170508593, 1.56392539979723, 0.696502137671886, 0.576809470068911, 
    0.881167250070458, 0.210029452242392, -0.546550249619004, 
    -0.05469092774324, -1.23380215986248, -0.248972608325522, 
    -0.488639524014252, -0.682607878852561, -0.959602271581224, 
    -0.393364612331646, 0.4949989752064, 0.731165867736756, 
    -0.218373983605735, 0.833264410889014, 0.20013039046944, 
    0.0171183064019065, -1.30833603828677, -1.44987521771931, 
    -0.961289593507835, -0.935994710358141, -1.41801050730042, 
    -1.72243106813314, -0.844047715445906, -0.471384264824102, 
    0.00519223561240789, -0.173729447261284, -1.03134464256848, 
    -1.37784252376587, -0.909921791768764, -0.940398102012514, 
    -0.117964612784798, 0.13602703346673, -0.176414890051628, 
    0.35008155696313, -1.04937706270889, -0.7101033210233, 
    -0.193303503734459, 0.705463143799679, 1.80709356243802, 
    -0.344646733730559, 0.381370038025559, 1.09319674946498, 
    0.979607118150608, 1.20943913631747, 3.32024302323322, 1.204795916498, 
    0.579425331578021, 1.31305358829087, -0.680815827265322, 
    -0.490506059582989, -0.502870576573047, 0.0505878852122699, 
    -0.0134789429292947, 0.100868299032193, 1.13306376317418, 
    0.505148507581641, 0.901304945022394, 0.334733678132717, 
    -0.732475562492891, -0.98102373223421, -1.35955398169652, 
    -1.17770807780107, -0.896058197781424, -0.696591899784154, 
    -1.31531894838986, -1.09670677861966, 0.162252834041916, 
    0.0273868456475945, -0.419654222570625, -0.418342218296011, 
    -1.34480886065546, -0.9965322212358, 0.109465120723233, 
    0.449447148704758, 0.507643586877955, 0.583600536522977, 
    3.88825748640375, 2.0645739572637, 1.89791551559208, 1.5936831181613, 
    -0.758379123673807, -1.06343125187026, -0.804192125992982, 
    -0.394451093906634, -0.456646867960719, -0.31925156385932, 
    0.0475835655035706, 0.0714544719515864, -0.175105411894045, 
    -0.603407044700597, -0.360716196295119, -1.23400827793703, 
    -1.57500037175352, -1.17609869986102, -1.17691319693994, 
    -0.608708090976018, -0.733308124061103, -1.0989663590691, 
    -0.0700942094479773, -0.234527027746361, 0.0674672909630525, 
    -1.33816619344569, -1.42546879810105, -1.07870789132325, 
    -0.228417660891793, -0.314191269185429, -0.774405914454253, 
    -1.02061679485535, -0.920431304283866, -1.18497037261359, 
    -1.64914258313149, -1.50322445007338, -1.50120913278908, 
    -1.58103924003251, -1.1900932632822, -0.602144436397429, 
    -1.46151964611246, -1.6802252838788, -1.45345316405423, -1.1299917299983, 
    -0.634551451873979, -0.567013437401749, -0.964062146835558, 
    -0.527366309990485, -0.0977143766880761, -0.284056093389027, 
    -0.435734291110643, -0.843444516219263, -0.0243261579311405, 
    -0.325376688826147, -0.864774387021923, -1.03233663609814, 
    -1.58157631764089, -2.14021849153041, -2.51506600751655, 
    -1.60616245906295, -1.93258582400492, -1.87816010904749, 
    -0.76024350536914, -1.15714016245292, -1.60599507680367, 
    -1.33254622208207, -1.54680713801715, -1.1903166376327, 
    -0.841561850331756, -0.390028622550029, -1.16174562015425, 
    -1.15201685395934, -1.55884327425443, -0.864921719862912, 
    0.0107206770456125, -0.83387629485987, -0.995408311814572, 
    -0.659705274914915, -1.83363004217008, -2.2842021527233, 
    -2.86709595449253, -1.23394568206853, -1.77274464371402, 
    -1.45011711490401, -0.661367910456785, -1.46556144688295, 
    -1.10578099128577, -1.75079187746441, -1.8239634120757, 
    -1.04631246069292, -1.09817140903429, -0.781818356848141, 
    -2.14786911096678, -2.62347875473369, -1.12912050212065, 
    -0.650915072796638, 0.936286694745569, -1.24860707006134, 
    -1.05591361368241, -0.387990686879753, -0.569511737598294, 
    -1.49662671300736, -1.52664040919829, -1.30687493164869, 
    -1.74347892706447, -1.4207571784965, -0.696442460995681, 
    -1.47346605628884, -2.36123462013103, -1.76756424287679, 
    -1.23711457209459, -0.92745352498119, -0.890166624974289, 
    -1.13306202234686, -2.49145502802333, -2.63993540119001, 
    -1.05296815748523, -1.15319597397002, -1.12293082769611, 
    -0.774492193866179, -0.299030734429948, -0.397515092028975, 
    -1.12962581203837, -1.61283457019784, -1.62784929784934, 
    -1.34127401091736, -1.13863988666755, -1.66015361197199, 
    -1.75942880112256, -1.56707962663132, -0.989861459708505, 
    -1.17742140522239, -1.24644498539773, -1.16572409127576, 
    -0.793495212896556, -0.90269920937017, -0.790549512571719, 
    -1.07046295863316, -1.37817532288016, -1.11223521288879, 
    -0.923230195477562, -1.68689009758457, -1.77700454453141, 
    -1.44135850606868, -1.16510789722093, -1.09629357763609, 
    -0.754078291810494, -0.927465952943174, -1.81141115957664, 
    -1.40689776715901, -2.00028794955097, -2.03656726901753, 
    -0.8567017271307, -0.97465097793545, -0.854553274730154, 
    -1.36339612219772, -1.39829647634276, -0.689800698771661, 
    -2.45740080551664, -3.31458501640432, -2.21847004561811, 
    -0.202438361696413, 0.0562817353637479, 0.44746123029471, 
    0.593875500153387, 0.436594775248871, -0.124817127578054, 
    -0.507343565962795, -0.869023285322132, -0.964695487022373, 
    -0.845433680154226, -1.37248947929489, -1.63013603395808, 
    -1.05425636111248, -1.99866967381472, -3.63060386359508, 
    -2.29129855835259, 0.367795445502415, -0.311225452153527, 
    0.711346004638505, 1.70019540267168, 0.220321979484037, 
    0.230450909423232, 0.433458315596975, -1.32736580710181, 
    -0.950115060411796, -0.188059351304255, -1.44737941684017, 
    -1.0818188956648, -1.66532387613284, -3.03331475455691, 
    -2.37811775955625, -1.08295143501154, -0.84349629223023, 
    0.445464417554096, 0.575576727563152, 0.583536252549415, 
    0.549854099528653, -0.632675243317236, -0.356788214418584, 
    0.384729586596788, -0.82630428958538, -0.65979699462539, 
    -0.494396996136253, -1.65878898539506, -0.940337955757973, 
    -1.06510200871203, -0.870108152441054, 0.0680813527799051, 
    -0.27691475537726, -0.208146720086155, 0.390027911743012, 
    0.57036213344956, -0.403708798991596, 0.23325630731005, 1.22265905825154, 
    0.897395369107721, 0.773178073511813, -0.591260430055383, 
    -0.233467572975989, 0.0287900316296064, -0.399339804166088, 
    -0.188206051636337, 0.404153493897921, 0.198519175965224, 
    -0.512448110729444, 0.54146828151151, 1.14345805012082, 
    0.281405702977877, 0.67098580309727, 0.0763228666504823, 
    -0.0465951627138139, -0.257794796561623, 0.502285791281403, 
    0.547084395313151, 0.0255811940794359, -0.283605144513519, 
    0.178733468528827, -0.169937459015022, -1.50576877915051, 
    0.0787609030906467, 0.634355057436622, 1.04215051441943, 
    0.435853570564033, -0.4842992657826, 0.244319228256291, 
    -0.401077388159261, -0.348768203088103, 0.659580100941941, 
    0.155009883208148, -1.7542658407424, 0.410300520297713, 
    0.357389431945019, 1.17625249641079, 0.409881175424309, 
    -0.382733236406239, -0.585530631206996, -0.360104965677852, 
    -0.197736486948639, -0.18776313872733, -0.829406563676098, 
    -1.33889786392341, -0.652237792189245, -0.429163660055654, 
    -0.405868390008028, -0.888518646108598, -1.21501092523384, 
    -0.562859398447837, -0.451724356996013, -0.624206247824461, 
    -1.70877972705889, -0.437438474622462, -0.830324022529183, 
    -0.972611856122363, -1.52706821419287, -1.64032648751388, 
    -1.18797141335881, -0.0876551668135894, -0.161685204611191, 
    -0.091332006552971, -0.380435503252046, -0.747343236313704, 
    -0.836501923800403, -0.489747331943873, -1.21272062846144, 
    -1.72974103760674, -0.164450854039511, -0.389721027498244, 
    0.151274323342512, -0.253831154262794, -1.08810931342324, 
    -1.67792576151414, -1.35359100251712, -1.15585945700906, 
    -1.02414330842699, -0.392994694124926, -0.873007741205951, 
    -0.741629198651403, 0.197868395941465, -0.726162403463504, 
    -0.708228188118176, -1.57449194631279, -1.07449663615024, 
    -1.07160143946225, -0.998634664496683, -0.952263097456862, 
    0.142878935680693, 0.732278296413624, -0.287885799890812, 
    -0.667700767091959, -0.761025732203021, 0.190134030511939, 
    -1.23937735434673, -1.01209359752449, -1.6077991520469, 
    -7.45172375188741, 1.1549513262704, -1.56050966376131, -2.31226245106552, 
    -2.98795750199713, -2.81111090763499, -0.466746653569539, 
    -0.511870795065024, -1.87952911879901, -1.92238871234138, 
    -0.825079229874826, -1.09701753747932, -0.2622892710701, 
    0.931889227675931, -0.476452786436483, -0.222723570464965, 
    -18.2237758790698, -18.3599023606526, -17.3642473444502, 
    -10.5752825194152, 0.0505198455966285, -1.04162530832651, 
    -2.04281640407443, -0.675441619762296, 2.85827534724632, 
    1.89618699084946, 0.415325613008122, 0.338249968275761, 
    -0.705057441346923, 1.20680539017926, 0.672549773824471, 
    0.607493441381024, 0.378200714263954, 0.322670338525643, 
    -0.399202907718177, -1.63900152592621, -1.17303291598988, 
    -0.51710048884912, -3.40970830068468, -0.467018583151062, 
    0.3392101309678, 0.934358086526972, -1.72181308727888, 
    -0.585827195744309, -0.317387938694066, 0.518135101874719, 
    1.80551983944772, 2.17562840528973, 0.500390431856892, 0.628584076649106, 
    0.842750897732496, 1.41608540445834, 1.24394704161474, 1.00084594199883, 
    1.71613259625015, -2.85929562008462, -2.71668796350895, -1.2407493468416, 
    4.21733397532975, 3.80021863820017, 1.65412244875495, 0.540354666074186, 
    -0.806590195496106, -2.49762515217853, 2.69476996200524, 
    -0.00454755118468597, 2.080046470995, -0.143791668033089, 
    0.891407444187564, 0.535687167042198, 0.301584279712586, 
    -0.43341343597163, -0.190935219748667, -0.126720949344872, 
    -1.02224302036404, -0.122035056365517, -0.686432637227181, 
    -1.66455208422828, -1.14430692790909, 0.500370563195691, 
    0.0378999480712672, 0.044090598823594, -0.415810930584382, 
    -0.813978427264486, -0.384647701072529, -0.139857488927086, 
    -0.368541112269636, 0.0443580264920485, 0.103669962707014, 
    -1.36747922875166, -0.297435342190382, 0.33199049811607, 
    0.407214105299381, 1.17096046156445, -0.212725377688185, 
    -0.219257333027341, 0.194040462497349, -0.243575952253501, 
    -1.0724149955779, -0.612285906815102, -0.328528435491946, 
    -0.596881489225849, 1.89455837140807, 0.457176749823316, 
    -0.333862065822284, 2.18229233470027, 2.95556564521055, 2.26805739071007, 
    0.307494671300441, 0.331716405795786, 0.736040107782001, 
    0.474192745018849, 0.631177485052801, 1.08085731747047, 
    0.441511526098801, -0.461741329306555, -0.413298631477401, 
    -1.23332753721181, -0.896951653945566, -0.813332167772818, 
    -0.840241443075724, -0.464616976759471, -0.180878003862093, 
    -0.354847633146358, -0.23739897262268, -0.276758647851154, 
    -0.507164662936583, -0.199096754877512, -0.617001367298, 
    -0.626677196804151, 0.0469033632164884, 0.336481838718106, 
    0.171338373549021, -0.628760843910703, -0.881559336892899, 
    -0.166997206561161, -0.288398818726918, -0.372794354580916, 
    -0.40706770671771, -0.334302744297736, -1.79497927029878, 
    -1.01235584058977, -0.043804132264964, 0.258387075970359, 
    0.568569225898474, -0.440127895766427, -0.55276245882697, 
    -0.274814893293844, -0.664423617332695, -1.33720261255344, 
    -0.833713398179148, -0.244488069445463, 0.398540875192674, 
    0.724692439186088, -0.248150008260835, 0.181304268049023, 
    1.12762560536495, 1.28283924635179, 0.205654845975096, 
    -0.915775297297574, -0.161191745282125, 0.0887809670620143, 
    0.225850258977713, 0.112885492472694, 0.580726583770934, 
    0.013648991380828, -0.378431988509953, -0.680608356901993, 
    -1.13697736271297, -1.39191071727719, -1.02836207287667, 
    -0.90125998767479, -0.208798259718783, -0.0966010759877056, 
    0.357878439517672, -0.215967795021919, -0.597025110004461, 
    -0.276692669455532, 0.0914095375165225, 0.117110537518581, 
    -0.896835968095173, -0.832222913528122, 0.166099705841551, 
    0.344498949346796, -0.647756836509412, -0.980839149113315, 
    -0.15542787174037, -0.573352823519198, -0.0588920151543526, 
    -0.89794187181981, -1.23413235788767, -1.39562959485276, 
    -0.470386820709643, 0.0672758789619277, 0.0752222758797583, 
    -1.25453269540299, -0.961796087251936, -1.16619449738739, 
    -1.34985324864286, -1.1640345860795, -1.19747746114812, 
    -0.27708428354746, 0.360152437505672, -0.0147749912578066, 
    0.01705771635697, -0.947379166610363, -0.809251601088112, 
    -0.204757741643187, -0.0408817613068413, -0.759607620674907, 
    -0.878343241708408, -0.272557639582951, -0.518411349132442, 
    -0.692579816182564, -0.407657487505233, -0.111047235369197, 
    -1.66107585630452, -0.572958695103107, -0.784756676406051, 
    -1.34757807923708, -2.3453568123257, -1.68945997419002, 
    -0.42849465687981, -0.260481709594282, 0.81535143421124, 
    0.195198738167499, -0.567123135925729, -1.21915100882337, 
    -1.06396669451078, -0.503290831198822, -0.649568022661011, 
    -1.30908624979284, -0.855837395505921, -0.418730345110276, 
    0.0927736131116408, -0.439722157076101, -0.615935688960523, 
    -0.448072122303662, -0.611857618642966, -0.0535661101310936, 
    -0.693711354535043, -0.968233965749135, -0.524065048560378, 
    -0.967980610614072, -0.0135622321135509, -0.870130791021166, 
    -0.321883838377932, 0.65618160751348, -0.293775051920782, 
    -1.27907702777557, -0.506262369144599, 0.0161447219231148, 
    -0.261132451744772, 0.660746073644152, 0.736499532104449, 
    0.230844281407814, -0.6301065078158, -0.0981264132352022, 
    1.05789722043785, 1.00507496307397, -0.0167186992290924, 
    -1.11287728236033, -0.0342067723577388, -0.793536501512944, 
    -0.166256376936396, -0.587915047769134, -0.482714060683995, 
    -1.43555728898985, -1.9083588742215, -1.35851185378755, -2.1631135455691, 
    -2.62936064593071, -2.02102026606515, -1.06021714909816, 
    0.0383032544393158, 0.0867570754738356, 0.00701303487605998, 
    -1.16546234562553, -2.41621602720318, -1.4815333077696, 
    -0.856168624804443, -0.594974544390441, 0.0140265579626142, 
    0.281904956158296, -0.588883460498035, 0.648220999197893, 
    -0.225691859215207, -0.57039376824398, -0.983067381726559, 
    -0.756377323489006, -0.269408122668331, -0.414376055875207, 
    -0.435028018731121, -0.374816308435784, -0.891288643378978, 
    -0.460476080222776, -1.46048271889587, -0.986376953445784, 
    0.0204079727918005, -0.280239763173391, -0.798277526722693, 
    -0.695458340272244, -0.0600508143526657, 0.590835919591886, 
    1.04327195599358, 1.08226240413248, -0.987325478367671, 
    -1.10134170080387, 0.0315078438391447, 1.58093637308858, 
    1.69186898975502, 0.670477775247851, 0.1249271131103, -0.545078588101551, 
    -0.710187058686538, 0.388495929240671, 0.50234479283513, 
    0.439342041861104, -1.46124840272273, -2.09101726354464, 
    -1.63770153753628, -1.93844854541482, -1.50663951150121, 
    -0.470346821848113, -0.162904011192171, 0.155151800585234, 
    0.132076417431222, -0.439760705782004, -1.30947407398666, 
    -2.14121893597568, -0.542940780140775, -0.286642279239988, 
    0.242644788714745, 0.197520409258125, 0.48820405863653, 
    -0.688983819250302, -0.223319221026861, -0.594608495892803, 
    -0.751331457253666, -1.21673416144065, -0.763925452844645, 
    -0.282083546016998, 0.0635915154594713, 0.370953579498181, 
    -0.141009377254755, -0.284038593728142, -0.0377687013293647, 
    -0.653591903531292, -0.93972087652054, 0.120745597271661, 
    -0.134210952738476, -0.0938910665582426, -0.281608452336899, 
    -0.0681027194511552, 0.605924431926059, 1.33239401025024, 
    0.731055102665508, -1.13251838453318, -0.844957162888118, 
    -0.334488442969074, 0.832576873318103, 0.620588769944224, 
    0.450370625010081, -0.571045622269457, -1.24680365096213, 
    -1.55415726279385, -0.677262200339595, 0.171544694991446, 
    0.622313859980816, -1.17112607857391, -1.84405270671736, 
    -1.48021422930178, -0.821647077315566, -0.828221220043304, 
    -0.170402317965039, -0.102071622433559, -0.0228334176160372, 
    -0.0658411194789688, -0.759976868064558, -1.1744842154514, 
    -1.82943555935563, 0.110541579250896, -0.578996895967645, 
    -0.568222283615434, 0.27310298161213, 0.248437962306403, 
    -0.878987480211428, -0.371843217421137, -0.401097137382349, 
    -0.506271603076529, -0.721577138662277, -0.464995940603257, 
    -0.470118525672163, 0.450886677354303, 0.219130390093687, 
    -1.38265281113069, -2.1320144511214, -0.17579304294573, 
    -0.571095267554576, -0.731371759221173, -0.866959966063305, 
    -0.526771731441471, -0.0188446982674861, -0.516154721894293, 
    0.0471492805734108, 0.607568636954112, 0.359997874081528, 
    0.339857189794026, -0.662047799656031, 0.452009082745337, 
    -0.147361024837851, 0.0124054720107036, -0.430646294628003, 
    -0.307959814936192, -0.381060228747265, -0.596347470778564, 
    -0.367138185391913, -0.112693896956508, -0.1646937395385, 
    0.54365137168682, -0.956536896908986, -1.12774670877263, 
    -0.955543955216704, -0.668382464884911, -1.10471902348187, 
    -0.414369511405548, -0.472851854978549, -0.583793822061418, 
    -0.535916794785014, -0.403327840926133, -0.506759110218122, 
    -0.985499135880752, -0.699989102799048, -0.790072038714369, 
    -0.508823065420581, 0.671406508335375, 0.0460166569248877, 
    -0.441468231570594, -0.30885860776606, -0.301331448365403, 
    0.164394864044755, -0.386977162848674, -0.997659176756169, 
    -0.656010136338661, -0.0511140493261086, -0.0328284385512001, 
    -0.892083737674665, -2.08413043084133, -0.387771108079358, 
    -0.733396645879614, -1.21220642558207, -1.04284479458641, 
    -0.433431146358658, 0.242096062687462, 0.305007898582543, 
    0.992367527000027, 0.281437366877983, -0.0575551803129359, 
    0.277269949181016, 0.171204851326365, 0.391163425281182, 
    0.554729676492536, 0.414304042035867, 0.0545476205401707, 
    -0.59575321517781, -0.739830853799548, -0.292727502143704, 
    -0.0586670028621761, -0.119057047961539, 0.275051493929195, 
    1.08478994079527, -0.618883235311363, -1.04381478770743, 
    -1.38257961395382, -1.01223697290855, -0.71991782599877, 
    -0.509675295113916, -0.267722520444678, -0.747438969554217, 
    -0.669793224861337, 0.221696280096531, -0.436718672372347, 
    -1.60371570016093, -0.648580260128959, -0.460913419307571, 
    -0.638246505796793, 0.113113238825706, -0.0132007329998984, 
    -0.0583924931215574, 0.135855591937855, 0.0244635635977009, 
    -0.0207067898847635, -1.35684030351326, -1.95555371243245, 
    -0.592741876487852, -0.76326090199097, -0.514646848530109, 
    -0.392087146280007, -0.0268566249318392, 0.0311307507441105, 
    -0.237154252899829, -1.31055911265728, -1.07200274544875, 
    -0.0322395046111046, 0.543635845972741, 0.748280384418685, 
    0.702748810097402, 0.0695303682493487, 0.269916629105665, 
    0.313585176361824, 0.585411846704611, 0.24688358452396, 
    0.191672591178347, 0.401132789754568, 0.365673308168413, 
    0.013517208748377, -0.354658951952671, 0.0480989913968077, 
    -0.870546835069486, -0.0311370704805025, 0.619184479204105, 
    1.0272148235789, 0.233729038823882, -0.853394484298104, 
    -1.94212194669309, -0.993057548590217, -0.506783180522272, 
    -0.448253320514191, -0.124644233737548, -0.712393801997271, 
    -0.121243052678865, 0.437228476482714, -0.429293357822645, 
    -1.90957696418527, -1.17483009521631, -0.345117374427568, 
    -0.0237180294066874, 0.415260911907369, 1.26229377232925, 
    1.11550505371848, -0.0163504946404558, -0.718408843780454, 
    -1.0856085986323, -2.01989505056313, -1.57266529929111, 
    -1.78282736469886, -1.65801214902175, -2.48865130779782, 
    -1.90445324032082, -0.216350835289515, -0.471101237150369, 
    0.151706564721579, -0.907720532917051, -1.00814862029559, 
    0.0377999641132565, 0.610784271744551, 0.909543593784723, 
    0.903312568351358, -0.125650110595896, 0.386206459804947, 
    0.418545068093215, 0.527385056231928, 0.78087297567258, 
    0.0198206218318564, 0.358682611848518, 0.521180807688477, 
    0.00262035641790614, 0.446401486600925, 0.505871098551243, 
    -0.394887718508596, 0.233989739708962, 0.367311842687066, 
    -0.636560633949554, -0.487347862175462, -1.57814001695321, 
    -1.04807524592681, -0.745517659216288, -0.716172967342597, 
    -0.0185978182293089, 0.072410517848005, -0.786254770282246, 
    -0.38768470846438, 0.259021702622397, -1.71588728292708, 
    -1.94044015692012, -1.44861954794673, -0.62087235243288, 
    -0.385056468133662, 0.619803824229423, 0.149462188564815, 
    1.00093740193936, 0.178005095519351, -0.285762777780407, 
    -0.761366714626357, -1.28854780402863, -0.813779541549193, 
    -1.69407159452188, -1.50532293852896, -1.78220554647454, 
    -2.42842500985595, -0.682842789554834, -1.20403068417266, 
    0.0378314022676474, 0.0309789458465426, -0.184108745613107, 
    0.0944111114127022, -0.158532874258834, 0.00629633322095202, 
    0.00304459307605587, -0.372137243316355, 0.473110498898963, 
    0.475706134921845, 0.743578524149822, 1.15396159910641, 
    -0.0839714905583813, -0.290943136186645, -1.14320242017928, 
    -1.03905657651451, -0.702666087579629, -0.726608251550256, 
    -1.06797955354735, 0.515923198457622, 0.6503711633147, 
    -0.733240588215782, -0.690679727316503, -0.854748715082283, 
    -0.585983437637383, -1.1409560731024, -1.32261092138816, 
    -0.758625480256216, -1.17697604538372, -0.707568496868518, 
    -0.628234294550092, -0.692160789656318, -2.1555655050674, 
    -1.80987256030743, -0.93522250275675, -0.414014086529368, 
    -0.212920341125864, 0.0147785070993667, 0.146335910819815, 
    0.0933057785824687, -0.245618070789977, 0.0110612005868393, 
    -0.552997701672475, -0.922677559352834, -0.471854178976905, 
    -1.08330573662445, -0.749328868230132, -0.293414678383614, 
    -0.680923466550993, -0.375503288366579, -1.19048773739425, 
    0.224279376882248, -0.285525925384262, 0.149380709232227, 
    -0.0399868645396007, 0.266537807390113, 0.185123498813895, 
    -0.24305525927613, -0.264433060289111, 0.541465514441861, 
    0.696532196178867, 0.190178455553802, -0.194090655288637, 
    -1.77886425792594, -0.107733256618254, -0.426262100553063, 
    -1.55787494347619, -1.9434219843665, -1.70030686881483, 
    -0.829174428303054, 0.021668313435641, 0.385883053487857, 
    -0.616465804434347, -0.889284051884949, -0.819407223344251, 
    -0.757416088290688, -1.3658482993996, -1.84053428149888, 
    -0.9266515135204, -0.86410119704905, -1.18383393919303, 
    -0.0184083636838418, -1.58088504517908, -2.30129061051092, 
    -1.89432488086285, -0.584492684444271, -0.569214406980683, 
    -0.223962767834855, -0.165731385114638, 0.0944800533832169, 
    0.517724316370165, -0.232495607694752, -0.171761971401878, 
    -0.848710731780491, -0.813521521327836, -0.676971257731656, 
    -1.1524783393861, -0.554558754148515, -0.622896800790493, 
    -0.751422538909652, -0.0560810273856172, -0.550942863070261, 
    0.296368643022991, -1.56853641632664, -1.46693778162269, 
    -0.767352775725043, -0.125985105842186, 0.566443367862686, 
    -0.0684406039673213, -0.421468003093164, -0.886860823168814, 
    -1.05238434640474, -1.05906602708475, -1.46916713568187, 
    -2.34578423173616, 0.281586162715959, 0.936085881280446, 
    0.402920436265681, -0.371216416292683, -0.357664331248326, 
    0.530525111921234, -0.585127042854334, -0.24553790760713, 
    -0.897381993933655, -1.3703182663187, -0.979541164135562, 
    -0.853958890429842, -1.36008598092804, -1.01496300549311, 
    -0.676566887221992, -0.886952516208281, -0.309805794004481, 
    -0.114222917264085, -1.78910795038365, -1.83461779611846, 
    -1.34708330733599, -0.57483918826617, -0.999044400488183, 
    -0.764240148698843, -1.11562894873226, -0.343451319372505, 
    -0.759289906383396, 0.112411994963999, -0.840942815431545, 
    -1.80006640656648, -0.992860611656954, -0.882575458418944, 
    -0.894633817835069, -0.59863479794303, -0.687973135307738, 
    -0.884066136882047, -0.252649174801927, -0.256507501683321, 
    0.460427378065402, -2.04275606500964, -2.52133162159865, 
    -1.52126629369095, -0.227035815270216, 1.24462576184849, 
    0.0104264758549322, -1.05947103757742, -2.30836493131618, 
    -1.01109775605904, -0.242710449757761, -0.74448629235182, 
    -0.871212305488632, 0.44504658361562, 1.28568634789544, 1.35400955520225, 
    0.969345848079803, 1.40057157690073, 0.442566202014323, 1.50235163360633, 
    1.078070241411, 0.832695232783189, -0.0189454272741063, 
    -0.146378088032204, -0.410086262625029, -2.189189341371, 
    -1.09735046340608, -0.493577344755201, -0.352199926335001, 
    0.701187041709104, 0.0490887098363279, -1.18468101751835, 
    -0.89271590198702, -0.465479793863262, -0.911238012773294, 
    -1.136113946029, -1.46556956004475, -1.38173676754048, 
    -0.592019684509575, 0.591921007675564, 0.243146045484313, 
    -0.414131897574719, -1.50719774846268, -0.44332698135281, 
    0.235598069555709, -0.54438350516226, -0.832591137780545, 
    -0.858071725263807, -0.589883855367956, -0.447507172117745, 
    -0.769381997823997, -0.0279850652158009, -2.18833701325796, 
    -2.30374787435426, -1.28086806477445, -0.435379812961383, 
    0.834031842720817, 0.028049491995672, -1.73052526935489, 
    -2.35480907646346, -1.00869947620298, -0.221018920664879, 
    0.206504128803218, -0.0625131097836018, 0.196904891943555, 
    0.847916094188972, 0.677011882036158, 0.0453743319796285, 
    0.697882390592843, 0.336427282127367, 0.727960015399685, 
    0.619535901368886, 1.06490371961112, 0.343067038472835, 
    0.222022178153019, -0.0961572239550446, 0.860353045452322, 
    0.569308061164935, 0.245372174027092, 0.516204581061142, 
    -0.383777664810716, -0.0701675052309536, -0.188286580623616, 
    -1.40223051396461, -1.38357845106018, -1.66086687660495, 
    -1.46313364039005, -1.40543865228852, -0.475410570772334, 
    -0.377274934120209, -0.641555633266471, -0.929642053224762, 
    0.636545914034436, 1.19429095812019, -0.107269033798221, 
    -0.843746854867335, -1.44035514073422, -1.10447968722792, 
    -1.23764213019497, -1.12982186469018, -1.33695492852234, 
    -2.10163990975778, -1.58716963792356, -0.965062541201465, 
    -1.44090223895017, -0.535408733342138, -0.00954810427038932, 
    -0.825389019998908, -2.25718380698063, -0.800778624748673, 
    -0.147598156429791, -0.868310671324588, -0.865382232295704, 
    -0.475741002094181, 1.41759245073229, -0.286942752789336, 
    -0.855725452593177, -0.734658180900655, -0.251098871748239, 
    0.612735992135396, 1.52771142559161, -1.05466187810588, 
    0.385220021414852, -0.104307214935075, 1.27539463017973, 
    -0.152704024933499, 0.603654879524607, 0.104490661239214, 
    0.576575324856607, -0.183376167775043, -1.1030918124498, 
    -0.286248134923742, -0.518264121719687, -0.283326674553046, 
    -1.9088026310761, -1.69447065758727, -1.71424527143865, 
    -1.80124202458332, -2.16284403657934, -0.436539529970004, 
    0.905907727256272, 0.00296678505675274, -0.867335680446444, 
    1.14920869976867, 1.91418437956299, 0.742892916838054, -1.42764248123069, 
    -1.76967771395208, -1.98925307980979, -2.10190046466492, 
    -1.54863011701942, -1.804293152669, -1.71400548583373, 
    -0.856636288473349, -0.414447449488571, -1.11839513254329, 
    -1.37486335002578, -1.00063658029231, -0.773255471188041, 
    -1.60143691418931, -0.066871160430213, 0.110734515343647, 
    -1.03326239615232, -1.10813526108437, -0.532527142696919, 
    -1.1175003706309, -0.653391758869495, -1.2370574738289, 
    -0.509206230374026, 1.52760503204854, 0.537970260447276, 
    0.448748948718394, -0.0399610403530293, 0.448473604704072, 
    1.04137376555847, 1.10239165888267, 0.155261351179101, 0.07846649065407, 
    0.593900093579387, -0.304034090322353, -1.17502207746918, 
    -0.642204887970487, -1.58515241529638, -0.57794116907556, 
    -0.799218416531913, -0.927991007809741, -1.02334767293108, 
    -0.420965675105838, 0.40304204730484, 0.106350984375521, 
    -0.775880167458034, 0.898453532928944, 0.23405840303024, 
    -0.131380034297344, -1.63867958873223, -1.72143892032983, 
    -1.24468305541834, -1.33591358347165, -1.74660141492426, 
    -2.09473710708139, -1.34658150914164, -0.906976940234947, 
    -0.443325423062748, -0.586486723870747, -1.4386674882, -1.68892717409849, 
    -1.1519289776915, -1.28372520656943, -0.609161208743836, 
    0.0911641237888761, -0.35380263909182, 0.245300503465592, 
    -1.22489266100796, -0.824471070053226, -0.277322427991291, 
    0.693147457732003, 1.6122547860223, -0.467717176012231, 
    -0.0438192773964996, 0.568488023634219, 0.341962649115305, 
    0.36946706569061, 2.70045356914801, 0.723189303119036, 0.122991702417764, 
    0.586577683017593, -0.929120103223919, -0.764546908662957, 
    -0.836321417351575, -0.134937544456273, -0.00906967187511931, 
    -0.039938426793622, 1.06751381012227, 0.66483950706802, 
    0.821609819157265, 0.314055282505059, -0.975567598223688, 
    -1.25331647714463, -1.56767555762906, -1.43628757695642, 
    -1.25348052730138, -0.978916252469375, -1.67168883520357, 
    -1.58409100535151, -0.482670354911305, -0.540562666241002, 
    -0.592178055159129, -0.63277284061821, -1.59771167314705, 
    -1.28201701350812, -0.144256514587169, -0.0545907423215786, 
    0.390273707446864, 0.376298387829457, 3.61737365149649, 1.59529129892239, 
    1.29188882022688, 0.840006548281096, -0.837591357178074, 
    -1.26767912764337, -1.05123013038254, -0.487960148380262, 
    -0.568644068841833, -0.435639345073642, 0.145429226402287, 
    -0.194252813855216, -0.926835571218803, -1.22812608212722, 
    -0.588749223546232, -1.57092505802562, -1.85880913702747, 
    -1.388789292022, -1.45836913971242, -0.936225646790736, 
    -1.06050360040364, -1.51945155000551, -0.698496794093986, 
    -0.629395419879515, -0.22960862264056, -1.57558800402626, 
    -1.76506663591036, -1.31927009294601, -0.588025922722539, 
    -0.287543926777625, -0.825051597678863, -1.13921054677286, 
    -1.1125167957922, -1.40450770757704, -1.89322822286264, 
    -2.08143000619336, -2.2178062362965, -2.14820358489212, 
    -1.30847732929713, -0.723906840294832, -1.72734733654666, 
    -1.94307606576805, -1.71854685951832, -1.40082041298366, 
    -0.849831453154177, -0.872115631463242, -1.36510799825656, 
    -0.964539710200563, -0.503028556916321, -0.568877255647657, 
    -0.739131493659535, -1.11577103253509, -0.125610920760484, 
    -0.596479218945616, -0.987124507036281, -1.21126169292369, 
    -1.87636717089425, -2.41809620528194, -2.76486525187578, 
    -2.08999185055794, -2.48696759093471, -1.98507699586537, 
    -0.986166117751814, -1.51219488499693, -1.88799971917142, 
    -1.70820696220861, -1.82743547346644, -1.4444824559903, 
    -1.07794010112466, -0.786376603217902, -1.7257992711219, 
    -1.6165661367485, -1.94694088014659, -1.16343238393197, 
    -0.373801897697752, -1.14710811303012, -1.24694532949931, 
    -0.961600503144373, -2.24102714270311, -2.83392568672321, 
    -3.07430892021674, -1.50428353738574, -2.1585403840511, 
    -1.57762382578472, -1.00532214242412, -1.87057868147796, -1.616954233201, 
    -2.15073312476441, -2.16071455643484, -1.31697006315528, 
    -1.30312983843675, -1.29875656970533, -2.88627832966537, 
    -3.0393865337616, -1.48303321029209, -0.756290082890607, 
    0.523864095784692, -1.35173000040942, -1.30574718013144, 
    -0.649713621044787, -0.903054030914148, -1.96315221392115, 
    -1.87034312450369, -1.48948044628171, -2.06671281493046, 
    -1.68540999062783, -1.26694237405361, -2.17792098147897, 
    -2.7516443119134, -2.10115589384665, -1.63947873943284, 
    -1.28339724140757, -1.12150394162363, -1.50663337058815, 
    -2.87776418180981, -2.82632788802036, -1.58766492318627, 
    -1.18058067483397, -1.38393767471119, -1.14876656152392, 
    -0.405781514418084, -0.742518237473382, -1.49845585292069, 
    -1.97913884357224, -2.07935600885988, -1.71364308041032, 
    -1.68596253725113, -1.98545187334658, -2.14752515746061, 
    -1.92988833806852, -1.4236349887093, -1.50933948067887, 
    -1.59606748074641, -1.62060191392117, -1.30224388977426, 
    -0.672714227280773, -1.06443448981394, -1.4512858359558, 
    -1.82135299958445, -1.5667155940976, -1.22563604288557, -2.1635278593911, 
    -2.79365137399998, -2.12367558757631, -1.68998951531789, 
    -1.39432363207209, -1.05582516196181, -1.28024283879674, 
    -1.86707362060903, -1.66976241899638, -2.19292841848624, 
    -2.17803586069674, -1.14562603740819, -1.32507976333252, 
    -1.39037681695437, -1.83225446359723, -1.77489927040784, 
    -1.0385078055251, -2.80043352582448, -3.82731817386116, 
    -3.02742059114323, -0.694949404932284, -0.38732155050262, 
    0.103603805294417, 0.33177636584905, 0.154129824432965, 
    -0.330263666456738, -0.601021851846788, -1.05435744424594, 
    -1.48924849623702, -1.28944345711986, -1.53920283685121, 
    -2.0490401001442, -1.35835996417774, -2.5111086802207, -3.95802353452326, 
    -3.09563478889888, -0.177972802344581, -0.776098858932666, 
    0.112278158836512, 1.42802683841198, -0.0817898216994095, 
    -0.225435109634229, 0.200265589247239, -1.88744592138441, 
    -1.11350143917196, -0.365119087780381, -1.88409557284856, 
    -1.41988185750335, -2.13756400949185, -3.66092295860982, 
    -2.94866291632403, -1.55523030012202, -1.38511672083794, 
    -0.092447795140167, 0.342480568502928, 0.39710811604158, 
    0.249239250667475, -0.999315527435014, -0.519919534400435, 
    0.0437581776131246, -1.55959089023368, -1.18340414283777, 
    -1.055223303438, -1.99954651842192, -1.36153109273313, -1.87045418478942, 
    -1.3867417027381, -0.306496104463916, -0.640767226862722, 
    -0.591383476531355, 0.166825834691009, 0.0692831507388147, 
    -0.831798638452463, -0.0161387256602152, 0.995504341609501, 
    0.329049488406916, -0.0227214483084293, -1.41869050308607, 
    -1.00079450243184, -0.406412157880061, -0.782780872459008, 
    -0.475419559399732, -0.102097189069648, -0.381490279789349, 
    -0.731438908587196, 0.209979808386875, 0.760567567852282, 
    0.00532115475169181, 0.120051728858308, -0.492415283491039, 
    -0.420149770827836, -0.706967376140031, 0.288847361342826, 
    0.208438073386104, -0.428639376514153, -0.605488036313129, 
    0.0508491694251267, -0.495836315811902, -1.82526585014858, 
    -0.175689474837566, -0.0153702948256385, 0.536145519951252, 
    -0.0933139776669023, -1.03194467674425, 0.133713443200776, 
    -0.538082549391721, -0.564996572040708, 0.262134114238801, 
    -0.318795644495147, -2.28326253894544, 0.141269363030259, 
    -0.0203401282751292, 0.619043261429639, -0.206108326728618, 
    -1.21600048832527, -0.660917381531263, -0.40479922057524, 
    -0.526944959451296, -0.81482998146825, -1.38131054108369, 
    -1.87279747941476, -0.990603326631048, -0.977935398730141, 
    -0.889770313556881, -1.54602124030876, -1.71159110989246, 
    -0.930559307506238, -0.855531812771519, -1.02242654446115, 
    -2.12265735491841, -0.74335627304094, -1.14611915819304, 
    -1.27274791567797, -1.75857535191926, -1.95317540469514, 
    -1.44997351576889, -0.53107753016068, -0.528024694776161, 
    -0.36169271077434, -0.838475546811717, -1.05260439624056, 
    -1.23191274588105, -1.06764615785679, -1.40521547120239, 
    -1.92473185605695, -0.366492652613859, -0.724065524584852, 
    -0.194434725193209, -0.306954344573889, -1.27163319485449, 
    -1.91806683438237, -1.85255454299076, -1.55183678587246, 
    -1.27254884646264, -0.621737478942856, -1.12878082093479, 
    -1.25152620466368, -0.137986353847861, -1.05267610290944, 
    -0.902488076208057, -1.5999303207377, -1.11479377693577, 
    -1.39696255809736, -1.3453732274277, -1.40105963923991, 
    -0.193956177249093, 0.463621990588594, -0.709763533946313, 
    -1.11222770071554, -1.66147667616262, -0.229160948882878, 
    -3.77105452402137, -3.64153020088867, -3.30385136315391, 
    -3.41612406009371, -5.61048437472182, 1.6326439187813, 5.24990762355442, 
    9.08734595404086, 1.5601451341483, -2.76482718210268, -2.52643613200492, 
    -4.18180489800997, 0.443576951263243, -2.08184100572137, 
    -1.81257776044387, 0.175950782436765, -0.444994492655608, 
    0.1730318075266, 0.233227934005047, 1.20082398787433, 1.51012543466631, 
    2.42116931300134, 2.62982955144554, 8.25346043597008, 7.97714089270016, 
    7.54914633502395, 8.00652473033736, 12.5574875500504, 14.1220350849387, 
    -1.34040319347193, -2.24851853805887, -10.4710522936223, 
    -8.20528628658934, -0.222783614132993, 0.124987836649382, 
    6.39288125993787, 0.157132586906528, 3.60819693543419, -0.24862729742452, 
    -2.13455865328172, -1.65311076580892, -1.93881150215702, 
    -3.80033000833677, -4.05523232682725, -3.16038659395943, 
    -4.37357450504265, -0.513462456703238, -0.1171367862122, 
    0.23092139468174, 1.41960757190366, 2.52352377820365, 0.81581670816848, 
    1.33328649657611, 1.94467607655501, -2.90265863438158, -3.40186773751047, 
    -3.76980340716541, -6.75731957579704, -3.0832003954084, 
    -1.50985958349493, -2.04446613134764, -2.17378657394058, 
    -1.29751951755857, -1.5146376667222, -1.30224188477014, 
    -0.668896879269871, 0.327344345320455, 0.0748327872829568, 
    0.944000101858309, 4.09893408310893, 4.59595569083433, 5.04417042684437, 
    6.30310182925413, 9.3489769364453, 3.93304405156876, 0.114078261162438, 
    -1.08314194634066, -3.25574067062436, -5.27689986361249, 
    -4.2666823786341, -0.746961787702105, 1.60184302827133, 4.03268417462002, 
    4.20759351986391, 0.892124536425598, 0.777443219682539, 
    0.686714399096644, 0.7942504017727, 0.734055766094599, 0.320638190335387, 
    0.622438365614641, 0.307748214679293, -6.39672578829539, 
    -17.275179202341, -9.85078858485121, -4.73111820031566, 
    -3.99017398837472, -3.47673379403812, -2.22851819428907, 
    0.645922815453888, 8.75434242953336, 7.64775620163926, 
    -0.582422304211203, -12.4398739110898, -15.0181970128226, 
    -8.90418125195007, -7.50286013988583, -6.57498613515374, 
    0.24231431558853, -0.419649069009438, -1.60927930998131, 
    -0.819968549193311, 0.74458919930473, 0.14693230791134, 
    0.108762799688726, -0.490217829720683, -0.599824415196144, 
    -0.26141915315419, -0.219349715449564, -0.364927129546126, 
    0.188159132073573, 0.312750196602227, -1.37795361350634, 
    -0.281479889733083, 0.539203526185612, 0.694139151095508, 
    0.858776423124672, -0.0217564112775381, -0.592916151893341, 
    0.384374207517428, 0.0666831546252089, -0.465227420616312, 
    -0.607257392323155, -0.551665873858522, 0.175274486144059, 
    0.818414055478338, 1.21296474545987, 1.11876383160737, 2.03569743215456, 
    2.77664650007598, 2.31190599590151, 0.0704227663922419, 
    0.0514024783286704, 0.322002745625807, 0.329008520158252, 
    0.149961699740753, 0.470928039162835, 0.251834173942669, 
    0.679269201308244, 0.789589562347026, -0.309924305850671, 
    0.0870610580277109, 0.0261152667172571, -0.0299929047123371, 
    0.134196343195052, -0.134409936805877, 0.199553726924147, 
    0.408176215905267, 0.278159965775115, -0.260580804405448, 
    0.076383663241435, -0.995683226346875, -0.583282293829308, 
    0.0624748344150117, 0.329485141349295, 0.309015158348904, 
    -0.577938994992273, -0.781172901668761, -0.154714714077819, 
    -0.514855169613675, -0.569682073798869, -0.204912365595771, 
    -0.0171049896914566, -1.7806150553196, -0.900536381638362, 
    0.115364582967099, 0.286244899466279, 1.05415882820394, 
    -0.0872994855196652, -0.776324347111035, -0.260236958936484, 
    -0.00569666941212077, -0.896217085571696, -0.8418731760811, 
    -0.126010782023678, 0.412299476831719, -0.293422194536626, 
    -0.150950335306925, 0.662544058284431, 1.68228147604919, 1.6427309539672, 
    0.610973260346639, -0.822179601816329, -0.367267189907499, 
    0.182510021646753, 0.0672982463326743, -0.288877073198197, 
    -0.135867649364014, -0.385791552604964, -0.264202699424541, 
    0.36931509618126, -0.191199433480636, -0.722368811487013, 
    -0.514979824491357, -0.155693452892858, 0.45473566790831, 
    0.363500356465161, 0.749979919066481, 0.201434394102988, 
    0.0511782097402547, -0.173174050244942, 0.623894463414052, 
    -0.0981782511307561, -1.16109885823311, -0.966098243908506, 
    0.112841042752869, 0.305963670179343, -0.68387309728303, 
    -0.926906206670179, -0.153999034791212, -0.701544835546901, 
    -0.140947713540314, -0.0381005091685394, -0.906940227467081, 
    -1.57058307152644, -0.808524317433252, 0.250713328160979, 
    0.383609940791079, -0.581136423304245, -0.847933932794906, 
    -1.09445903883343, -1.29717486047927, -0.860025339437605, 
    -1.00657843714004, -0.538718874516779, 0.402464629364272, 
    -0.279069983402431, -1.17080143336334, -0.471553720289473, 
    0.413895420238748, 0.445041868416975, 0.0995295176420097, 
    -0.897090527836668, -0.750518896509842, -0.634928283861322, 
    -0.519697114150404, -0.486967476493732, -0.674175588824344, 
    0.0162894722456475, -1.22411983536568, -1.12212120944443, 
    -0.911394505757075, -1.01814029155264, -1.64578945930263, 
    -1.1887008396051, -0.00852181302720467, 0.399732973820286, 
    1.20564611818794, 0.678288076715927, -0.162434290794233, 
    -0.762099487098782, -0.605202197417594, -0.184248979090968, 
    -0.757658590835844, -1.49496645529706, -1.02474856659109, 
    -0.466434528652373, -0.223245482930574, -0.501757496575204, 
    -0.340722628898917, -0.286469644562555, -0.866311176619523, 
    -0.201714296015174, -0.369895371501059, -1.20921148186547, 
    -1.03463284399846, -0.801280916530129, 0.174514087192708, 
    -0.98976055801514, -0.61954600376389, 0.482624063146626, 
    -0.290830465543976, -1.58306617225458, -1.10487790610911, 
    -0.413370666082882, -0.451456611583425, 0.481857994458545, 
    0.0183339985131159, -0.643520722642075, 0.0176997641634902, 
    0.435673653068411, 0.747712451199138, 0.224125355589484, 
    -0.419148039974182, -1.07337541701432, -0.449035395205386, 
    -0.809964592775558, -0.305546369666869, 0.23195735651298, 
    0.450014493921191, -1.30181855580911, -1.99332452107719, 
    -1.67963960208391, -1.50853176518941, -1.52931408389318, 
    -1.5359428112036, -0.567420711478128, 0.53909278732053, 
    0.344176506612799, 0.799192990416282, -0.807572934275065, 
    -1.22553070822255, -1.22933944031239, -0.96356439697268, 
    -0.475022673722432, -0.207971446027084, -0.0257894766294342, 
    -0.850127708706383, -0.16478136093049, -0.547591124041924, 
    -0.662310527996977, -0.85802746532909, -0.976413071970175, 
    -0.229120123632733, -0.334817770287454, -0.736199885525513, 
    -0.657708815991613, -0.95603015185048, -0.675965579914299, 
    -1.79981155281177, -0.852994641828824, -0.00526353934283463, 
    -0.323753973295218, -0.699857543952871, -0.847654883358389, 
    -0.252957824711157, 0.271147706620694, 0.758786052713791, 
    0.429980277282285, -1.25668004032177, -1.09964148009033, 
    -0.160141026502503, 1.48095713672304, 1.30501972014583, 
    0.218782414558194, -0.471601916857853, -0.625725287613248, 
    -0.615258535405783, 0.355717861463973, 0.800473211074895, 
    0.935515990711959, -1.27575910061116, -1.48973129204706, 
    -1.98562292218642, -1.34764611795554, -1.11981457956363, 
    -0.0197022724876694, 0.195861595186124, 0.177197541218423, 
    0.244010776760226, -0.112536110496104, -0.952137366757304, 
    -1.27931833031887, 0.0497472530465703, 0.0244060883323893, 
    0.295159969184828, 0.0377197990483502, 0.129256950369134, 
    -0.900976237265363, -0.895351975768577, -0.684493934429939, 
    -0.424621108373029, -1.01395227765853, -0.539876007811078, 
    -0.141049758213447, 0.433722142201032, 0.187323794994367, 
    -0.303147469487532, -0.156957683584098, 0.0684816039066893, 
    -0.90740159643206, -0.793332072142876, -0.151257887004097, 
    -0.29399109310404, -0.172226170110537, -0.369516751852768, 
    -0.0210472789602933, 0.605038023566022, 1.11605357935406, 
    0.576170741445847, -1.03345383230641, -1.0618940561678, 
    -0.492170934469112, 0.602538061286149, 0.634414196548279, 
    0.231306579382164, -1.01816960768405, -1.03176210928414, 
    -0.901290532414576, -0.119423187760646, 0.157831451317194, 
    0.778873089267988, -0.399785055784561, -1.20681476251668, 
    -1.0776700066971, -0.620184665252363, -0.340751699390656, 
    0.0452131701052272, 0.49446419922206, 0.153895944117544, 
    -0.115548964096295, -0.200424022163901, -0.26045242660754, 
    -1.30566355277927, 0.45275737987386, 0.23438606345092, 0.375299760443113, 
    0.0162419185779772, -0.10432845200727, -1.22768761416134, 
    -0.757639450421745, -0.703208071151673, -0.470986577792631, 
    -0.52640416107169, -0.42115275260409, -0.227717857836125, 
    0.656281463761728, 0.0344005407779013, -1.60104850344971, 
    -1.75505040207723, 0.0751461290971639, -0.514239084293804, 
    -0.756828865518928, -1.11097383806121, -0.840292058786569, 
    -0.156962800786649, -0.307962770010137, -0.0965530467744458, 
    0.807348434540271, 0.682292347509654, 0.322274923257466, 
    -0.891368331332227, 0.445932123882247, -0.149135092187249, 
    -0.0510917838392588, -0.203353934133554, -0.245174154591736, 
    -0.35714527277491, -0.362221587918334, 0.329101780303698, 
    0.0686550842139644, 0.120907432105035, 1.25975568540608, 
    -0.69277898805737, -0.862818841156376, -1.13100353339225, 
    -0.401491379040806, -1.00939114529177, -0.260251455541716, 
    -0.207951833112117, -0.213013311168919, -0.0869860584148618, 
    0.0928872312390272, 0.612393250017793, -0.742544267944845, 
    -0.387784493819368, 0.548516477128933, 0.590359074490312, 
    0.643909275536227, -0.225621026725475, -0.925425147674321, 
    -0.590258992683972, -0.667231772837886, -0.164289537491316, 
    -0.551622123422937, -0.724381075728058, -0.31895850960491, 
    0.267884407888292, -0.0305410911115445, -1.79393221733574, 
    -2.28708442248147, -0.241978178153626, -0.762573689820329, 
    -1.35233362088191, -1.23854556400912, -0.638973382585717, 
    -0.0909237645289496, 0.0306869455207037, 0.34744383356113, 
    0.552705243506924, -0.0417166399392244, 0.267842194033023, 
    0.125668620760009, 0.30489082015714, 0.443829134030476, 
    0.513376809693828, -0.0756163133027821, -0.324434442387633, 
    -0.557123169717282, 0.00413793178578814, 0.162852884867117, 
    0.134977272033723, 0.642867683691586, 1.25341770027775, 
    -0.427651947378043, -0.778827927955166, -1.00435984550685, 
    -0.416225176360833, -0.465277422803663, -0.19701922912573, 
    0.352376895513524, -0.356404359325184, -0.200044579512744, 
    -0.0151505388464912, -0.211317896844568, -1.73005708048632, 
    0.465229229017847, 0.849123794135647, 0.382952326241943, 
    0.294087551410085, 0.076548879839109, -0.0336092654249676, 
    -0.0948743971044586, -0.227580563287848, 0.235519596371949, 
    -1.44343509926526, -1.37361308178515, -0.506704922285603, 
    -0.920079739768793, -0.287460220079505, -0.852015798268693, 
    -0.191546807066329, 0.0894208762519799, -0.271754988807729, 
    -1.46866500116437, -1.16370386039682, -0.237947329697752, 
    0.378698029373212, 0.414326209486369, 0.705226788652333, 
    0.245701675573122, 0.0199886089428691, 0.458048887385929, 
    0.530497696233407, 0.511222602009087, 0.223255450464386, 
    0.828474311055056, 0.449726391574443, -0.0367700344659827, 
    -0.15009550943164, 0.471036032907479, 0.316667745400507, 
    -0.0199730066661141, 0.63235170112641, 1.17129706183464, 
    0.290617561934039, -0.568169111673633, -1.64296358342745, 
    -0.877180749230941, -0.096128991845208, -0.269125701100772, 
    0.284033124203118, -0.291644810001097, 0.126390508845855, 
    -0.155476536778685, -0.844688290487362, -2.03377814441576, 
    -0.393865604828063, 0.553958091276492, 0.770890455840298, 
    0.601915674482347, 1.63404953659299, 0.982408220655957, 
    -0.25421088488879, -0.91939961845299, -0.851299909669043, 
    -2.23120501739507, -1.95238608366608, -1.58727454181976, 
    -1.63099917965162, -2.35637150735302, -1.74003126361174, 
    -0.227349424432207, -0.30027147897151, 0.172787928977001, 
    -0.984149362036333, -1.02498244324422, -0.129488398129554, 
    0.373793269430105, 0.841325902269232, 0.551928557254029, 
    0.0502156850786006, 0.125154558441953, 0.603843568162645, 
    0.486696243633169, 1.15258214782752, 0.667758149952293, 0.47842081339887, 
    0.180924786642609, -0.0136995239220106, 0.382702043891436, 
    1.07410663389442, 0.370989206957861, 0.349522923277723, 
    0.374982449285408, -0.333907685503845, -0.154710642546845, 
    -0.494748156721103, -0.870717240365151, -0.780176777245156, 
    -0.179149985905549, 0.269152878683552, 0.136515977760179, 
    -0.297005758271758, 0.358795131793621, 1.296582478347, -1.55497285989826, 
    -2.10486755375098, -1.51118677716774, -0.20044537040909, 
    -0.0710292105573482, 0.507421578899709, 0.520634929258472, 
    0.7910251911761, 0.195461556345338, -0.447379896548332, 
    -0.838242834610639, -1.53841146727069, -1.24536293687359, 
    -1.71373862886061, -1.5317933822609, -1.75277986647193, 
    -2.73961179540246, -0.71300183585291, -0.985499860549055, 
    -0.0406774797158915, -0.107591297256397, -0.331347410062408, 
    -0.138507364314013, -0.227723687897079, -0.00446108028891334, 
    -0.0659203077026271, -0.398234826501729, 0.201824159231263, 
    0.531956893282466, 0.796284481907334, 1.19425728806836, 0.6202524389697, 
    -0.0445916519976652, -0.540791367394728, -0.813717330143753, 
    -0.702882185498042, -0.490372841290672, -1.00175569303159, 
    0.443248406729255, 0.815908395423368, -0.532188028230514, 
    -0.578298373153125, -1.00036451126321, -1.15355016919053, 
    -1.07911138138553, -1.27508529975694, -0.74152558692874, 
    -0.56463948322969, -0.334282200748315, 0.13664782352, -0.674377540879831, 
    -2.28881023973121, -2.00235133769641, -0.791394258600269, 
    -0.28479044163543, -0.480548715845366, 0.0475689931832068, 
    0.147664813600006, 0.0725140624067855, -0.466478350725126, 
    -0.212300070235942, -0.697071176776332, -1.10966000533127, 
    -0.442051448984793, -1.30564951363593, -0.810342494800178, 
    -0.395623614778176, -0.955393597681411, -0.643097520035831, 
    -1.31428921496701, 0.0834917724655337, -0.539766424986765, 
    0.0671511664453517, -0.265485762407329, -0.0697326287320532, 
    -0.0838035223783429, -0.464531422408556, -0.437704618369201, 
    0.0727507024491603, 0.710605577698726, 0.331301139003086, 
    0.32591974423783, -1.12097586029707, -0.273053202463811, 
    -0.0551655616109281, -0.982236954850757, -1.84541858623184, 
    -1.96576198087816, -0.831795363845953, -0.174114655410516, 
    0.00122415117677743, -0.614440714590581, -0.812259923615719, 
    -1.13725329030011, -1.41715737783805, -0.986003526629031, 
    -1.76739909535536, -0.768878133682684, -0.509066258941058, 
    -0.577029594202489, 0.299834561238977, -1.65977969929281, 
    -2.45517668912723, -2.0157478664397, -0.334965689861173, 
    0.32976501851901, -0.303378419346432, -0.374179764663625, 
    0.593057625932767, 0.552676330687172, -0.308192016429762, 
    -0.451063953180104, -1.12885063424817, -1.08290886616261, 
    -0.307829187919144, -1.41192745682116, -0.667710337221084, 
    -0.815301531369061, -0.618358044855412, -0.226663067094681, 
    -0.686822336705046, 0.136701044663345, -1.7878386637407, 
    -1.65418655107551, -1.00400864182574, -0.327364136375063, 
    0.458662066243845, -0.247513027943973, -0.502133590594829, 
    -0.615174186833842, -0.949821049194517, -0.619988790096109, 
    -0.793232701676732, -1.94162565676436, -0.455053925757829, 
    0.623531360071392, 0.280184346503982, -0.793082214010017, 
    -0.31269306503602, 0.394381274136002, -0.513147012471986, 
    -0.403656536888297, -1.27047214671052, -1.56175765390534, 
    -1.25913504501945, -1.75162881289612, -1.63810468624617, 
    -1.18541562914903, -0.949043932405602, -0.276002201630967, 
    0.437153139343605, 0.132097720756454, -1.94798205933302, 
    -2.0238916164205, -1.5934002684704, 0.120225462909271, 
    -0.0926917241149727, -0.144156066235954, -1.6127737520074, 
    0.294141849167957, -0.607788080679592, -0.27436553238104, 
    -1.06193475433627, -2.22445796302337, -1.39622249246134, 
    -1.0569541014378, -1.11459374293055, -0.528540447718551, 
    -0.793819614112286, -1.00392379397267, -0.343708452694864, 
    -0.21954216106268, 0.406872134152239, -1.64820986070221, 
    -2.64971646410827, -1.48390398558302, 0.0493944037541816, 
    1.40536744586554, 0.0120220326441389, -1.12138722552106, 
    -1.60643780447799, -1.19814036429432, -0.702034644299174, 
    -0.857942179265305, -1.32365231888561, -0.387122121136474, 
    1.08587557495039, 1.00606494359279, 1.06148102052154, 1.0981760068802, 
    0.365826306737302, 0.750942671993537, 0.575129667445635, 
    0.324708068932482, -0.325016134134013, -0.714717415831099, 
    -1.82127484184102, -1.0929362102851, -0.308531091837354, 
    -0.0660006352529097, 0.474931606038722, 0.0540180041177092, 
    -1.50704850282159, -1.08777715291388, -0.645088906420637, 
    -0.197184817298277, -0.360315713510042, -1.02556598770852, 
    -0.960173820963215, -0.448731758342165, 0.408197591619404, 
    -0.109378805546942, -0.805126650851395, -1.88788268142142, 
    -0.51989380788219, 0.177287279078926, -0.681781332382725, 
    -0.758521297208472, -0.966972481605932, -0.747513782127744, 
    -0.542942117556815, -0.755153075361217, -0.116691308187584, 
    -1.9873591363626, -2.59570651698335, -1.31024657142745, 
    -0.446249331677371, 0.986424606778273, 0.266660459513965, 
    -1.91460416555672, -2.59465197194773, -1.45731116455938, 
    -0.326729897087521, -0.272719647572299, -0.47850698907892, 
    0.389771969753783, 0.957164391812046, 0.39440094618314, 
    0.127084642169396, 0.156382072222918, 0.36637270549098, 0.54562782804783, 
    0.470398759600967, 0.865748320165451, 0.719647218690653, 
    -0.360764745869426, -0.380631783935117, 0.437079099426769, 
    0.654722052856561, -0.0603052558609729, 0.104547018605499, 
    -0.954553724615614, -0.456829989771306, -0.52031616679542, 
    -0.567111772211319, -0.76908919626459, -1.43475948284621, 
    -1.57167651050809, -0.823814812976575, -0.342697266385938, 
    -0.321172539677557, -0.925368068931069, -1.21109584558349, 
    0.442115618449574, 1.21535606461445, -0.163428161160626, 
    -1.00172830005033, -1.59483388618748, -1.21229640316271, 
    -1.52961743539819, -1.40143794378382, -1.49306323922048, 
    -2.00415384979074, -1.71811991511673, -1.0149880395904, 
    -1.29761315891057, -0.65377475751327, 0.0116118557487832, 
    -1.22194368782089, -3.24319056252059, -1.37271994564143, 
    -0.352873696707716, -0.972034322541866, -0.778028619372471, 
    -0.651736994697858, 2.01349837092393, 0.270449142873832, 
    1.42489702088529, -0.343331471269053, -1.5161127123518, 
    0.351114803435255, 1.36696787875276, -1.22873984780368, 
    0.0179764344156164, -0.412843815205135, 0.948927154708255, 
    -0.552856676872056, 0.563921251209787, -0.214433848736522, 
    0.149965389836799, -0.4810379008777, -1.59851484726036, 
    -0.443477430473658, -0.840648502499191, -0.355342737464809, 
    -1.02842947306478, -1.13754634069445, -1.02438254396912, 
    -1.64406135727506, -2.05549467500318, -0.573705100921229, 
    0.590596085958444, -0.220242305916285, -0.859148580638331, 
    0.799046926586571, 1.92903261228524, 0.72709170475084, -1.64464275661061, 
    -1.85707394210546, -2.23121092076915, -2.42696846593858, 
    -1.89250562604946, -2.05409428639169, -1.93529022267043, 
    -1.26594426419037, -0.514185754559162, -1.07344447264203, 
    -1.34841402471089, -1.31642097860388, -0.983203796522134, 
    -2.63870346735233, -0.810724897621881, 0.205607946724249, 
    -1.46010890027113, -0.850601760509763, -0.532903348119742, 
    -1.33945420919872, -2.86283122279451, -0.430938160407893, 
    0.317126454502619, 0.372027937851009, 0.359619991224882, 
    -0.308816914421426, -0.378794306892081, 0.540520524012917, 
    0.630569842954767, -0.422615075008559, -0.540188382560935, 
    0.325128546711176, -0.648870135169058, -1.56043073620898, 
    -1.08161428485501, -1.04191335563153, -0.629495106142635, 
    -0.577995447731325, -0.572495810508613, -0.696377967582262, 
    0.401916524157016, 0.231100857941886, -0.217120617775635, 
    -0.970993447866562, 0.705817673750753, 0.248162700918595, 
    -0.101413209280716, -1.81847127247529, -1.92610129099395, 
    -1.47342150421831, -1.70296691194386, -1.95808840758225, 
    -2.24574486228896, -1.65956059612232, -1.22789929168188, 
    -0.735889642982888, -0.707669619337166, -1.49581809762758, 
    -1.83365218126821, -1.41703202580998, -1.96686313679479, 
    -1.25172889099271, 0.106683592882821, -0.606464278816237, 
    0.231635947483768, -1.28376764837448, -1.4575105729704, 3.41473567507468, 
    -0.915936846790537, -0.48987515743006, 0.0399532492281418, 
    -0.244822511742797, -0.473394569341798, 2.14504405552535, 
    0.351316477126722, -0.232607288807187, 0.0930717857436527, 
    -0.588031364393604, -0.0236030513315377, -0.270729019136509, 
    -0.0268279350117417, -0.233965825852147, -0.0471809511843713, 
    0.658344782034677, 0.591016191315283, 0.777212865156578, 
    0.191487453821813, -1.1020910329381, -1.33420871973061, 
    -1.68056830817566, -1.45695670886262, -1.44851254876085, 
    -1.20375134666808, -1.76255896237713, -1.73323589192042, 
    -0.712079134676902, -0.882773505051433, -0.755266552602665, 
    -0.996429316288108, -1.88288864739772, -1.61872754372967, 
    -0.581785334168985, -0.233955867995834, 0.172603786547736, 
    0.44558307441946, 3.28976817135586, 1.24040095060379, 0.747451172819877, 
    0.295941110297546, -0.115309760526783, -0.131910117158176, 
    -0.458161909776535, -0.280632025399354, -0.460419943947974, 
    -0.205777461065306, 0.607019533666193, -0.314145725406161, 
    -1.3359927899275, -1.50444841969686, -0.776670707343432, 
    -1.77688862721831, -1.88888635065291, -1.41184701298521, 
    -1.5133451911544, -0.999166519908181, -1.22834461460649, 
    -1.6520903295985, -1.13557536061659, -1.05351741952074, 
    -0.488404843666297, -1.95062524989605, -2.07629002942856, 
    -1.54752730010108, -0.912192485396597, -0.200398897832104, 
    -0.491660551444504, -0.743860924890436, -0.743604668531983, 
    -0.808431418315521, -1.00088696901063, -1.89708753445718, 
    -2.59727027600959, -2.51096830896734, -1.44493357052367, 
    -0.866015496554779, -1.99811010717811, -2.0737467965526, 
    -1.89585453355699, -1.40679328793849, -1.24961321228135, 
    -1.01609739020069, -1.57938110664614, -1.52065500473067, 
    -0.811050613733495, -0.943159319350642, -1.04292440041319, 
    -1.51782112693093, -0.599637756181646, -0.561015997753707, 
    -1.03430420974173, -1.02871286417155, -1.51748448535881, 
    -1.72419859403014, -1.78650231728589, -1.54516301465612, 
    -2.36916962081839, -1.98849513704281, -1.18237184183756, 
    -1.6693746807523, -2.10249278597598, -1.91682213717213, -2.4627247592307, 
    -2.10570789970409, -1.31058729421026, -1.13611874269591, 
    -2.13899674669493, -2.26564923267109, -2.46564722943778, 
    -1.5259169045347, -0.768766317831897, -1.15237336200743, 
    -1.02722666535747, -1.282866472915, -2.30197393636899, -2.5639258986977, 
    -2.26551848261996, -1.08750907766259, -1.88692446229994, 
    -1.69407534797953, -1.10028434947748, -1.91947992823451, 
    -1.74049146817937, -2.70000059924847, -2.80394603044097, 
    -2.19005805691309, -1.48166893425608, -1.68578084478392, 
    -3.35552367958769, -3.58054451218028, -1.80418736926629, 
    -1.28999797203892, 0.337117599228485, -1.47219094834589, 
    -1.49273684690984, -0.87201557666738, -1.39302341644171, 
    -1.94469951319996, -2.11110057763049, -1.10610299700185, 
    -2.07186819239669, -1.76762804366188, -1.09128751068386, 
    -1.82813219470503, -2.22260712030433, -2.50325185224821, 
    -2.21503265506188, -1.91075402854103, -1.3338225244795, 
    -1.66772616269111, -3.07372488241988, -3.00921620923429, 
    -1.73823319573171, -1.25246899269776, -1.66080546550705, 
    -1.47300934328585, -0.81324809215257, -0.974482327945707, 
    -1.82851908064295, -1.57953781057436, -2.10536642968555, 
    -1.81046046481607, -1.40874028116846, -1.44912575759291, 
    -1.62351593478821, -2.48691853664435, -1.74507951280064, 
    -1.86934205617338, -2.21802851257663, -1.99469068283509, 
    -1.69298535708071, -0.747039894324608, -1.48403173842486, 
    -1.95606331075702, -2.28292750385635, -1.96797850045157, 
    -1.45422254485592, -2.46147871581049, -2.84833531523333, 
    -2.28933519132816, -1.86683122885542, -0.959693005916646, 
    -0.640446433837463, -0.92255085541157, -1.39370807628318, 
    -1.8058665714545, -2.04793161347421, -2.35367362191315, 
    -1.49617514467542, -1.4799836422095, -1.48281255205096, -1.8987654333238, 
    -2.33539215254463, -1.5952851205334, -3.13803164781149, 
    -4.07452026317494, -3.37679062763589, -1.02410828673196, 
    -0.40259325760144, 0.133153168237254, 0.59200312130363, 0.48576683690543, 
    -0.336766295047082, -0.517869930280574, -0.97123942056534, 
    -2.01093479355794, -1.45916652281733, -1.60737241091225, 
    -2.60196201150611, -1.55525442991625, -2.73064730063953, 
    -4.12046044337119, -3.33917179059943, -0.598265784828991, 
    -0.968140829486175, -0.266196276276931, 1.33489835622521, 
    -0.0231832922357178, -0.549622912968748, -0.211096177543899, 
    -2.25612764562725, -1.27926586889627, -0.493262216377794, 
    -2.35434265043228, -1.70241710059465, -2.36835873179472, 
    -3.88063916621177, -3.16796454369366, -1.92969787176665, 
    -1.68176822081317, -0.475086252368531, -0.0251903460658642, 
    0.41071930910173, 0.406632178586057, -1.37878967149967, 
    -0.581081169880235, -0.207449639171537, -1.77064750154888, 
    -1.55746702230976, -1.34916708256761, -2.32573777257786, 
    -1.70920396854349, -2.22681906027562, -1.62946235944332, 
    -0.490468220990388, -0.848841645680509, -1.03497163525802, 
    -0.0947969946391236, -0.297333976049852, -0.917861407115184, 
    -0.223440010816347, 0.733828272968537, 0.0679532470836364, 
    -0.169848383364268, -1.66929968349819, -1.10109221172294, 
    -0.558472879814498, -0.684702149500191, -0.946291719283847, 
    -0.620686378277195, -1.10147886920784, -0.907951838936083, 
    -0.0344649033335465, 0.643345131024526, -0.10973721371673, 
    -0.0206730833982416, -0.81324873787636, -0.581451365893551, 
    -0.890719418307477, 0.124234916425898, -0.298961354766893, 
    -1.08095958082685, -1.12877231354608, -0.251064769955032, 
    -0.93050792561018, -2.03604410568241, -0.349175032972067, 
    -0.370928541083835, 0.147587524796573, -0.237910167427322, 
    -1.22974977668099, -0.170826594729556, -0.878599379600424, 
    -0.916865994286771, -0.141037549393559, -0.96322311958827, 
    -2.69684762570519, -0.248950657719225, -0.452997103311761, 
    0.140867660628463, -0.410540083684694, -1.50599191395918, 
    -0.753457807994513, -0.885371895988558, -0.972678479810938, 
    -1.59317737813879, -2.13192541891404, -2.34294564625719, 
    -1.41326809868243, -1.52326995266649, -1.30362850276872, 
    -1.8019459062032, -2.01229438750314, -1.43956542396831, 
    -1.40751910100447, -1.50018427331941, -2.53181634259433, 
    -1.30887002380091, -1.59014246350432, -1.83570012715168, 
    -2.26731457995824, -2.24794749079547, -1.889361213558, 
    -0.318305227100706, -0.867097274422259, -0.432986971239346, 
    -1.23065605217402, -1.58009056929358, -1.74582508401137, 
    -1.63667231139216, -1.88498535621851, -2.27799570275991, 
    -0.253568495781824, -0.940916959001132, -0.289987643039482, 
    -0.230585382850723, -1.40434759588836, -2.30589844808472, 
    -2.24401975315022, -1.88288853966603, -1.68045199862216, 
    -0.691066493951968, -1.10391459693917, -1.85962390230955, 
    -0.812771588669094, -1.15976072325973, -1.2508865857981, 
    -1.85574648672434, -1.62662386661052, -1.58157052988631, 
    -1.7957846751738, -2.25226256075055, -0.840922993348601, 
    0.253857236984749, -0.930798813549143, -0.595654117905768, 
    -2.38951378328321, -0.0698255831869416, -2.46414006831358, 
    -5.91606840357928, -5.84135782038949, -5.24770246668172, -3.182288814572, 
    -2.04153396888525, -5.34278807943021, -1.35864296685977, 
    -8.08299460839507, -5.85960977303057, -4.42300047106117, 
    -9.4718766035028, -4.32973224234006, -0.317449997178728, 
    -3.32012332497331, -1.06866599687174, 0.920341717054125, 
    -2.79172025940768, -1.78829701917629, 1.37915953033347, 
    -6.85917661054006, -6.77767142840285, -6.27347296728553, 
    -4.56371207041299, -2.30402475707065, -0.63213485726984, 
    -2.14686678014273, -0.121393955335645, 1.16396039794594, 
    3.11880384654703, 18.8447289524061, 22.8377617668197, 25.964468031424, 
    23.5033845081495, 7.34263177040759, 7.5514219076986, 7.88592195962323, 
    11.8563840073456, 7.22052691173189, 2.42726427848297, -6.50073229714039, 
    -3.24279740026398, -2.42847896605257, -1.94449725369504, 
    -1.56898676335976, 4.26641745029215, 20.3375644295255, 8.35161650393662, 
    7.78073072614335, 5.71601207517345, 5.18986188552617, 4.79299439150367, 
    4.51863479140471, 4.86385602135329, 9.36662533492836, 7.67109175648031, 
    -0.324814220443918, -2.80763701704153, -5.36030320334026, 
    0.133202335536433, -0.495528498100741, -1.57148691109581, 
    -0.844696218019205, 0.745595429067167, 0.231121234801277, 
    0.187480467601828, -0.320313785400232, -0.319760914328029, 
    -0.117538090311884, -0.0563892812667444, -0.220706575443028, 
    0.454305730440847, 0.504641342044705, -1.29744673782288, 
    -0.309890105303472, 0.659687243900318, 0.728146863268511, 
    0.295172979283893, -0.263785374682932, -0.730565373494825, 
    0.39296661077143, 0.0913121595574973, -0.450348513085661, 
    -0.772644104530449, -0.751067606212414, 0.00689198791177681, 
    0.767853128764133, 1.55516563157792, 1.41085546152128, 2.4424623357238, 
    3.22045222689229, 2.62834546234848, 0.275591950552059, 0.679038778276646, 
    0.669240164150477, 0.552971599346415, 0.453170719945799, 
    0.540199279970972, 0.445194732395842, 0.548952033260344, 
    0.555816683935935, -0.432383627718362, -0.287842028226972, 
    -0.380823324522575, -1.39710636982374, -0.532047818039856, 
    -0.465479039110495, -0.271990075819031, 0.338302447411474, 
    -0.19401582978432, -0.182777878587732, -0.0251564929366754, 
    -1.09939333805414, -0.697534060006735, 0.0862336429264499, 
    0.581205078136326, 0.379551559886719, -0.347075565899688, 
    -0.462120100552488, -0.0467021383855748, -0.394026701282106, 
    -0.424259178408084, 0.0846985743862128, 0.224988245974829, 
    -1.65161539385713, -0.831974858825202, 0.21468346944201, 
    0.400633914818029, 1.00256526212868, -0.230319645328994, 
    -0.962465606820602, -0.154136874369244, 0.294318411529768, 
    -0.660091740161985, -0.951293093497618, -0.243603902385598, 
    0.428106782718141, -0.210703641078118, 0.406948283990292, 
    1.06926953065532, 2.00116269127751, 2.02233249092552, 1.07958619132628, 
    -0.479350066891513, 0.137736803079451, 0.683171033848318, 
    0.413206861337621, -0.122019373044928, -0.0294446849932939, 
    -0.0680228867976496, 0.0704093006170003, 0.268614346163609, 
    -0.276968253386922, -0.797464977634443, -1.32492021554297, 
    -0.938109232278763, -0.133916377283936, -0.476277605289948, 
    0.151389969056166, -1.00937337775433, -0.602915347757862, 
    0.191987250879277, 0.714640707624055, -0.220133944393437, 
    -1.19837933775985, -1.01489661472845, 0.21222290936163, 
    0.354796001566324, -0.442665649397203, -0.521283089661981, 
    -0.00215212093147343, -0.426910978528605, 0.0743344650176958, 
    0.154037963369098, -0.445365192440739, -1.58244491156144, 
    -0.797775881274365, 0.177018849646338, 0.353776645621067, 
    -0.390217529307466, -0.906135394243508, -1.13729261617287, 
    -1.15001809571237, -0.773370454934801, -0.841159671315346, 
    -0.453813642789163, 0.364906466074011, -0.318961770219746, 
    -1.24960079584205, -0.0587222580470703, 0.854638112940527, 
    0.499026330479801, 0.363090132473629, -0.679234339754795, 
    -0.330433200352012, -0.32883935206486, -0.0274661528369213, 
    -0.0964799805771621, -0.552147286236804, -0.0237154483914193, 
    -0.993608205173864, -0.911287742264397, -0.60735277198432, 
    -0.832078422847515, -1.59553441066299, -1.7170075612292, 
    -0.519945340426751, 0.109731063918241, 0.455104424481676, 
    -0.704801172137066, -1.17238750659978, -1.69102145411548, 
    -0.10661984784428, -0.0556394868516374, -0.850764279306917, 
    -1.51651819792525, -1.08392408042958, -0.410605686755039, 
    -0.14677967827434, -0.283946038613525, -0.00165112677112056, 
    -0.212777131928794, -0.606505650892002, 0.0242159278805598, 
    -0.234778199098344, -1.02411298596333, -1.08215235077265, 
    -0.707182964981463, 0.0842458290965986, -1.18933192027706, 
    -0.558177442495527, 0.582018637718429, -0.0174401182609918, 
    -1.30374891118058, -1.14175510968936, -0.502221934317659, 
    -0.269327924258151, 0.434209779395176, -0.34248153490108, 
    -0.931148163585593, 0.0265278645357947, 0.557416235642032, 
    0.945120036986178, 0.239525908884493, -0.312637796951947, 
    -0.790254657841407, -0.24048287268895, -0.530185114593458, 
    -0.363625511882018, 0.0724537513056855, 0.225315835130346, 
    -1.43376280187701, -1.7729458574801, -1.06931485534849, 
    -1.54436935136208, -2.13750541122125, -1.54442283003997, 
    -0.938109278464156, 0.332395580747922, 0.0329286172520149, 
    -0.0957473963801577, -1.82257545575254, -1.19178962727389, 
    -0.843528952355985, -0.714300771980945, -0.561510802516558, 
    -0.339864751169277, -0.0538097268112026, -0.852460055690383, 
    -0.15172849185765, -0.344056913773505, -0.409107265936424, 
    -0.783578160198388, -0.812077251608367, -0.0632467041668594, 
    -0.273720632893015, -0.83275934131839, -0.701603241629862, 
    -0.726740623501763, -0.877871937246968, -1.82592057617359, 
    -0.635321913452986, 0.069934411477468, -0.234750720446675, 
    -0.656151196607762, -0.875967370462085, -0.260211589337489, 
    0.339035814781461, 0.867353353280604, 0.0513826520993721, 
    -1.32675993783612, -1.01662731480936, -0.133391660131301, 
    1.5924819959368, 1.35963028270017, 0.329245512971603, -0.643287674347781, 
    -0.676682983774515, -0.583123914064756, 0.390083961274921, 
    0.869258193860984, 0.746976955412362, -1.58401182893479, 
    -1.61945516945413, -1.53212519561576, -1.56079959415058, 
    -1.25315422357803, -0.140648039204563, -0.101081561976035, 
    0.357199136068296, -0.155932101145071, -0.525057223444865, 
    -2.20234409814074, -1.28383423934564, 0.610719604781433, 
    0.922357879431724, 0.583274609516886, 0.533454842670258, 
    -0.0541113760541378, -0.997677028686415, -0.916133943571653, 
    -0.617586053169306, -0.306050071198691, -0.894524223322741, 
    -0.440820742307744, -0.0292312778468151, 0.511705317997357, 
    0.165214221240206, -0.0746674493356014, 0.259481789900384, 
    0.466953083199977, -0.845239939230376, -0.744154859557882, 
    -0.380697427722461, -0.404886681718688, -0.223829406979261, 
    -0.36772167898969, 0.144306441818598, 0.959411295993902, 
    1.32030406965734, 0.577561327294389, -1.01189734512574, 
    -0.849010957836964, -0.484758951339135, 0.710226529321574, 
    0.879063348759348, 0.333870323655896, -1.01661479923107, 
    -1.00344049760148, -0.839969575469555, 0.0462323608595261, 
    0.36589558807659, 0.917250700664769, -0.837685564347619, 
    -1.31108245317479, -1.18833704820668, -0.817681149923244, 
    -0.249884973573278, -0.01675505448123, -0.127476194748386, 
    0.117731820797369, -0.0427864345124496, -0.47522364039732, 
    -0.865038719769832, -1.40716065405702, 0.765562486012499, 
    0.543119969100099, 0.871859425800015, 0.00637314626272811, 
    -0.254108397399531, -1.52999748784323, -0.83467349552262, 
    -0.655703510868912, -0.4722895355789, -0.485531213221675, 
    -0.465249098075553, -0.149406527645306, 0.849394419994085, 
    0.200941762418489, -1.06770078125094, -0.82626664658533, 
    0.665655650977354, -0.389630884247238, -0.875790174944466, 
    -1.26978740143778, -1.04474205537773, -0.179968678753091, 
    -0.219262538481502, 0.0338493723674071, 1.2781679957994, 
    1.23188895189526, 0.528548543296514, -0.995575178188433, 
    0.40055027080832, -0.479312231318856, -0.0231886897715139, 
    -0.144517722865349, -0.140058597779404, -0.358985249986561, 
    -0.209012616297213, 0.409318664359257, -0.101990049624381, 
    0.116700498661171, 0.841715520185478, -0.406166002552344, 
    -0.752698476101505, -0.980244997922579, -0.708533820867792, 
    -0.844446166336734, -0.367265811840998, -0.641264423046279, 
    -0.178691257013552, 0.156970692997671, -0.233256324390974, 
    0.429597401143815, -0.458485810407536, -0.204423337148922, 
    0.379468176262785, 0.478645320874707, 0.648020536759919, 
    -0.238440278031069, -1.21749363506495, -0.746733915451072, 
    -0.787377178160895, -0.234414142750268, -0.672037634305216, 
    -0.770643315660613, -0.172428799745479, 0.436751942949196, 
    -0.184857280538666, -1.98710112774686, -1.76188880866209, 
    0.375804064477969, -0.620962638248215, -1.36909894335931, 
    -1.32932797855275, -0.623244690823332, 0.102373950374415, 
    0.0424678772887166, 0.182581234688719, 0.964537815497093, 
    0.511741137514772, 0.458987535996784, 0.13721813068813, 
    0.255063471281325, 0.347802208440102, 0.688178752437651, 
    -0.0941926950766137, -0.316317088563718, -0.359659464047648, 
    -0.00466161853335478, 0.191971527333408, 0.306309695468543, 
    0.700393079158341, 1.06836608735802, -0.341088824979243, 
    -0.645183177180177, -0.532437527545353, -0.603113597032854, 
    -0.917263269700532, -0.463465998937314, -0.258093587546915, 
    -0.37664153260049, 0.156376454723128, 0.212951201883516, 
    -0.318880662292576, -1.56138223446657, 0.399252349002772, 
    -0.103542494074604, -0.15269094516392, 0.705565353723845, 
    0.173348502564004, 0.0132915611348444, -0.293968241085105, 
    -0.370430338943355, 0.0333641659465167, -1.71846189741171, 
    -1.71180615505427, -0.603569268371555, -0.801692134411813, 
    -0.333957922632955, -1.40939766939487, -0.247436430406119, 
    0.331154385073855, -0.206213777289213, -1.53712480173621, 
    -1.27483091812265, -0.222781099778868, 0.423898714218023, 
    0.445570113379574, 0.70994840134857, 0.683452727242124, 
    0.296668018789878, 0.585090683707858, 0.713579893075353, 
    0.611953205503477, 0.314482179277698, 1.35848740791832, 0.48585453790305, 
    0.15144731179225, 0.0915311509547445, 0.319163055202938, 
    0.588715481251278, 0.585829589672207, 0.685052917489477, 
    1.24484444143674, -0.00140955183409286, -0.401248866170825, 
    -1.13000895929331, -0.96973690143578, -0.997181541583032, 
    -1.05068791469864, -0.482938089107083, -0.29467118605853, 
    0.669975994654131, 0.228303019839746, -0.808941530573755, 
    -1.55600976503519, -0.508587528439266, -0.0916759037615034, 
    0.0229792634561932, 0.821448233146018, 1.82515565252794, 
    0.78785874984594, -0.552718774810659, -1.12419830056107, 
    -0.936915785526309, -2.1777039747365, -2.35372876425957, 
    -1.76368701006298, -1.62793685165639, -2.11131098065867, 
    -1.6246902486626, -0.134331969757085, -0.123456639920825, 
    0.232757338168579, -0.947024907784675, -1.03574235264615, 
    -0.131561365799358, 0.488394861209684, 1.08711719760788, 
    0.708191916957168, 0.181029757063267, 0.262711856339011, 
    0.752434231447636, 0.6765610564528, 1.41082461638519, 1.05007024874407, 
    1.0139827824075, 0.562605524446953, 0.155545784404003, 0.740797784520666, 
    0.749984646391773, 0.705420067887159, 0.492547453375054, 
    0.0832827770968469, -0.5178325086891, -0.333463808266932, 
    -0.404474543641782, -0.375918744921373, -0.504692687409785, 
    -0.655385620317417, -0.192795767142111, -0.213480035897606, 
    0.240475839313983, 0.669469441749149, 1.85638866872471, 
    -0.769485682247577, -1.39202822280148, -0.932427191132872, 
    -0.671486575736546, -0.170805785343333, 0.208007159416104, 
    0.660645564575022, 0.715989215487456, 0.164738699820344, 
    -0.732696871553031, -1.12604688897718, -1.64864078337512, 
    -1.68537819453284, -1.97451397993767, -1.79543024487874, 
    -1.91745825449521, -2.75819610164409, -0.675446958610768, 
    -0.895876426147706, -0.098704231819422, -0.133929887450681, 
    -0.307677965506663, -0.256645288384054, -0.148820355322838, 
    0.133606183296702, 0.219291949258551, -0.0198951430876981, 
    0.43211034507737, 0.739073197058877, 0.733578584278769, 1.3727345945046, 
    0.711843338536067, 0.158901345996183, -0.510221574791334, 
    -0.571596090119115, -0.690431866551363, -0.655194923932811, 
    -0.836670398702468, 0.578777691548096, 0.907436167054647, 
    -0.536200370931672, -0.274548436527082, -0.676922049510038, 
    -0.481313948597153, -1.05324243896133, -1.26804181331256, 
    -0.372417846052024, -0.685071896923315, -0.0895289648036401, 
    0.519344399395383, -0.178539671915629, -1.45096157979293, 
    -1.65018312708257, -1.10372224315801, -0.234586604832794, 
    -0.426517124224617, -0.289668323874421, 0.166065243893705, 
    0.581212382566489, -0.789971687902851, -0.423004847279227, 
    -0.282674946206232, -1.35043820138967, -0.582446507041494, 
    -1.64066903155151, -1.06786727525668, -0.662838030135973, 
    -1.24476699645908, -0.853840330882534, -1.45857868849481, 
    -0.0234269810930687, -0.668444278901936, 0.138020527600542, 
    -0.505081582372333, -0.206394134236318, -0.228068761115714, 
    -0.470097725293095, -0.144739659837594, 0.13369417013263, 
    0.991994680938597, 0.861072355439552, 0.934542713487638, 
    -0.431584354174239, -0.40035396433181, -0.450308401303836, 
    -1.0208479932096, -1.64794922150064, -2.09843713927047, 
    -0.828317626735027, -0.101793995010571, 0.287827699438234, 
    -0.325452472596699, -0.385501815226679, -0.82302064369502, 
    -0.49998923793348, -1.14569176015471, -1.30426540421206, 
    -0.628767763747189, -0.713578813676334, -0.395612016432825, 
    0.768727581010231, -1.42683913128048, -2.02107920337747, 
    -1.53434124199889, -0.544497778925921, 0.203335652308372, 
    -0.34703450403903, -0.560291638707904, 0.293471789151987, 
    0.79258774862045, -0.335147237949363, -0.7159191234547, 
    -0.794499181862536, -1.32378590394511, -0.400990232520257, 
    -1.68528138231506, -0.963571903317431, -1.12159105287278, 
    -0.934500994503455, -0.411966928158161, -0.86057373766133, 
    -0.0142491705081227, -1.98666345064078, -1.72484575228208, 
    -1.12285580239601, -0.635708513319653, 0.117285781896479, 
    -0.600497022090107, -0.465208034960729, -0.12691452278685, 
    -0.557332566692454, 0.292229111002538, 0.366262636001546, 
    -1.02965259398681, -0.397650105597123, 0.401033651123548, 
    0.0787773658770297, -1.25088655681006, -0.708295673590018, 
    0.22684062319374, -0.0598821316122722, 0.00844435715937397, 
    -0.605599421539367, -0.97191227997329, -0.976582281266229, 
    -1.67807801400767, -0.76207232150713, -0.954057105758133, 
    -0.504706023294248, -0.0207494403395225, 0.272812590153193, 
    0.0779922204305983, -1.05363126682897, -1.54191348735525, 
    -1.24773357924449, 0.0158099949486346, -0.028082576256665, 
    -0.120020827167249, -1.00059065582821, -0.0404429820534702, 
    -0.467213779798445, -0.867336346003356, -1.33688583043225, 
    -2.25187836451129, -1.70708896299917, -1.1353632666924, 
    -1.46259539834359, -0.748250291463251, -1.17766096232192, 
    -1.32863556490701, -0.389356375081689, -0.317246158467706, 
    0.28316170204949, -1.66322762400713, -2.65907328714552, -1.555142500756, 
    -0.101887509367273, 1.2838170931196, -0.259069765926885, 
    -1.22391782667284, -1.2496937958573, -1.36548442921173, 
    -0.151329099656148, -0.38645368661459, -0.352379552405303, 
    0.607923731815622, 0.994921098824415, 1.07599576145236, 1.0137721905234, 
    0.918678078767671, 0.984603800475714, 0.309093171388617, 
    -1.49450172728686, -0.426722964978135, -0.271368446558728, 
    0.40464481501382, 0.0569855431295085, 0.208425460380459, 
    -0.0295492595264735, -0.927747305439497, -0.582573185119615, 
    -0.534933237588948, -0.532061076509009, -0.598084540312849, 
    -1.41897319967386, -1.3467895136657, -0.566408156509235, 
    0.173038953091922, -0.158777814115858, -1.78028273721559, 
    -1.93118951350606, -0.0578407364332278, 0.172048881701992, 
    -0.779569080902816, -1.07066577843268, -1.41827708002508, 
    -1.07622311003563, -0.673970645410926, -0.900886996822505, 
    -0.137998577651652, -1.94215767170869, -2.73310937552084, 
    -1.4362004941834, -0.657573056113527, 0.753714172590851, 
    0.0136135808356252, -1.96375273437889, -2.59864654057477, 
    -2.37330531395831, -0.368846413104653, -0.297363643069124, 
    -0.0439042984321736, 0.673464178235825, 0.710668260053846, 
    -0.0137337940599142, 1.34348638226708, 1.60000222531914, 
    0.639935048580953, 0.345620503765374, -0.0691726552290373, 
    0.238820272892494, 1.21682950806643, 0.317758210548016, 
    0.244204141432953, -0.736367054721239, -0.666973912649418, 
    -0.534915966287874, -0.072137757272297, -0.747526619723082, 
    -0.988788858658429, -1.81479281586296, -1.88387646401172, 
    -1.0303624650665, 0.102983429363279, 0.163609429030336, -1.0246609789174, 
    -1.6182038707868, 0.44486222937361, 1.3614755416013, -0.196498331394031, 
    -1.29371304394684, -1.9643664749681, -1.53086103281026, -1.5856097244051, 
    -1.39383562534223, -1.49287539877, -1.94668969651831, -1.70466487019758, 
    -0.952833675705484, -1.37774446573224, -1.19810808432247, 
    -0.339537117141178, -1.50022998005058, -3.98570040969422, 
    -2.02615210855947, -0.313445777057519, -1.23304310284752, 
    -0.942223099121891, 0.707024897654556, 0.955310308666988, 
    0.326562613237744, 0.506379471310492, 0.700624562031193, 
    0.246111182937527, -0.179082315254774, -1.71104242557189, 
    -0.958932070743315, -0.909969416508472, -0.0848159019987623, 
    -1.23265477083108, -1.33553944686815, -1.31294392223115, 
    -1.78727566857407, -2.0695745901367, -0.796761054665724, 
    0.405781445591495, -0.310530245117926, -1.29059576188857, 
    0.607693030620657, 1.94508072719137, 0.756924821088062, 
    -1.96709065485105, -2.21422527996013, -2.58878366869562, 
    -2.81854760050002, -2.09023148753078, -2.21277595835258, 
    -2.17204201403478, -1.34960557289351, -0.549646860241841, 
    -1.12076095469053, -1.55035367144293, -1.57423497042719, 
    -1.72088053994532, -2.79177424525774, -1.08876937212633, 
    0.496126643547985, -0.949766016854644, -0.616780182395649, 
    -1.6035910291161, -2.81182319753896, 0.442532905476503, 
    0.784169554557264, 0.670265461486803, -0.317250765466248, 
    -0.372253866383283, 0.349063011655949, -0.532358160348712, 
    -1.20700078812852, -0.647300924400185, -1.22510083828018, 
    -0.800653337529438, -0.719213824499221, -0.777629066838146, 
    -0.81332245005227, 0.354237518045672, -0.056210105274177, 
    0.081442952377806, -1.34241389616253, 0.223564274397692, 
    0.453201057019399, 0.136457434077784, -2.21108997945598, 
    -2.14412668460033, -1.70613751624495, -1.73535006235481, 
    -2.08710679479424, -2.43950619897781, -1.74491688675516, 
    -1.41833123427713, -0.674406305025204, -0.852782119494186, 
    -1.81027105485136, -2.12731876897664, -1.73813482349357, 
    -2.20238143068291, -1.62337659407937, 0.637620992473331, 
    -0.039644859908492, -0.572199189447267, -2.37790943481158, 
    -2.81182319753896, -0.401903222378488, 0.0974623937030072, 
    -0.0235697562838915, -0.193480103913179, 2.37115328362846, 
    0.657957399356358, 0.0876855060577542, 0.42667126988835, 
    -0.862623805544791, -0.171790095244111, -0.29989152080554, 
    -0.269216282697355, -0.495323190071284, -0.158717880627739, 
    0.336773918045585, 0.388721479716887, 0.483811045517832, 
    0.144223216065016, -1.0632338738337, -1.36611816933292, 
    -1.95406030299144, -1.77972952432939, -1.74472018421894, 
    -1.35342859420474, -1.84560191438384, -2.01864267525874, 
    -0.933349736580116, -1.30462229955308, -1.41089226457458, 
    -1.3950776954827, -2.13015385834338, -1.89133412483956, 
    -1.00393361632392, -0.377427757893285, -0.138207712191987, 
    1.13430801272911, 3.48291140334569, 1.64922042829879, 0.85945868539896, 
    0.6204869995817, -0.39834271570248, -0.259948762078315, 
    -0.659829867280806, -0.484896197107085, -0.509893285570895, 
    -0.126295266427143, 0.401417962818238, -0.645767614339214, 
    -1.58782504545711, -1.54106503716332, -0.634473782277749, 
    -1.85333896349936, -2.06404909236626, -1.57336581795906, 
    -1.71900038621922, -1.31359421452126, -1.4371102370221, -1.8866881892367, 
    -1.5854433752311, -1.73053214335144, -1.27124743572588, 
    -2.18741846218628, -2.26381040781408, -1.77064670704575, 
    -1.27074522507655, -0.456056938004741, -0.681903057522879, 
    -0.987141923429635, -1.01805063999948, -0.914375324753398, 
    -1.11361572456811, -1.98852901073264, -2.88548254103326, 
    -2.79803871642783, -1.30815935351848, -0.655651734909921, 
    -2.22393248954482, -2.21576356753126, -2.00603596069404, 
    -1.55916520726584, -1.57469727337083, -1.43063482675536, 
    -1.95662437883612, -2.00060356907455, -1.301374579724, -1.60743669891426, 
    -1.24219975798173, -1.46123455472555, -0.382721726665687, 
    -0.772723891138547, -1.23417468281245, -1.26485188462124, 
    -1.80497058865047, -1.85260546804516, -1.94614508889895, 
    -1.66211425668816, -2.60647025930977, -2.03523011442694, 
    -1.20856759993247, -1.56698050342455, -2.26229574649354, 
    -1.92934850166492, -2.10642732840944, -2.17357705545436, 
    -1.62935798521441, -1.38893148964018, -2.57031089092172, 
    -2.87482598978551, -2.96493539368584, -1.345238703834, 
    -0.0552846629085561, -1.1401558242136, -1.17155488973373, 
    -1.1398180771225, -2.61643568060482, -2.61028246899446, 
    -2.21904765336033, -1.23227275841661, -2.09871282272862, 
    -1.82810816501639, -1.33290160001381, -2.07514076346023, 
    -1.97839996784741, -2.79283613377381, -2.56012353813919, 
    -2.13000740973912, -1.34663390431551, -1.72595384429288, 
    -3.85219897451621, -3.94437676622354, -2.02379614663522, 
    -1.45873433758203, 1.14072156853383, -1.48501507482526, 
    -1.59331305595761, -0.77296057981056, -1.55295827163307, 
    -2.43394754891766, -2.2145441092048, -1.20815846811783, 
    -2.18940256181997, -1.8836942103774, -1.31163781235402, 
    -1.95972375534204, -2.28226517832931, -2.46110122972337, 
    -2.51115889303419, -2.29213223572479, -1.9638863136929, 
    -2.15061816785158, -3.39952914612048, -3.40721866595097, 
    -2.00037086790434, -1.3163008494008, -1.6582458341908, -1.25171633775299, 
    -0.62354038503956, -0.951545120889499, -2.15202086190749, 
    -1.6011198931202, -2.28829890383134, -1.87808552366312, 
    -1.24737254372548, -1.33207872350554, -1.59248117852993, 
    -2.24543911681728, -1.78784938838476, -1.98932085565063, 
    -2.73697835519558, -2.20710045178775, -1.97572436804933, 
    -0.939326843078887, -1.62429321415128, -1.81649514662447, 
    -2.19174905185118, -1.78299657346815, -1.48368117466235, 
    -2.78352081448571, -2.83214317730117, -2.15921568103156, 
    -1.60767086833455, -0.627141643439528, -0.413073898472156, 
    -0.764540630530632, -1.1107865803967, -1.72879790767197, 
    -2.03414003621306, -2.56397026929008, -1.60332376318985, 
    -1.36906191709682, -1.4320273951301, -1.948424109327, -2.50989780152714, 
    -1.8393667717786, -3.50785153257994, -4.03956027078782, 
    -3.28222758962689, -1.24254679919174, -0.301546841759208, 
    -0.0335379123606128, 0.504961808288886, 0.678451033397569, 
    -0.0758480678600293, -0.117110613594158, -0.615943441863708, 
    -2.12664685094849, -1.29597061261951, -1.30521405533839, 
    -2.69035053272471, -1.47810056071674, -2.95570975575402, 
    -4.23903240739921, -2.9676976538665, -0.751733888731625, 
    -1.01619373442495, -0.540428291750632, 1.26794623545892, 
    0.386154393464766, -0.184088769279915, 0.0918859234308167, 
    -1.98204926132131, -1.01194469367262, -0.343398285467105, 
    -2.42515151680553, -1.70242289160372, -2.27182879329269, 
    -3.84716440367228, -3.076821335228, -2.13091418521124, -1.80504101385962, 
    -0.530890781771385, 0.120793650214992, 0.553234689191715, 
    0.513312810468571, -1.25059770025099, -0.350415686786922, 
    -0.335342160803545, -1.7690031751241, -1.42856413492443, 
    -1.13897537638922, -2.13638850151523, -2.34424111316993, 
    -2.40436898030356, -1.68750722422415, -0.63296642892265, 
    -0.797900286614914, -0.723552533185989, 0.0231730076067382, 
    -0.489794779839405, -0.607884271190273, -0.0806680603998977, 
    1.49930846365409, 0.750356945712363, 0.0830242484437485, 
    -1.49177506097839, -0.632506150502699, -0.0933038441344314, 
    -0.434280600679888, -0.717656025857702, -0.712712752035003, 
    -1.3787187437013, -0.819686473248815, 0.158071592980948, 
    1.05231144230694, 0.350124664538463, 0.534428054909686, 
    -0.207323162977984, 0.244307268389035, -0.370135662639153, 
    0.119168612995981, -0.508715509722331, -1.09682726924244, 
    -1.40127512814321, -0.132218940995381, -0.702872899451115, 
    -1.44241239304574, -0.323726588498103, 0.220140737963539, 
    0.77552806223391, 0.560362463145943, -1.01811404327641, 
    -0.416399083752941, -0.934282326009588, -1.13250353307257, 
    -0.288644118137937, -0.778599612557787, -2.46590632731679, 
    -0.280970083489103, -0.367592400809915, 0.0970179547239525, 
    -0.218017858569723, -1.54228579201507, -0.736581624645387, 
    -0.99117279087217, -1.05558123713094, -1.74709072061395, 
    -2.05640148667163, -2.51788353032701, -1.66901379478296, 
    -1.52183086221691, -1.31477331860058, -1.93836100915279, 
    -2.09161191036371, -1.28598618250203, -1.84552749997561, 
    -1.8826821245933, -2.59604862472014, -1.77588788537894, 
    -1.88160545928802, -2.05570961548389, -2.60052073457212, 
    -2.30097568750238, -1.71539459551683, -0.880611761369847, 
    -1.71269897178979, -1.54851969071024, -1.4343087694599, 
    -2.04793657184811, -2.39783486499, -2.17622255589883, -2.17287612557712, 
    -2.35304635954199, -0.740576389450207, -2.21323187502485, 
    -2.30903888939586, -0.999553042930952, -2.24200326332847, 
    -2.96825399725926, -2.4331969272268, -2.0966703239479, -1.69259054336587, 
    -1.90659990881458, -2.45193702372426, -3.47175226673742, 
    -2.23942223217374, -1.60507945275446, -1.23518262553889, 
    -1.72325892177482, -1.4369889951343, -2.54271359433808, 
    -2.96147147613101, -3.28297170190339, -1.3653610870045, 
    0.0816145625067044, -2.19470036272942, -1.63801730459876, 
    -2.62326426703748, -0.201924417731298, -5.81242609591001, 
    -4.02157229791401, -3.32341523609815, -3.09213971470065, 
    -5.59089083570127, -0.448545724739821, -0.793030323019632, 
    -0.414668451145392, -0.435439976451916, 5.04731541430132, 
    4.8235817337364, 4.56132238870595, 4.73663595257108, 5.57738428804697, 
    3.36561073829228, 19.4449554844084, -0.187002193625411, 
    -2.04161896780595, -1.85205506023488, -0.982102427529803, 
    -0.349994125336757, 0.451998431456371, 1.10076013790817, 
    1.33279474632114, 9.0057056355819, -2.61639237349242, -3.13444542616892, 
    -8.9189467893886, -8.44857696393164, -5.01806325111794, 
    -1.19997236019487, 0.662045758608736, 3.33486417126799, 
    -11.0366152447575, -11.1626945438658, -11.8621381583019, 
    -12.1078372158841, -10.9996814728277, -0.828823234592517, 
    -1.20773416250039, -1.84681150342119, -4.80504294600139, 
    -21.8139000821211, -14.8040495607695, -9.17511320698878, 
    -4.36112777496263, -4.02554046491517, -0.801441055812546, 
    -1.41980716137903, -0.945347198533593, -0.630786781707181, 
    0.0718167023083555, -0.53345478375523, 0.503445288184047, 
    0.398592217331217, -0.235119556801038, 0.872453599609292, 
    -2.15960078025205, -1.20336247731611, -0.268529825582066, 
    -0.872014819371469, -0.982275117220301, -3.35068542478096, 
    -1.44612716537114, 0.55871129901878, 0.145062566914762, 
    -1.52797061116967, -1.34582788033664, 0.591677482662437, 
    -3.30974623090603, 1.11664594783874, 0.158522198694742, 
    -0.574705108583876, -0.369671510814658, -1.61906763748206, 
    0.705230187898934, -0.111598439583827, -1.69812577792521, 
    0.0128563349579391, -1.00512365037197, -0.967165617424863, 
    -0.404194317574386, -0.854945292001664, -1.10635543119082, 
    -0.148956160516349, -1.52438657775102, -1.43421004803318, 
    -0.829718843425795, 0.0179400340865263, -1.05958566312239, 
    -2.03927659055139, -0.602210910611307, -1.93462649085661, 
    -1.23061159978322, -0.518549247596724, -0.545232047180383, 
    -1.09931648027544, -2.68257834485517, -0.496042804261627, 
    2.07751107947197, -1.33287225428627, -0.433995245231366, 
    -0.517310484880765, -2.30247228651369, -1.39354235997349, 
    -1.28823672824546, -0.151457486134418, 1.39554128217568, 
    0.0313661573045479, -0.205127450059631, -0.470694414425595, 
    -3.08373423428528, 1.19705570824633, -1.01499362023814, 
    0.804834975232859, -0.517552184430607, 0.574736024497588, 
    1.22602906175329, -0.840419524634792, 0.245505422184612, 
    -1.2677931069135, 0.710516193379931, 0.155817123408476, 1.15055109411787, 
    -0.873617639159556, -0.145270185019963, 2.06978956218542, 
    -0.019124475410192, -0.903701369751821, 0.615869019464338, 
    1.48989882021212, 0.950302545128613, 1.32178866552688, 
    -0.144175046479919, -0.370067729951513, 0.0710945184936043, 
    2.37381859902792, -0.756213311603862, 0.17418122983263, 
    0.309429541092217, 1.84966732116429, 1.0525689869113, 1.94947327753612, 
    -1.94915741849222, -0.846708716989854, 0.0455535916987701, 
    0.595754228793915, 2.0828903648882, -0.583704125484855, 1.30328899246574, 
    0.0299158670543323, -0.0326634181114963, 0.707331909004227, 
    2.54986381538891, -2.11725342812485, -0.0393913327636289, 
    -0.0483661109750178, 0.387734186192173, 1.4564320164458, 
    -0.262619644367142, 1.84599075548674, 0.0214399211960939, 
    -3.57975142652727, -1.23737866897257, 0.0249304950804358, 
    2.37777028950745, -2.1374611391392, 1.28166502601877, 
    -0.0149737612833697, -0.270142855866366, 0.840487564151, 
    -0.267151647718916, 2.10171149902047, -0.383272368610989, 
    -2.94503519864215, -0.89317335574423, -0.557180236243496, 
    1.40201919422657, -1.9871143246418, 1.91416636298107, -0.428269572027941, 
    -2.43127800996426, -0.765933946716266, 0.141786081265304, 
    -0.874352699919472, 1.86248575228524, -1.11383592606764, 
    -2.67345411106953, 0.381489428876503, -0.444936376355186, 
    0.433565100575985, -1.09085517868008, 1.82451818033284, 
    -1.40223407038688, -1.33806871505031, -1.22319804521434, 
    -0.352510041427016, -1.65316688557887, 0.80622692519898, 
    -0.660112388010552, -2.13396874390777, 1.37274802423669, 
    0.000512843896697396, 0.177595164352071, -0.398190373279492, 
    -0.734708470582987, 1.10918050682736, -2.05481655859399, 
    -0.716118354920332, -1.20091278867453, -0.322070830872671, 
    -1.64624738964693, -0.190671784697929, 0.476495597626712, 
    -0.77777878465987, 1.41968625759284, 0.525817793096728, 
    0.0210517558459078, -0.747407193133334, -1.48947831155387, 
    -0.000526385864965673, -1.21542115805009, 0.266802756229283, 
    -0.781192725313287, -0.187507059020582, 0.565762995528478, 
    -0.307129005957357, -1.06392916801169, 1.14379889326943, 
    -0.164228228955032, 0.546172846180978, 0.282632160616684, 
    -0.854752994133866, -0.558610950516986, -2.04582795001633, 
    -0.725072377942261, 0.0279932057597548, 1.44105211598808, 
    -0.189926282402052, -0.592250605375011, 1.17476174405408, 
    0.634897339338561, -1.09169677387277, 0.978590817824296, 
    -0.837806268261344, -0.461888454550412, 0.698158654555083, 
    -1.21538691373958, -0.0418838704661376, -0.670150674532069, 
    -1.04238827662333, -1.20605724321911, 0.382070215758015, 
    1.31633936397384, 0.0904991424647894, -1.15772553683386, 
    0.661341430615518, 0.131879934093003, -0.676690174479427, 
    0.413177733561362, -1.46956391895344, -1.03688203825409, 
    1.87820373887361, -0.905355387866646, -0.0129179260081311, 
    0.529737322273157, 0.44714007697524, -1.1028831978398, 
    -0.211888145974513, 0.278767847971947, -0.151963640613674, 
    -1.31256090525994, 0.74921218555478, -0.437032293334659, 
    -0.252296997402192, -1.36685244328342, -0.251915855779656, 
    -0.78550439233836, -1.12082765172015, 1.62932880437024, 
    -0.203190613880301, -0.276963939843693, 0.51111801370222, 
    0.655220648017654, -0.981212941755437, -0.913692977135674, 
    -0.179785934764953, -1.07880266566753, -1.24709596960253, 
    1.73924140965262, -0.489885020971625, -0.0267981282384228, 
    -0.032885938244058, -0.543052904748403, 0.567105614119541, 
    -0.920718698200523, 0.024812724448417, 0.0419707907520314, 
    -0.853333827404019, 0.234843003906009, -0.0528426692438466, 
    -0.992380398310858, -0.63722044107027, -1.67542082124696, 
    -0.0354977693590053, -1.88017689219569, -0.947456851176004, 
    1.37951252557445, 0.020809522661662, -0.224872290651412, 
    -0.721660766245181, -0.835166174855578, 0.975033830035552, 
    -1.11589169375621, -0.898066707875462, -0.514134415468587, 
    -1.33274797718406, 0.357510728877734, -0.532268113384858, 
    -0.972469985765568, -0.157406382663455, -1.96922360718204, 
    -0.0514798440574241, -1.73815204918791, -0.583316023550001, 
    -0.504882424882463, 0.433809383624052, -1.06073825943713, 
    -1.88906011701424, -1.44812318730069, 0.209709815202865, 
    -1.51784842201058, 0.334993862724211, -0.643443255603553, 
    -1.27517290460286, -0.807583209610549, 0.2169542094607, 
    -0.204263567067146, -1.2008399936169, -1.86048727193592, 
    -1.92280436866797, -0.466553301445848, -1.33640803741125, 
    -0.626456694562098, -1.55726135668502, 0.429178623685002, 
    -1.92032951751821, -1.98754587798403, -2.05437611027217, 
    -0.547520116587234, -1.52400569552052, -0.191003642592391, 
    -0.45959997282925, -1.39947149471144, 0.431219919063978, 
    -0.704197619359222, 0.485531863265058, -2.21093739091942, 
    -3.11155603244859, -1.92027529079187, -0.828532663371816, 
    -0.89770848850868, 1.20812573660057, -1.02335174196512, -1.105403882886, 
    0.174223294550846, -1.28261534294428, -0.996355066318499, 
    -2.00200086292136, -0.435724669842649, -1.63540318021864, 
    -2.06603232121819, -1.04672382479447, -1.14378023028444, 
    0.814732507051625, -1.30196341846767, 0.658155529659638, 
    -3.30450993419358, -2.58949708092517, -2.06567760002695, 
    -0.838816747585158, -0.258078118325055, 0.229825982246078, 
    -1.01802119443571, -0.6024780437065, 0.16007872457211, 0.654303468956027, 
    -0.364910798263184, -1.68480544034266, 0.267672038628067, 
    -2.66419491088499, -2.91016435349258, -1.46511762010956, 
    -0.747799589089873, 1.78080558288307, 0.0158921108144749, 
    -1.01928570219051, 0.598274831314932, -2.81943523216899, 
    -0.773846343516325, -2.12753166276758, -0.81785892026896, 
    0.0220302980309102, -1.19416761436718, -0.809920448834315, 
    -0.986538961846675, -0.0185948759441698, 1.48975818225486, 
    -0.430573165579, -1.02231180761064, 0.363245540060508, -4.06394738287696, 
    -2.21947690314366, -1.27720093645711, -0.15877043519009, 
    0.273851180810694, -0.837750385023289, -0.569873831139969, 
    1.02350983319692, -0.569558809533111, 0.139882915392344, 
    -2.45131982225313, -0.671373997399502, -0.963792121262409, 
    -1.72653643238774, -0.222359034051491, -1.35017006191908, 
    -0.590978061501097, 0.877694911741468, 0.547295853693961, 
    -0.75053080950726, 0.00689568015230565, -0.0682071655128444, 
    -4.06277102383625, -0.101124145702933, -1.31381929281156, 
    0.353415022875863, -1.00104131408734, -1.00263882548033, 
    -0.51142179469729, 1.01978222105681, 0.922677325723147, 
    -0.102225351095069, -2.48941365057671, -0.830531326604544, 
    -2.91160134647101, -1.34365023525724, 0.31045362095886, 
    -1.46712562703325, -0.749543586899589, -0.573879632278296, 
    -1.51967922240334, -1.22485682419456, 1.19344081519398, 
    0.293280043254115, -2.12219437826501, 0.995992433728947, 
    -1.12610479917733, 0.107710445677628, -1.33087623703137, 
    0.177711429598137, -0.452959701792864, -0.120087543869342, 
    -1.11043099317105, 0.220109193108971, -0.809075863875942, 
    -2.03791324043762, -1.98528757127455, -3.78364331221066, 
    0.30967411609015, 0.145535245268257, -1.80792549026768, 
    -0.218285418519279, -1.8810167021965, -2.90803189356513, 
    -0.903197214607098, 1.74407615573104, 0.663256238116985, 
    -0.347814817753487, 0.60092710361612, -1.20341919291632, 
    -1.19375201326753, -1.05422442062959, 1.6117599322182, 
    -0.984737436065741, -1.01192020827814, -1.75594919823163, 
    -2.22280346251803, -1.95815045614043, -1.5008424629349, 
    -2.09748354355156, -2.24489319413995, 1.74571207256683, 
    -0.0149899108935762, -1.57884370200756, 0.162338286580193, 
    -1.58528048401281, -1.38078901560408, -0.220940403855798, 
    1.71645236346865, -0.399933120710486, -3.38560735347821, 
    -0.0928441653172594, -0.443110682608605, -1.86035105400781, 
    -1.80066393258019, -0.113848486029616, 1.88270339280773, 
    -1.89451590275858, -0.951720397759301, -2.30105625604912, 
    -4.15874009987425, -2.35377627125043, -0.845623194945514, 
    -1.5882055474208, -0.075276002681636, 2.36327826100872, 
    -0.685669836664766, -1.15981356351, -0.371414198451364, 
    -0.558107393467758, 1.214689701182, -0.827136766352988, 1.19554832755781, 
    -1.5316558231184, -2.42253412364202, -1.50661249052669, 
    -2.31688964872631, -0.655816652925934, -0.439801776036869, 
    1.36341157674059, 1.34392906737813, -1.66764393884607, 
    -0.885945511790439, -1.47617643779079, -2.79319737143996, 
    -1.90443431665642, -0.0078250998005177, -2.41483613391753, 
    -3.58628763305101, 0.906868829153129, 2.29353421521109, 
    -1.90832146003406, -0.602273368722921, -0.526777633102408, 
    0.278057717393006, 2.39296174822626, -2.45440842905026, 
    0.0548810500882475, -1.73567332098834, -1.49383828996671, 
    -2.66394996443957, -3.94386373457755, 0.669972303011798, 
    1.28222364775462, 2.69865487547224, -0.500963080496257, 
    -0.648542800223783, -1.26768946653384, -0.104386534704403, 
    0.256235866951811, -1.94733569068448, 0.388926212608167, 
    -2.93138238687613, -2.60618664028895, 1.21751515835453, 
    0.0683746901468094, -2.94340348172779, 1.52280071249564, 
    0.402883215948449, 1.00175675490719, 1.79284158858852, -3.03451623430015, 
    -1.03045164696505, -2.37003496850454, -0.716392124514495, 
    -1.864310922507, -4.1483867411901, -0.370490126568424, -3.02676074435718, 
    1.37370138116231, 3.36959472986127, -2.83290321876037, 0.362342167843682, 
    -1.34581243857171, 0.179379383573167, 1.87615727211375, 
    -2.74654723647668, -0.339405492742491, -2.45932538673513, 
    -1.33967434070716, 1.79008413565255, -3.0305571322609, -2.53507044917318, 
    3.17832045069604, 1.15699548100957, 1.16837450414743, -0.524967267714781, 
    -1.6407313164196, -1.91605621521781, -3.10638874649026, 
    -0.481863305123839, -0.0719425941264382, -3.56920836499679, 
    -1.39166619315188, -2.68113411307792, 1.07681759884039, 2.56076102406469, 
    -4.02262915308334, 2.05960483245008, -1.01975106691561, 
    0.0986153121668368, 1.47522599826979, -3.21582613685109, 
    -1.60247725646461, -2.71109636193214, -0.571810617210836, 
    1.81429816098352, -4.30256984580051, -0.37104496032622, 2.07025922522325, 
    -2.36111468140239, 0.612660206795792, 0.648586563973103, 
    -3.3009451638052, -0.288286296961572, -2.34852734504719, 
    -3.27310013281294, -1.66868071438478, 1.0463336957011, -3.15036129236602, 
    -0.724591353844108, -2.17522543641361, 0.943262761639789, 
    0.244378680788191, -3.30308117149574, 3.48512400812733, 
    -0.466334160384932, -0.178722437026558, -0.194947901037941, 
    -1.83021060264658, -2.877131380304, -3.54208313844469, 
    -0.888800295896039, 1.0204033958201, -4.00292642810441, 2.04795867344475, 
    0.400475270890688, -2.31253216403532, -0.315772845812757, 
    0.711935930186276, -5.0671822169556, -0.029452733468853, 
    -2.10121170782533, -3.1471916070393, -1.85633000523601, 
    0.931385210717704, -2.98935145199532, -0.0408122291283401, 
    -1.44872527903559, 0.61318810163586, -1.76267368175157, 
    -0.819431018960779, 2.97518906606179, -0.96696792014821, 
    -0.440998534899772, -1.17268180690788, -2.31179872076318, 
    -0.278503445004128, -3.65588807178943, -4.25884761262462, 
    -2.82751651055169, 0.104649676141818, -3.47875468630108, 
    2.09284834778357, 0.980180619344909, -1.99948252675746, 
    -1.01140038320352, -0.099029144737969, -5.22869003991181, 
    0.273629426901892, -1.37939215130911, -2.17402069842908, 
    -1.22853009065231, -0.0249708316627406, -1.82008016561436, 
    -0.572020842850768, -1.34323459065225, 0.011229752786851, 
    -2.33252883230332, 1.84851452923055, 1.594532452466, -1.06433072427135, 
    -0.959454884367075, -1.03462429043842, -4.30898533394693, 
    -0.0395015068721002, -3.67694032290719, -4.47496308332037, 
    -4.33746327067385, -0.179737337704994, -3.22082412357909, 
    0.134111458171161, 2.33345039085126, -1.52093204722126, 
    -1.39457183756232, -1.47421915813159, -3.33838116514373, 
    0.638409361014559, -0.937034898008889, -0.247873350259074, 
    -0.975810395411118, -1.48485325565325, -1.02862042586814, 
    -0.632763795025383, -2.20052054809305, -2.70287971689601, 
    -0.721833886867389, -1.93247275766847, 2.36016955486672, 
    1.74786739477825, -1.0954083072824, -1.1305659692716, -0.863392254057475, 
    -5.46526966881754, -0.0524111137058945, -2.75233640187939, 
    -3.14313204642587, -4.07120380833398, -0.235094205973205, 
    -2.45879294362638, -1.39660841092989, 2.2377820504366, -1.35579731938344, 
    -1.41978466828432, -1.83877310244299, -0.893194748823275, 
    0.402902709386991, -0.994174780442899, -0.135376135910418, 
    -0.389920617412581, -1.52633198494628, -2.26372973044992, 
    -0.324410511501224, -3.83541366364809, -3.92448236918169, 
    -0.747722857002293, -1.55692805317392, 0.816938202423978, 
    2.98859251493497, -1.08965917414887, -1.11374416415522, 
    -1.88391220909416, -4.79892103224257, 0.293200817742195, 
    -1.53963996259505, -1.55971677258997, -0.985506387972017, 
    -3.8165535118596, 0.088026012020017, -1.7516093828195, -1.65948381035935, 
    0.220603275257363, -1.94418168472423, -1.83341721308829, 
    -1.26197216895333, 0.228183229791111, -0.202349648714897, 
    -1.67555439882074, -0.634655384999889, 0.00150742737968015, 
    -1.2429612599528, -3.90568376162425, -0.193040390598888, 
    -3.46982292980818, -3.41900771446052, -0.288184633442529, 
    -1.43615077614008, -0.278050345874872, 3.19774262950611, 
    -0.957952802116005, -1.47064094482012, -2.27988727522624, 
    -3.4618066437528, 0.365428929742138, -1.64140517331228, 
    -1.65698159854086, 0.229619254230114, -3.72768622252553, 
    0.465556731724421, -1.3572319774801, -1.68156427378949, 
    -2.54897741221771, -2.50638952488308, -1.98777630954787, 
    -1.14848500124008, -0.341532224809673, -0.159107543136221, 
    -2.02626219960606, -0.146424098633628, 0.295221139305867, 
    -1.4523611001054, -4.64889297508078, 0.31718395105207, -1.6975295680229, 
    -1.32585062363817, -2.25607288035677, 0.147446794532767, 
    -1.56970407569682, -0.130374171395098, 1.35703928044355, 
    -1.27654859504967, -2.65037351231771, -1.56896130863451, 
    -2.34992310995135, -0.615248259208313, -2.70471213702398, 
    -1.68887416997713, 0.45587884155654, -2.36326834693595, 
    -0.17594659601945, -0.903941165254755, -1.49262891962239, 
    -3.53243465343236, -1.97171984954866, -1.22817404120573, 
    -1.46516322093179, 0.0175580931644529, -0.021144139039371, 
    -1.70788170800668, -0.296327312150021, -1.90330212436572, 
    -4.23070430380171, 0.787425130448065, -1.27150870374872, 
    -0.299442694793606, -2.23235745715393, 0.518118709767187, 
    -0.976049124873728, -0.379550072707656, -1.42724150441851, 
    -2.25066445728618, -3.17419420210508, -1.23781537585881, 
    -1.82248747455431, -1.50832178059297, -3.29431019114212, 
    -1.64697348133128, -0.320703308583195, -1.51243381569545, 
    -1.93002542661699, -0.429228497954687, -1.72759265410537, 
    -0.925832655764159, -2.30954589692761, -0.927096384141193, 
    0.0603038744159547, -1.5952437706385, 0.29454860026129, 
    -1.11709848451752, -1.90512123930674, -1.56833728055142, 
    -1.80138373324685, -3.39574075683388, -0.0720936166779595, 
    -1.77899054919314, -0.566582635256805, -1.87499210100554, 
    -0.417963088826002, -0.385370251390438, -0.687444389420552, 
    -2.80745992299032, -2.93907146965919, -2.31625998968159, 
    -1.29399003896478, -0.860065841337666, -1.25686653335313, 
    -2.92411152095216, -1.22921266878121, -1.92966670313868, 
    -2.30943992966817, -0.0620137076610051, -1.37303112642212, 
    -0.6798696360332, -1.59238735170356, -0.680126846287107, 
    -0.0428383613355475, -0.852179014725437, -0.435550083992736, 
    -1.93173509859587, -3.13510000342351, -2.3032548365984, 
    -1.34436047365337, -2.68318490292914, -1.42183488639112, 
    -2.75781875018791, -1.20315600951501, -1.70254568990851, 
    -1.95776083171899, -0.455443896474001, -1.89991443697047, 
    -0.818614170851758, -2.38008490399725, -2.58364482358603, 
    -1.13621949466292, -1.15356075008426, -0.246317082523297, 
    -1.56214178241268, -2.77189026871712, -1.07989630456348, 
    -2.71576017303369, -2.37784740390093, -0.529536138170007, 
    -1.54935334029391, 0.579661162087237, -1.71604299338729, 
    -0.941785134496493, -0.663851852117858, -0.203931792063594, 
    -1.43343772360831, -1.65061750160009, -4.22586924434808, 
    -2.36419261532508, -0.313181564301971, -1.59091099571082, 
    -1.28512487312241, -3.22078985278726, -1.82801321476327, 
    -2.57147990201807, -2.05126375413034, -1.12209216319555, 
    -1.99851298316591, -0.930497171447278, -2.22556856664154, 
    -1.32589397995117, -0.628643371526058, -0.546996100362935, 
    -1.02875195481132, -1.78193765071123, -3.55881862674223, 
    -0.46970745194083, -2.18435616508889, -3.04700611729286, 
    -1.35844590182899, -2.29927610375816, -1.42910335615007, 
    -1.69534700713667, -1.75855160121818, 0.0701497451770103, 
    -1.5769282611271, -2.19471424627873, -1.06002863247531, 
    -3.75746936402222, -1.63372859938459, -0.0886651551370173, 
    -0.866559188999251, -0.643548092065505, -3.16866399819029, 
    -2.10789923042536, -3.46857602851781, -1.92349849637429, 
    -1.50030414105054, -1.89435649254601, -2.4337844631159, 
    -0.807673419984188, -0.618206884900853, -0.136035700900575, 
    -1.54733784732968, -4.35043427302761, -0.0546679246369544, 
    -0.465063378879042, -3.2243149470919, -1.45740659202469, 
    -2.80004486539315, -1.19359897359074, -2.9683512213834, -1.8821263310106, 
    0.0497182602424704, -1.82525631358528, -1.93528900535685, 
    -1.48420561688013, -1.79087597245483, -0.641169400824774, 
    -0.186367195325107, -1.97801280722148, -0.309359692482308, 
    -2.86021475451915, -0.626145711717421, -2.21183638919487, 
    -1.31741021880761, -2.31667260548622, -1.23358502690408, 
    -1.70578358730481, 0.336064836454936, -1.40448301071627, 
    -1.20215907089718, -3.86072738449997, 0.042591785426864, 
    -0.19225203870461, -3.097609412425, -0.46703224966641, -2.76668135984053, 
    -1.42959307924764, -3.43642800179354, -1.72703806621333, 
    -0.113259942264376, -2.10532648718068, -2.07549154546084, 
    -0.675371780018518, 0.112174434142156, -0.301608726839331, 
    -0.352707183084378, -2.26156237734913, 0.443408238245796, 
    0.311785466379595, -1.33178222709391, -2.64757319169367, 
    -0.627604421240157, -2.3861509803935, 0.949519802153586, 
    -0.917609862412149, -1.57201156253756, -2.11236655309854, 
    0.73143566206654, -1.72308005113855, -2.96712450912602, 
    0.698744222487523, -2.26608095577694, 0.0453951499972904, 
    -1.08723563740776, -0.616951928777546, -2.86865555954285, 
    -1.9871758212649, -1.23198987170216, -0.0426979638678941, 
    -1.59202951025395, -0.849179020799107, -2.0384241442223, 
    1.35383476331414, 0.372532802759021, -1.16485405234294, 
    -2.42026163989037, -0.713284752030874, -1.7881688205009, 
    1.02251552935365, -1.4305253032263, -2.12159705923559, -1.18821324555837, 
    -2.05274171608966, 0.957240643744637, -1.62439323844321, 
    1.66272922656205, 1.95271441784862, -1.02590444735246, -3.29209453235342, 
    -2.02809798994846, -1.35349600310736, 0.431854181449996, 
    -0.275325157420876, -1.73425623474151, -2.35407170303324, 
    -1.36206734946192, 0.340953383701019, -1.85868007607853, 
    0.659163773434046, -0.374326417986438, 0.119780906088988, 
    -2.50141802942273, -2.08489966172792, -1.48328678692248, 
    -0.438327064871238, -1.45503015818914, -0.091965435967338, 
    -1.54301652396925, 1.72315182914627, -0.948150166254774, 
    -2.33511301344465, -0.858183379894096, -0.59167827946886, 
    0.639406499110166, -0.535426889334825, -2.84239041371001, 
    -2.77442787464832, -1.44033004326228, 1.56214296805605, 
    -1.46172403284955, 0.109216017126446, -0.611435670348453, 
    -3.11481044426849, -2.10929301623842, -1.26932473521283, 
    0.553866416313525, 0.788454051601646, -1.81123063647397, 
    -1.71875844771804, 0.00342401653588981, -0.167050601663248, 
    -0.649677279245477, 0.881233559658374, -0.531340795432135, 
    -0.497736681335252, -1.72002703992886, -2.81645308757261, 
    -2.61481287188871, 0.00297520170277343, -0.557899634727981, 
    0.987290653809811, -1.41204637090047, -0.642709722557737, 
    -0.584716778985874, -2.05508993669022, -0.435840204017464, 
    -0.690672405603151, -0.644094931133207, 0.819319449167319, 
    -3.29488962094813, -1.77379174603864, 0.00997477576819977, 
    0.273086337101371, 0.0666730238904678, -1.71079059720761, 
    -0.936403752586216, -2.34531616755034, -2.255088724057, 
    -1.73637946614907, 0.400657567587841, 1.08985889692963, 
    -0.581153426547974, -0.960249414179951, -1.61909776581355, 
    -0.38786762448987, -0.0036604532544688, -1.2002009881696, 
    -2.59847018058199, -0.456471533790478, -2.81820090646589, 
    -1.89716551818248, 1.00815873215992, 0.352999923130497, 
    0.210036726253163, -0.531363947221796, -2.2909672517635, 
    -0.201221377452437, -1.41828146871538, -1.24868532207409, 
    -1.20013577758447, 0.663222361533345, -2.57028728770503, 
    -0.295178598791597, -1.23529441131386, -0.493581576688421, 
    0.950687690412935, -2.87947848883768, -3.18029894475052, 
    -0.804987406643984, -1.39943328447394, -1.9690180292748, 
    0.554459615187476, 1.40896942516329, -0.653401688967193, 
    -0.994449606649431, -2.13684209985172, -0.162603415920604, 
    0.593108257590389, -1.86802128952968, -3.18550076614505, 
    -0.561387411381405, -0.614555340934274, -0.572018529897254, 
    0.43780951889237, -1.14546903692243, 0.255297004738648, 
    -3.66420935818551, -2.07472790904336, 0.142241525104263, 
    -1.89082831379771, -1.50443700551746, 1.24857564387656, 
    -0.649314542101295, -1.88905230336708, -0.750176868029419, 
    1.62564841354706, -2.8871116284994, -3.72149680234679, -0.55266508692889, 
    -1.65682615888965, -1.41478875864303, 1.58956985522924, 
    -1.71695255957415, -0.769163461347169, -3.13501665075, 
    -0.637926933721236, 1.35017513433292, -2.02180845833786, 
    -3.37528146016308, 1.20276566381504, -0.184241387072181, 
    -2.07776203283231, 1.22892846960699, -0.883496248608212, 
    1.22068284558463, -3.15739726637691, -2.67252184879103, 
    0.385152689518612, -2.16779803620272, -2.36215126498514, 
    1.75773910108254, -0.951817538315203, -2.58416622541754, 
    -0.471323050789599, 1.63679508184445, -2.40759010597062, 
    -3.32247245395689, 1.24332655159031, -0.154175773382644, 
    -2.47086110251706, 2.48573666132463, 0.494732368389039, 
    -1.71727192134767, -0.977956894243632, 1.21883690088376, 
    -1.77223477781338, -2.25947204152711, 1.99022382673892, 
    -0.578678004303332, -3.04650478703427, 2.43378634698859, 
    0.49475988076535, 0.549027340687213, -2.33745800463993, 
    -2.75239647109822, 1.09956874112329, -0.301575932956257, 
    -1.88191082737041, 2.60530466010373, -0.0934679912443365, 
    -0.163759293312933, 0.938305526220872, 1.20083298015654, 
    -1.45201317223908, -0.836328951922322, 1.98745341284692, 
    -0.376039329233328, -3.18210556324884, 3.83455261552685, 
    -0.662767443150541, -0.550143401484422, -0.569414942986262, 
    0.695896394111791, 0.235727644134314, -0.315101508017163, 
    2.20845311918272, -0.490373558439094, -0.680095158485436, 
    1.46443058681273, 2.2891377814732, -0.257574229727237, -1.39758201886746, 
    0.0373013398320292, 1.57552090030681, -0.255513142073945, 
    -1.51834404564575, 3.3476631760529, -1.27820205947662, 1.50763576175298, 
    1.85284886943441, -0.227533524015618, 0.58125708073991, 
    0.884741181619653, 1.79826743019442, -0.88079728188792, 
    -1.76511268464911, 2.56090464094426, -1.72907266698972, 
    -0.199367987642445, 1.49658997596335, 0.66881360232432, 
    0.408211090475478, 0.724793284022543, 1.39347988255543, 
    -1.45221307648387, 0.868803456120699, -0.292731382573886, 
    -1.76359166713985, -0.393844613680686, 1.0673950267927, 1.41214770135698, 
    -1.02579159095923, -1.41683995588829, 2.38544222170949, 
    -2.04391197697848, 1.70732939500965, -0.739944264114876, 
    0.558376386787012, 1.19009716045323, 0.0212189511806675, 
    -1.58391401612172, -0.978810350109602, 0.493497150070361, 
    -3.13942678246991, -1.50478956310847, 1.26681162992852, 
    0.494164097316788, -0.434428165468179, -0.666993610908852, 
    0.662134506584577, -1.76105348423301, 1.07840734149033, 
    -0.37331683862713, -1.97092826966133, -0.870125382108963, 
    0.561269145902549, 0.0929048397063668, -1.67991507399174, 
    -1.53302723179882, 1.31366392998666, -2.95952228021802, 
    -1.40480124190567, 2.21660788145358, -0.760625460577309, 
    -0.153971572323054, -1.65260717540469, -0.613133161188473, 
    -1.54190879946835, -0.801734197197082, 0.025962870440209, 
    -2.64523544233777, -2.73932935270671, 0.0244779495493085, 
    0.306073684753963, -1.65981025942748, -1.12910335399114, 
    0.924417550317727, -1.58277924664632, -1.63682658170037, 
    -0.788472464784942, -1.41055234511493, -1.23726191719084, 
    -2.06868878054208, -0.234179281892047, -1.56775751714423, 
    -1.71725790482918, 0.907491157734924, -2.08418477502286, 
    -3.51393334294018, 0.698549818428812, 0.0347166073839363, 
    -1.29333288753725, -1.96778295806951, 0.288211824093769, 
    -0.438120408452766, -1.27400998531436, -1.80615811647785, 
    -1.34779279374366, -2.88798374306438, 0.177052738771001, 
    -1.76031760632701, -0.928879292745158, 0.558509343145766, 
    -0.692842764077243, -3.43654804894354, -1.09911036806597, 
    -0.142700527702185, -1.21063124040312, -2.37655033602907, 
    0.0834852708786683, -0.0144463225490256, -0.71170518237537, 
    -1.03426755624074, -0.864410087888937, -3.73131020788826, 
    -0.122809874569367, -1.69891735328859, -1.11724202607488, 
    -0.318519514136813, 0.221555120107621, -2.22911744824676, 
    -3.50225108811066, -0.0912606086567732, -1.30785907994815, 
    -0.133208697247832, 0.0328774364880095, 0.15244113675258, 
    -0.983538257443754, -0.366221737636531, -3.35537520309196, 
    -0.802771505468937, -0.641770237473907, -1.61874922247829, 
    -0.772899842258547, -0.994046153020075, 0.630555236869474, 
    -0.799849075561002, -4.06000122474407, -0.197454632675751, 
    -1.62963444426059, -0.844626249527069, -0.119037264869097, 
    -0.280232238016344, -2.27913976792685, -0.45911152099909, 
    -2.02617449308026, -3.2663547782836, -1.00879831161863, 
    -1.28463974732797, -0.982493115448323, 0.803953716696724, 
    -0.0923521197144658, -3.80976475557336, -0.764124457347805, 
    -1.26073931982987, -1.85017135505824, -0.46939709355491, 
    -0.576092067780094, -3.23052437048626, -0.422529673953997, 
    -0.774779056851271, -4.40958103878749, -0.999348322769603, 
    -1.24079833069049, -1.05208542795737, 0.611151742473706, 
    -0.976271428547868, -4.2209886753261, -1.33827187220091, 
    -0.310838826989308, -2.29575403175575, -1.25638876091122, 
    0.262664538195653, -2.83223601024313, 0.0815211629307193, 
    -0.824730297415988, -4.10610612042259, -0.835471973008012, 
    -1.32274426639594, -1.55468289978024, 0.0967950037933596, 
    -2.52229029526472, -4.36689493117315, -1.12108976936922, 
    0.563062082918762, -1.82319625540722, -1.46300349353349, 
    -1.95277801685504, 0.435282210779296, -2.33151136866143, 
    -4.14397617129742, -0.755852270807461, -0.882291079330925, 
    -1.74632565162032, -1.06172696831473, -1.05710659340471, 
    -3.63393422833901, -0.447816199583408, 0.619161323399845, 
    -0.827473829600196, -1.16820587147802, -1.54123989927974, 
    0.130092105669952, -4.73895204908567, -4.16111795791626, 
    -0.478214722004571, -0.200092011941105, -1.51512894247762, 
    -1.12044733901215, -2.7398251921718, -0.183485888708196, 
    -0.734612294868432, 0.0756112658430022, -1.48565479756675, 
    -1.38456548121185, -0.765156538772585, -3.2744456171915, 
    -3.58409850318321, -0.137284273427858, 0.718260648914269, 
    -0.949986318642091, -0.50349848369448, -2.37350075578534, 
    -0.471779262754501, -3.00473390838594, 0.619822773694442, 
    -1.67255877068658, -1.61283175808833, -0.571571815173279, 
    -2.84002269904879, -0.422724680045568, 0.691019325755137, 
    -0.251533192997648, -1.06236837579148, -2.16221665292154, 
    -1.05999060824075, -1.93965019391714, 0.242985330580277, 
    -1.2297285106527, -2.01320899861121, 0.0552815967616513, 
    -2.4694087539085, -1.00643418511793, -0.272946135707283, 
    0.198870803232864, -1.61655052458545, -2.34495239360569, 
    -0.795298039569408, -0.828063758708958, -0.467926618403714, 
    -2.02247373360032, -0.765110738935971, -2.38943909373079, 
    -1.69330154739948, 0.753865160515552, -0.305381045662987, 
    -1.38690068067415, -3.01305496589518, -0.634339179707914, 
    -1.74540654846969, -0.235147092063801, -2.07066341338562, 
    -1.29740713833216, -1.77598403459927, -1.36437313561761, 
    4.04356809131269, -1.08426546942589, -0.551929416156758, 
    -3.29758419106273, -1.49266458499764, -2.31831863982754, 
    0.150364249786481, -2.6129540063417, -0.862328808776344, 
    -1.8387631419389, -1.18524234655374, -1.46461072964831, 
    -0.177435366264608, -4.00566074805969, -2.29513521863333, 
    -2.02187204756914, 2.57709905615756, -2.20768393892932, 
    0.172856535374781, -2.88622973744221, -1.75469436922222, 
    -1.58979546787126, -0.223863531399489, -4.37126955555025, 
    -2.41077073535027, -1.7466086150253, -1.26438803777872, 
    0.762214796353854, -4.42535703622188, -2.52585823353635, 
    -1.30373547307519, 1.7735469125505, -3.39587669807236, -1.59429291383045, 
    -1.1798886199303, -0.866981450563242, 0.408904458611145, 
    -4.50616755901967, -2.89452937727045, -1.16642543244946, 
    -1.95613101421256, -0.402944265977139, -0.532891934720996, 
    -0.658924956916966, 1.85190092041122, -2.89183081767836, 
    -2.50752418783209, -0.503332346320161, -1.18110588575401, 
    0.68702045749357, -0.21946453638018, -0.817842904101733, 
    -1.61731264345078, -1.55571701980413, 0.527204845810478, 
    -0.83145212437772, 2.96753157524781, 0.383509632422001, 
    -0.55429844751492, -1.48041849327292, 0.150018404492575, 
    0.703338657259517, -0.711502412667067, 0.876442825885933, 
    0.206710752768062, -1.45295455040465, 2.96762948738678, 1.23569777365766, 
    -1.09004161361968, 1.48167267560471, 0.140502613746042, 
    -1.21373001420339, 5.20025866121111, 1.89958891053138, -1.29746019081608, 
    2.98479194124444, 0.766646272267045, -1.61455509671514, 2.46066515023738, 
    -0.611907166994381, 5.78723540153079, 1.20163741486258, 
    -1.88271848389783, 3.95919160098665, 0.364595316894506, 1.94597121675894, 
    -0.446485755776342, 6.60187978198992, 0.646769077620851, 
    4.18025753856767, 1.05559972829607, 0.775599385912471, 1.48286935463306, 
    2.99947753091509, 0.895203854974942, 5.95472633368029, 2.48348275187945 ;

 NLcost_function =
  10457.7055852316, 2263.75352520979, 0, 0, 0, 0, 5640.64048697727, 
    2553.31157304456, 0, 0, 0, 0,
  3237.34685094907, 415.281719759614, 0, 0, 0, 0, 1516.04369292778, 
    1306.02143826167, 0, 0, 0, 0 ;

 TLcost_function = 10457.7055852316, 8435.32259328932, 6488.86257662177, 
    5247.24540629257, 4213.68920600726, 3806.84974599203, 3271.03113653136, 
    2958.4635974877, 2698.75337892342, 2475.99322492623, 2245.93939466651, 
    2074.68625877632, 1908.63503562244, 1750.4717021438, 1640.02696812922, 
    1558.86047205107, 1472.65439659831, 1421.55343616495, 1378.53964850306, 
    1339.85344540683, 1306.79957287655, 1279.40061528664, 1262.70034042738, 
    1248.57264257308, 1236.03976072109, 1224.56258336222, 1217.11550446172, 
    1210.91593965177, 1206.59478632267, 1203.42617175139, 1200.97478176555, 
    1199.00141438448, 1197.76109699686, 1196.79829402133, 1196.08444900022, 
    1195.5066244591, 1195.18284435356, 1194.91112322915, 1194.71645586882, 
    1194.6132582183, 1194.54041805797, 1194.48333263843, 1194.43535788622, 
    1194.40351082301, 1194.38147232162, 1194.36502006591, 1194.35389074546, 
    1194.34785036665, 1194.34353763125, 1194.34028909083, 1194.33812858943, 
    1194.33812858943 ;

 back_function = 0, 3.11396602399619, 15.5455835354681, 35.4982752667702, 
    71.0113504945423, 93.2587214344107, 136.688173376378, 171.808997426075, 
    208.531211431843, 246.86421405536, 295.185591698408, 338.378111755483, 
    387.395964349506, 441.803122279072, 484.699375317241, 519.014402018616, 
    558.472271490882, 583.536805519425, 605.797481556441, 626.833623311485, 
    645.658176581959, 661.966814099471, 672.27177746976, 681.245339606457, 
    689.437608117917, 697.161733539388, 702.306709543374, 706.689444800455, 
    709.807682673028, 712.134396505301, 713.962781531381, 715.456477911228, 
    716.40769497792, 717.154875102982, 717.715328408461, 718.174137615239, 
    718.433667768201, 718.653316658099, 718.812068113387, 718.896853666287, 
    718.957068632815, 719.004550212142, 719.044722379091, 719.071565250732, 
    719.090249820258, 719.104278801689, 719.113820890214, 719.119023001699, 
    719.122751983337, 719.125572387632, 719.127455730403, 719.127455730403 ;

 Jmin = 3.06902585039813, 2.47643039158131, 1.9088505238906, 
    1.55032829979731, 1.25743229831308, 1.14456594788744, 1.00006436094138, 
    0.918641994105291, 0.853201640603157, 0.799077751718736, 
    0.745744676849571, 0.708162691278591, 0.673816874533219, 
    0.643367520006713, 0.62354404796668, 0.6097945338429, 0.596075324457575, 
    0.588434406950661, 0.582343985343948, 0.577164216791876, 
    0.572988334397214, 0.569733654992256, 0.567856821099675, 
    0.566344235415859, 0.565070394376818, 0.563968985150876, 
    0.563293386355125, 0.562760200866389, 0.56240718092317, 
    0.562160108072396, 0.561977274628594, 0.561836505442613, 
    0.561751663088709, 0.561688384189086, 0.561643368278409, 
    0.561608440814185, 0.561589585362219, 0.561574303708656, 
    0.561563763457727, 0.561558360054172, 0.561554654934934, 
    0.561551836493198, 0.56154954666627, 0.561548078084736, 
    0.561547093805394, 0.561546382646396, 0.561545916840991, 
    0.561545670834437, 0.561545499520053, 0.561545373874823, 
    0.561545292537002, 0.561545292537002 ;

 zeta_ref =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, -0.000159060948906429, 0.013673910803881, 0.0160926893912428, 
    0.0132446340833114, 0.010315316828801, 0.00969144308471488, 
    0.00886926280492229, 0.00277516430233557, -0.00489991356365215, 
    -0.00576368931800111, -0.000733858995061766, 0.00431468554332382, 
    0.0068159845225507, 0.00675267959182694, 0.00451825646183626, 
    0.00360522182287072, 0.00746121916907461, 0.011577044491648, 
    0.0100995018309415, 0.011753385409234, 0.014491825933484, 
    0.0178347933084365, 0.0136482481565119, 0.00638400183611861, 
    -0.000375100997789568, -0.00328860891039923, -0.00284233677201645, 
    -0.00430892596370287, -0.00868203338294476, -0.0126329310384841, 
    -0.013122920821751, -0.0087410709532008, -0.00194741011347665, 
    0.00618915331448503, 0.0130044756837716, 0.0140387043974101, 
    0.00852808659786121, -0.000527780096031716, -0.00779749060657101, 
    -0.0144777412757372, -0.0208224811954473, -0.0199651363727974, 
    -0.0137039772303316, -0.00313991931888989, 0.0033115903579544, 
    0.00259704652004861, -0.00373762255592912, -0.00728692582942897, 
    -0.00783883880437669, -0.00573303449434986, -0.0121700115718127, 
    -0.0139313954250775, -0.014353792935076, -0.00639084158887991, 0,
  0, -0.0010462100678213, 0.0247044525910482, 0.0479412260278583, 
    0.0456920436162593, 0.0381299653928739, 0.0287901187970671, 
    0.019367540291966, 0.00686970839004419, -0.00792058554757884, 
    -0.00668907195239949, 0.00324601154360612, 0.00884148808576429, 
    0.0103024777564694, 0.00875342566886284, 0.00538184358749446, 
    0.00398378760694434, 0.00781637828454632, 0.00966210971207084, 
    -0.000278048282625941, 0.0011348863996023, 0.00799617922508818, 
    0.0175627024618318, 0.0140765638208986, -0.00412927525217435, 
    -0.0239354017810475, -0.0387224483446389, -0.0461963967574461, 
    -0.0561073866606127, -0.0693331715244771, -0.0732037462495482, 
    -0.0617481232534194, -0.042880084944956, -0.0173913720904776, 
    0.00932332376782411, 0.030749386639018, 0.0353885590206936, 
    0.0106284495497612, -0.0321452071932125, -0.0664553453072798, 
    -0.0902644070010637, -0.107468459430814, -0.096727313673908, 
    -0.0712600742025809, -0.0405823478965354, -0.0228133791408865, 
    -0.0244646586106245, -0.0336363498578712, -0.0382148036116927, 
    -0.0307279225238522, -0.0248772316345747, -0.0342792572481319, 
    -0.0427018698594024, -0.0437663916120157, 0, 0,
  0, -0.00125906557392963, 0.0200977278497454, 0.0420824445815106, 
    0.0440004778143824, 0.0348117572381584, 0.0176669159185685, 
    0.00255329077804416, 0.00105688379735974, 0.00585708317385793, 
    0.00793100372112389, 0.0113105420726382, 0.0101411764057218, 
    0.0141346245190525, 0.0191956834458047, 0.0193742174751473, 
    0.0156379397573578, 0.0126247457217522, 0.0128487008174886, 
    0.0139241482247521, 0.0215635722265146, 0.0461683370170887, 
    0.0544609545897762, 0.0451090063016134, 0.0200437464437252, 
    -0.0010431098655617, -0.0188043663452061, -0.0343911963036265, 
    -0.0517085619475406, -0.065324682578552, -0.0608831049255055, 
    -0.0344286520166794, -0.00568692432026508, 0.0175666713756436, 
    0.0407031607251418, 0.0616648368078518, 0.0593845998384459, 
    0.0224253806170833, -0.0286836212173579, -0.0648771375852368, 
    -0.0910271654322957, -0.113554518903137, -0.109235308427472, 
    -0.0804356932190945, -0.054513020216619, -0.0424914058066991, 
    -0.0385078130199638, -0.0464200889953039, -0.061408684529419, 
    -0.0598254792691222, -0.055886120787995, -0.0584921820223134, 
    -0.068066804007002, 0, 0, 0,
  0, 0.00233844804027245, 0.0200984715138796, 0.0205838632673946, 
    0.0132548477367016, 0.0128638954915552, 0.00558049748879909, 
    -0.0123640890243118, -0.0128172644098489, -0.00235953053757842, 
    0.00442276236040061, 0.00368537248616632, 0.00154979032421306, 
    0.00869413874611191, 0.019107192862947, 0.0266540905349521, 
    0.0264724676264394, 0.0219313325001814, 0.0190399911714246, 
    0.0219734442808696, 0.0373742860856312, 0.0654441664743482, 
    0.073007697073456, 0.0566237058044607, 0.0338854427892437, 
    0.018290894253241, 0.00178313213185693, -0.0162540818534865, 
    -0.0399674610925515, -0.0518858712449954, -0.0353630046242047, 
    0.00160081708306761, 0.0331033099191999, 0.0472808156661538, 
    0.060588676021747, 0.0732598853471994, 0.062722452406701, 
    0.0266556550858951, -0.0121767095216263, -0.038532401387079, 
    -0.0591655464335469, -0.079232530056261, -0.088683295634555, 
    -0.0759721318839706, -0.0571312586747078, -0.0419235082604875, 
    -0.0390823929260848, -0.0508423573143728, -0.0772876168325593, 
    -0.0776703633236329, -0.0758802317506565, -0.0731314407031505, 
    -0.0814229958729939, 0, 0, 0,
  0, 0.00074991052012677, 0.0150060353185743, 0.00612335822260639, 
    0.00799303489328136, 0.0196349109193641, 0.0202690746123212, 
    -0.00169193270638371, -0.0145899001864508, -0.0140889146736742, 
    -0.0122793769319827, -0.0108656806794574, -0.0048602652665801, 
    0.0118144015168318, 0.0222003553836527, 0.0334438342831538, 
    0.0332160860290534, 0.023567991641242, 0.0174817497399133, 
    0.0244949501622308, 0.0346275965279152, 0.0585001171098434, 
    0.0700755126509727, 0.0631761655813548, 0.04899596973659, 
    0.0385667807405394, 0.0274837822436971, 0.0111470000599527, 
    -0.0160755595951645, -0.0316086159906321, -0.0175630840122148, 
    0.0221947155175029, 0.0486893627622298, 0.0488405597912713, 
    0.0420025260066715, 0.0476287729533445, 0.0542809573150426, 
    0.0403228732845537, 0.0212224857860827, 0.00353701600808142, 
    -0.0107321048852068, -0.0267386972500712, -0.0478415743318644, 
    -0.0544833170012883, -0.0453671959376033, -0.0360322404380895, 
    -0.0312386824574107, -0.061045076658108, -0.0815657930411274, 
    -0.0937470233609828, -0.0883639196488446, -0.0831146148714816, 
    -0.0811308559851325, 0, 0, 0,
  0, -0.000458429674936386, 0.0105626838584882, 0.00880366400772009, 
    0.0101660848704182, 0.0229722618500492, 0.0286912457584614, 
    0.00856423808744866, -0.00398427564290723, -0.0119925720749795, 
    -0.0106357729175717, -0.00388905815812981, 0.0107612171506671, 
    0.0223783066340654, 0.0379365596575637, 0.0478700140019147, 
    0.03863324580068, 0.0210427343709493, 0.0122169562440981, 
    0.0133792300185275, 0.0209898750106084, 0.0360606715276162, 
    0.0490420146104165, 0.0559061672552854, 0.0537366026708151, 
    0.0508384865477101, 0.0469784884582058, 0.0383769090326841, 
    0.0148784282566769, -0.000732143603712517, 0.00217437180171671, 
    0.0281305105531537, 0.0403431140326417, 0.0180539771334802, 
    -0.00695704675810761, -0.0128497235014633, 0.000825627325898899, 
    0.0165536526897446, 0.0317335828010668, 0.0364369336222939, 
    0.0326262398505043, 0.0186977527323777, -0.0112010057245331, 
    -0.0344793160875913, -0.0367498787160755, -0.0298822629868306, 
    -0.0459052334003382, -0.0616335739773131, -0.0886092864240825, 
    -0.0993531876728611, -0.0946976648572862, -0.0891975433685508, 0, 0, 0, 0,
  0, -0.000289214787087966, 0.0107502310641713, 0.0154476820959108, 
    0.0176045724994278, 0.0304564787776926, 0.0199896386174668, 
    0.00340928001714354, -0.00373990218769735, 0.00215929653517255, 
    0.00350184513896237, 0.00574307108842477, 0.0148358350991029, 
    0.0303028283394906, 0.0484542058951063, 0.0692374054495794, 
    0.0633398098195467, 0.0358759850586135, 0.0140708605100052, 
    0.00501067724412472, 0.0094492144186433, 0.0252065972193193, 
    0.0411961731025526, 0.0472575783979944, 0.0517405711393588, 
    0.0501637199973162, 0.0537610491896326, 0.0541762966780802, 
    0.0418631423044849, 0.031010963601894, 0.0295973914055222, 
    0.0330194871546699, 0.0123733447120565, -0.0423808537456994, 
    -0.0842741107004708, -0.0968686277037605, -0.090523644278607, 
    -0.0707498321270664, -0.0367712139825201, -0.00226535208359737, 
    0.012463002626322, 0.0101255248430706, -0.00166032222056984, 
    -0.0219664179405637, -0.0429818436662452, -0.0524612681321419, 
    -0.0636053422109744, -0.077126303920689, -0.0938679396715358, 
    -0.0988906946714461, -0.0967362800150732, 0, 0, 0, 0, 0,
  0, -0.00533168246315232, -0.00117663378069783, 0.0243431087260654, 
    0.0294460970183758, 0.028404617755387, 0.00738679908855122, 
    -0.0086638202883521, -0.00899863259006788, -0.0053359828789333, 
    -0.00321541133320082, 0.000208007013115243, 0.0104077683508742, 
    0.0255696650312561, 0.0477683832380097, 0.0677967721998566, 
    0.0732094621111304, 0.0471163548388029, 0.0217820736511935, 
    0.00538545487916703, 0.0132664535032446, 0.0239430069884686, 
    0.030963235695813, 0.0356928429474194, 0.0352700781188403, 
    0.0337125989299045, 0.0351401429427095, 0.0405520891375653, 
    0.0457712234466653, 0.0455587952627113, 0.0472094179430691, 
    0.0328106670117503, -0.0287905424300113, -0.114841855220907, 
    -0.166286041926022, -0.178036620002187, -0.177303502232858, 
    -0.165275820054648, -0.130050933867285, -0.0836694079990751, 
    -0.0553881412892827, -0.0414304170825978, -0.036433867217451, 
    -0.0535262052483695, -0.0702065630344053, -0.0781744647524939, 
    -0.0813997288775866, -0.0926827369701371, -0.0970820095656227, 
    -0.0982643092635963, -0.0994675098000206, 0, 0, 0, 0, 0,
  0, -0.00531592812940382, -0.0137537337449695, 0.0273033171772903, 
    0.029937898254686, 0.0171578258636285, -0.000571154942001913, 
    -0.00824885598802378, -0.00231925971314857, 0.00877696432080612, 
    0.0149292011864483, 0.0167658093129844, 0.0223955111977638, 
    0.0345613913196971, 0.048883359283348, 0.0595406566093635, 
    0.0602881468361405, 0.0387353023312329, 0.0163213050640694, 
    0.00182085997164947, 0.00128817461727189, -0.00144459732640698, 
    -0.00485789339177677, -0.014084924620652, -0.0217390170748778, 
    -0.029175973468105, -0.0254855155507933, -0.00987400411599026, 
    0.0116441120462029, 0.0310198453828014, 0.0382987303481248, 
    0.0130948809314201, -0.0750575979835224, -0.177258472939132, 
    -0.222561005619771, -0.225761807991906, -0.226589395611178, 
    -0.218218046246146, -0.181204356364851, -0.131151403075231, 
    -0.100055343550168, -0.0826281691273168, -0.0849449061002546, 
    -0.0988804343967696, -0.0950686168070111, -0.0940125513815963, 
    -0.0917610451474081, -0.0937599146742855, -0.0941822551599345, 
    -0.0939313534215339, -0.100616004284997, 0, 0, 0, 0, 0,
  0, -0.0029020788198307, -0.0179068139457025, 0.00353437886706895, 
    -6.96375249293992e-05, 0.00442493937814688, 4.10228905618643e-05, 
    -0.00196258720780011, 0.0107017832677942, 0.035223827020311, 
    0.0488878931733085, 0.0501313997224494, 0.0503625795592362, 
    0.0549368663821534, 0.0605962554981881, 0.0600439967841528, 
    0.0498061999696036, 0.0305181826136029, 0.0143191104388104, 
    0.00278308839923953, -0.00836284153289136, -0.023837481012098, 
    -0.0450823573688242, -0.0664302481361389, -0.0855957698021339, 
    -0.0948369615643676, -0.0806981879707517, -0.0556995063261495, 
    -0.0304371327617801, -0.00558365287975514, 0.00965906759329462, 
    -0.020402654816227, -0.107799734165407, -0.196367146211933, 
    -0.230443792707054, -0.239049114516059, -0.249853617560477, 
    -0.24279242335985, -0.19875155492594, -0.151044712521748, 
    -0.121397577679583, -0.116372766285926, -0.109738840357963, 
    -0.111594946132511, -0.109881675292739, -0.0957062861789277, 
    -0.0863581367485855, -0.0870420814823505, -0.0915675051325271, 
    -0.0933651854839396, 0, 0, 0, 0, 0, 0,
  0, -0.00368724861420403, -0.0361473912643087, -0.0344624134383807, 
    -0.0222915568568134, -0.000981016807109487, 0.00355584569965819, 
    0.00615197055150224, 0.0172193461810295, 0.0383968354105398, 
    0.0617452395250991, 0.0695340677283779, 0.0667644680179683, 
    0.0699779543808928, 0.0713947716727939, 0.0664585839754234, 
    0.0502750446672613, 0.0327797139308251, 0.0203887427525495, 
    0.00688097272803583, -0.0140154501442007, -0.0425261012239712, 
    -0.0749700356594932, -0.103328718887373, -0.125971294123772, 
    -0.128372797579999, -0.101726445325002, -0.0734424158634028, 
    -0.0546919734482949, -0.0358145899857882, -0.0260837282866502, 
    -0.0548468105082758, -0.114422726293588, -0.170161744588594, 
    -0.198289833677829, -0.221436091973328, -0.238452683729903, 
    -0.234841959762177, -0.197356093149307, -0.160510044626077, 
    -0.139252185982664, -0.133459909110386, -0.127664353394422, 
    -0.122098502115012, -0.115538502286683, -0.100808534038733, 
    -0.0916559906142875, -0.0928055336024805, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.00299654082407326, -0.0474719326342507, -0.0640125467145864, 
    -0.0489766693863208, -0.0176131229568289, -0.00167153604023011, 
    0.00712910800990538, 0.0215035752056343, 0.0400973565350545, 
    0.0561876629722237, 0.0693201914359979, 0.0792839170024278, 
    0.0790586676958007, 0.073536882941254, 0.0673449390682587, 
    0.0565772035578726, 0.0434593388607818, 0.0265749062818859, 
    0.00626200745420793, -0.0235684282030984, -0.0644691172934502, 
    -0.101706141620184, -0.126483610911859, -0.143390929986825, 
    -0.138126955435682, -0.104954731801192, -0.0786085879348311, 
    -0.0665368272597023, -0.0672598376610818, -0.0766359647862954, 
    -0.0975351319114164, -0.128210667614208, -0.148848719109961, 
    -0.162504986263132, -0.185922502115702, -0.204651710514828, 
    -0.209300464254602, -0.193675108253733, -0.1654968283816, 
    -0.15684820201894, -0.153716504431191, -0.145255488217127, 
    -0.134383489799792, -0.120482191235762, -0.109846659802057, 
    -0.103462270037933, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.0094056722981523, -0.0249152107976491, -0.0440406535785211, 
    -0.0497497658186273, -0.0358487090304848, -0.0185529751871304, 
    -0.00122972203110452, 0.0143315123671017, 0.028399332965215, 
    0.0423872067026037, 0.0582356711655851, 0.0744453790165982, 
    0.0766802954955735, 0.0789249630693817, 0.0784756979167577, 
    0.0718474784263129, 0.0545575554677124, 0.0327246692304118, 
    0.00816241786552748, -0.0263879826736914, -0.0764654593180895, 
    -0.118586984166214, -0.14096495538178, -0.152665235031676, 
    -0.138806032447094, -0.11055006399736, -0.0975711249357752, 
    -0.100240077993249, -0.119313856043932, -0.143997737258238, 
    -0.16253619183674, -0.174683698012134, -0.170607892278752, 
    -0.160579646809704, -0.168937680425725, -0.187415035718217, 
    -0.203031223333834, -0.196991389105296, -0.181845667922361, 
    -0.171935642966382, -0.161990330655707, -0.152556168769358, 
    -0.145039449261315, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.00740195225198748, -0.00954251220885304, -0.00772416960782518, 
    -0.0172037547130994, -0.0206323476904488, -0.00487853605895627, 
    0.0107988888048355, 0.018494099048518, 0.0200271106751368, 
    0.024866066830272, 0.0358861925178585, 0.0481410671475527, 
    0.0552100900956458, 0.0604291767574267, 0.0652914912087822, 
    0.06523030327877, 0.055105593865553, 0.0367011492847978, 
    0.0174581684175203, -0.0103846629249175, -0.0585414596449915, 
    -0.104745784840176, -0.127831436330993, -0.1352794490063, 
    -0.11988744594485, -0.100647856140131, -0.106491845348429, 
    -0.129674087857226, -0.157917026449634, -0.184843991331001, 
    -0.20307360506177, -0.200795558988082, -0.183065704501192, 
    -0.174717805954925, -0.172180410930852, -0.187745790561051, 
    -0.208297623735156, -0.201349947468765, -0.198335373738538, 
    -0.188981589928297, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.0040503931312687, -0.0127110225248399, 0.00665456210411853, 
    0.0067940149124947, 0.00971548317931155, 0.0177800037800493, 
    0.018594915659763, 0.00835054196204241, -0.00228765006001871, 
    -0.00324070418894368, 0.00480618569836305, 0.0174613952027476, 
    0.0280398021436389, 0.0348052890672815, 0.0384947887971392, 
    0.0412691840583128, 0.0391340091266831, 0.0298210000697322, 
    0.020198158564546, 0.00945189185052389, -0.0246466650493764, 
    -0.0722146875040189, -0.0998043069472485, -0.103548794072211, 
    -0.0878852647667885, -0.0766536276543487, -0.0943873202915581, 
    -0.1233553387244, -0.153262319789385, -0.183554312127462, 
    -0.204749100614426, -0.200170499618013, -0.18506747083796, 
    -0.176576814748988, -0.175559125014764, -0.1928403428173, 
    -0.19915832600316, -0.211690889464938, -0.198975676850678, 
    -0.187362420016329, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.0011416367159785, -0.00918383634142598, 0.0186400255769524, 
    0.021797190375169, 0.0161883289754911, 0.0040336833429127, 
    -0.0116747423021934, -0.0291439816084774, -0.042340928900057, 
    -0.0448145375528884, -0.0375088208489951, -0.0218361839559113, 
    -0.00232651604649169, 0.0132907238018414, 0.0220212531846099, 
    0.0281071556326908, 0.0307000871681461, 0.0204300355585407, 
    0.00840534865999853, 0.00714687344596954, -0.0190842792353123, 
    -0.0690759954278698, -0.100184301160887, -0.101087685889756, 
    -0.0820206189627853, -0.069217641857936, -0.0871261281317695, 
    -0.114986915160676, -0.136056824216488, -0.165336368599696, 
    -0.19558781219541, -0.197023374153916, -0.191667972774357, 
    -0.186547363252189, -0.182188533265266, -0.183216990428448, 
    -0.201983437354674, -0.205947969568984, -0.198839869260358, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -0.00401231539939224, -0.0210298833688071, 0.0160361158905199, 
    0.017708768407371, -0.00703649019513484, -0.0303473320116357, 
    -0.0377145711407019, -0.0452295459379222, -0.0564829191874115, 
    -0.0563642889106743, -0.0397613674194183, -0.021376501325466, 
    -0.00668061352743205, 0.00358441595744751, 0.0107493706989707, 
    0.0199888589575959, 0.0233232819296682, -0.00647606081173791, 
    -0.0346565554321134, -0.0359101302564665, -0.0632433841997543, 
    -0.120140215917913, -0.152267628463644, -0.141899261354416, 
    -0.113486754005442, -0.0998389364352911, -0.118923074479801, 
    -0.14369917766208, -0.15297206985489, -0.160922932319724, 
    -0.180279855543199, -0.188055430034499, -0.19121255611176, 
    -0.189828508040601, -0.185296211655829, -0.182910620647857, 
    -0.195893598102551, -0.20323992042682, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, -0.00720939664899104, -0.0432064456402054, -0.0109303891746655, 
    -0.00442313286025693, -0.0280172993464745, -0.0418285032820404, 
    -0.0282256799319323, -0.0266515922055501, -0.0376624817598675, 
    -0.0369268230832208, -0.0210346242370344, -0.0102204285518941, 
    -0.0133481567198552, -0.0109734982752189, -0.00507986711548656, 
    -0.000795647099565924, -0.022444813867561, -0.0756469122486532, 
    -0.116526285745093, -0.126187979927146, -0.148015759662316, 
    -0.197193619282901, -0.222964205689863, -0.202629686436093, 
    -0.166356069820669, -0.152070130106787, -0.169680102139119, 
    -0.186509649984243, -0.184988872202437, -0.171417112506127, 
    -0.16944899962788, -0.16814348226675, -0.17225347318289, 
    -0.179941425987035, -0.192560356517141, -0.18764074875688, 
    -0.190318606470463, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -0.00781652802577529, -0.0562905036367304, -0.034119080633897, 
    -0.0185683171165487, -0.02972909869989, -0.0304671087488068, 
    -0.00946214811679989, 0.000311506247456324, -0.00337014497848966, 
    -0.0124143278363539, -0.0165145255653897, -0.0274729644662768, 
    -0.0351709386170949, -0.0267283820945335, -0.0259172004796519, 
    -0.0498011995606512, -0.106032731855423, -0.166968212257662, 
    -0.206082988391386, -0.218254921553038, -0.217788400396666, 
    -0.234892563862213, -0.246135285294387, -0.229187055443657, 
    -0.202014664593733, -0.192181883614458, -0.208965606089104, 
    -0.216247341788455, -0.206950147719663, -0.18745131413366, 
    -0.17585233875828, -0.167988531083607, -0.171158125466747, 
    -0.182239063823218, -0.201421800701049, -0.202855701919087, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -0.0062202877899089, -0.0460831323343643, -0.0281196842225539, 
    -0.00920162811036545, -0.0189825431127402, -0.0255895151711745, 
    -0.0198469567257025, -0.00415824642546648, 0.000462599859355859, 
    -0.0174841139756156, -0.0394320832933725, -0.0492796633452929, 
    -0.045391530598268, -0.0419335097194373, -0.0565291154404851, 
    -0.105850643722493, -0.174496366068467, -0.218259930688404, 
    -0.225260322616882, -0.218676319817776, -0.206317356550768, 
    -0.201942625214246, -0.208474548579532, -0.220728614210652, 
    -0.225878601224715, -0.221606038542574, -0.230510650462587, 
    -0.229463649055071, -0.210772096876572, -0.188663256343501, 
    -0.179862479669866, -0.171988663097369, -0.155201343369957, 
    -0.161621142550302, -0.194053040767564, -0.190183340173258, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -0.000364820876989899, -0.0209695742235442, -0.00843577968124123, 
    0.00374860272657576, -0.0124775489077276, -0.0391215066088227, 
    -0.0603276656536602, -0.0525846463519827, -0.0539374309005495, 
    -0.0819327829839914, -0.108510874390695, -0.110588387231984, 
    -0.0906391679951433, -0.0730810867208825, -0.0767738637550327, 
    -0.113054646105158, -0.158131095573559, -0.171942794005322, 
    -0.143079266900671, -0.115221873720376, -0.113814856746813, 
    -0.126394212753114, -0.150858983212337, -0.194348575596165, 
    -0.232631418910371, -0.235507206261597, -0.233579425899605, 
    -0.2254120225593, -0.21090614869267, -0.196294167599232, 
    -0.181334113214002, -0.164331217052085, -0.14387358157916, 
    -0.155273722617381, -0.174437511533192, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.00477364205636986, 0.00217299685333094, 0.0125062976746569, 
    0.0124205265977305, -0.0108955848092438, -0.0496183160863359, 
    -0.0891725934485183, -0.105544262322688, -0.130991993211436, 
    -0.177246541548177, -0.20066402505077, -0.184957462394395, 
    -0.149262566303607, -0.108073346330358, -0.0781825319657365, 
    -0.0738870521876532, -0.0830477302730806, -0.0825518046560952, 
    -0.0520673650441905, -0.0245990294276662, -0.0299543086925268, 
    -0.0521522502206632, -0.0907379047085776, -0.154962403117024, 
    -0.212438466080148, -0.226366546043785, -0.219399610647402, 
    -0.212335628018482, -0.204169647585472, -0.197376943390295, 
    -0.173665105441384, -0.159562633504424, -0.152830051773923, 
    -0.162462459468163, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0.0110490023174978, 0.0160636139117801, 0.021773334546471, 
    0.0160877288403801, -0.00565351320945193, -0.0356595737792716, 
    -0.0739965776192137, -0.110524698488812, -0.159158300313697, 
    -0.206758810230943, -0.210132980499195, -0.17691582762027, 
    -0.135727581445766, -0.091261894424708, -0.0516111003843263, 
    -0.0274499812616141, -0.0176738091198976, -0.0136070511229875, 
    0.00568982507554355, 0.0213605831558666, 0.00726116999035322, 
    -0.0208222948356319, -0.0554134757291627, -0.10392801981791, 
    -0.146287582753965, -0.17534350559358, -0.194645604229769, 
    -0.197050538255658, -0.191607596874035, -0.196791761599044, 
    -0.176923575021131, -0.175472935878097, -0.169676672074857, 
    -0.169844059986325, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0.0161433445380042, 0.0164248232590632, 0.0149141604139882, 
    0.0109018613686524, -0.00060999957155575, -0.0162593528550061, 
    -0.0419204085783166, -0.0830424615291374, -0.14519267935707, 
    -0.204473439748649, -0.215340907250042, -0.166557011424131, 
    -0.110935748914797, -0.064804255668223, -0.0311612434506563, 
    -0.0133042064494206, -0.00618703348906341, 0.00270463103291649, 
    0.0191573973270363, 0.0270240660825959, 0.0113890053316127, 
    -0.0186382767646551, -0.0507915298193476, -0.0814133218480911, 
    -0.104945477755102, -0.130738169296939, -0.159464961890119, 
    -0.174279080426119, -0.180963573367597, -0.194987805480911, 
    -0.191759929640001, -0.18331123062197, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.00806157088963978, -0.00268644706698442, 0.00565362729239925, 
    0.00209431794082155, -0.000885448883646368, -0.00557666577383069, 
    -0.0153820018622676, -0.0406427365481443, -0.0976752018853343, 
    -0.179426099775161, -0.221221858983818, -0.184804271372111, 
    -0.12047748542116, -0.0713024917085979, -0.0412780854142894, 
    -0.033138100748691, -0.0330170041653554, -0.0218163721871416, 
    -0.00184750643436106, 0.00734280812268698, -0.00594681114277229, 
    -0.0355257123347959, -0.0685749068707577, -0.0923430456096856, 
    -0.109713046404488, -0.134553448790079, -0.151888599736661, 
    -0.162186683682724, -0.167711755355018, -0.184230294011774, 
    -0.188855826226722, -0.1828754655075, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.000159555946762603, -0.0338398559703723, -0.0206762684759601, 
    -0.00685298901956099, -0.000681824688129207, -0.00266548130461802, 
    0.0065814817209843, 0.00758229924816185, -0.0226521022684009, 
    -0.0956155733797534, -0.165236128464468, -0.164252516601463, 
    -0.111830105390508, -0.0691621928567464, -0.0481997093320319, 
    -0.0424765785041713, -0.0407175165938616, -0.0360395204864626, 
    -0.0309869212230974, -0.0379260193715879, -0.0577459721878975, 
    -0.0830491214609445, -0.106505920897097, -0.116850384779354, 
    -0.123550683829839, -0.142142506620489, -0.153540184522261, 
    -0.152746599371163, -0.16245695614285, -0.177953556898988, 
    -0.184038484156127, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, -0.000875863980285943, -0.0356064015084589, -0.0192153889498858, 
    -0.00407238262703955, -0.00566344530328925, -0.00742359879223595, 
    0.00311088507558404, 0.0133318309475527, 0.018420421663339, 
    -0.0128596738660651, -0.0737965047736408, -0.0915261091931554, 
    -0.0580499713559402, -0.0286793901785967, -0.0206011689741616, 
    -0.0218554259619612, -0.0350757296120166, -0.0619265160163588, 
    -0.102187995380513, -0.14377826956508, -0.171000129369289, 
    -0.180514901182447, -0.177772574298765, -0.165086801736673, 
    -0.15480160250188, -0.170563931614465, -0.186400910594846, 
    -0.178778363075475, -0.185919933427965, -0.188037687967851, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -0.00141782306180556, -0.0239050841591091, -0.011753819417765, 
    -0.0073284507037806, -0.000859521567093844, 0.00263233222267986, 
    0.0101644760297507, 0.0123335985242928, 0.0203164918541965, 
    0.026904932847345, 0.0155691401891689, -0.00643878459964545, 
    -0.00694797984667206, -0.00588372996241086, -0.0116888799030686, 
    -0.0320012356340374, -0.0825505392861135, -0.149978873984617, 
    -0.226892249188172, -0.286355811855329, -0.298237457508822, 
    -0.273279463458499, -0.239893355698391, -0.207666429022979, 
    -0.190722463969829, -0.194899162403114, -0.221288529976326, 
    -0.2325935451045, -0.219886050103537, -0.206978203985328, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -0.00419908773185676, -0.0256164058651286, -0.014251152426268, 
    -0.00806736641099442, 0.000589713330769563, 0.0195355057152185, 
    0.0353619110046491, 0.0385573909019647, 0.0369483416708943, 
    0.0453403069525955, 0.0580425873105101, 0.0356901329062996, 
    0.00456534900844467, -0.0249961860419821, -0.0558112971294267, 
    -0.103155743484387, -0.172868521569328, -0.223755639774186, 
    -0.272587741790085, -0.311309463545095, -0.308087811667022, 
    -0.275750582506315, -0.239694707063925, -0.206343542818799, 
    -0.195044594415813, -0.21095257540145, -0.236218707682508, 
    -0.242139014589928, -0.223645239605403, -0.206095251403718, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -0.00241277847523811, -0.0233678620667373, -0.00961102802363489, 
    0.0127922736569092, 0.030937688619943, 0.0367720309475558, 
    0.0404812953283352, 0.0460890108884413, 0.0494801145154791, 
    0.0567870665795796, 0.0532202846059679, 0.0286361701791327, 
    -0.00782797229693523, -0.0502748628989004, -0.0950558257125829, 
    -0.146640601294469, -0.187077725552953, -0.190334154002339, 
    -0.203134555382775, -0.236444554876082, -0.241789745975685, 
    -0.22358616792504, -0.204639428038272, -0.192979598076744, 
    -0.200724647985755, -0.203646818459106, -0.233155752206234, 
    -0.228818435342463, -0.205809674779921, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -0.0010470655225473, -0.0109886241089416, 0.0152663318780403, 
    0.0419502542839353, 0.0515828465593307, 0.0406011176634265, 
    0.0339199414104578, 0.0357846293534481, 0.0447217286213254, 
    0.0544562008163242, 0.0491235892179033, 0.028992622977146, 
    -0.00561178150533431, -0.0523907322505486, -0.0960681625282149, 
    -0.129655955787821, -0.140729098303303, -0.137476041626791, 
    -0.139020343851262, -0.162762459428273, -0.177589667503001, 
    -0.182504862442046, -0.183514258596526, -0.185291561014427, 
    -0.209359514348179, -0.214046310085821, -0.224120026000302, 
    -0.218587056884372, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -0.00433143280163714, -0.0165433867366032, 0.0154203489174487, 
    0.0436289235397168, 0.0411454513546906, 0.0412322157080308, 
    0.0372855690696953, 0.0372801846611827, 0.0361148170339874, 
    0.049614079599452, 0.0503679128596674, 0.0399209253684991, 
    0.00279221064040629, -0.0442240142367597, -0.0752077913148766, 
    -0.0982859037968211, -0.118850877027342, -0.130507832722863, 
    -0.114511091964049, -0.104310424851884, -0.116464115916725, 
    -0.145902733273091, -0.166796653251538, -0.169976234161031, 
    -0.189449551773323, -0.201145899556563, -0.210433515877876, 
    -0.210303151751051, -0.204713480298208, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -0.0036328379095124, -0.0244449040917213, -0.00540937156859158, 
    0.0140245592638988, 0.0173512580867386, 0.0276057517929257, 
    0.0254070226065413, 0.0183515858413136, 0.0152066450539076, 
    0.0247563725592626, 0.0285642042377055, 0.0202680349953332, 
    -0.0195193300526538, -0.0682355563630555, -0.093451523357101, 
    -0.106921304735141, -0.124093995006101, -0.133724488695619, 
    -0.1183859248887, -0.0907634583140728, -0.0938976340089321, 
    -0.129644128475676, -0.15924776925165, -0.168580733121128, 
    -0.173445513153709, -0.190968829214765, -0.204203025209615, 
    -0.210132845014231, -0.207010942102688, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -0.000171544772935114, -0.0184498673915661, -0.0144800254560342, 
    -0.00578679109731116, 0.00467380921313643, 0.0119988616245785, 
    0.0040033877651056, -0.00460880448972547, -0.00626281392849921, 
    3.14481356770787e-05, -0.000942484798145868, -0.0153261556653697, 
    -0.051604675067961, -0.0871041097839941, -0.103023282046566, 
    -0.118925354307036, -0.139958172705974, -0.15119127857262, 
    -0.14690331339028, -0.119490161397964, -0.104708199668348, 
    -0.12665705636, -0.157923936162623, -0.175796759942387, 
    -0.178685147098101, -0.197718231827906, -0.202190474076474, 
    -0.204845228378153, -0.202581591301036, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.00482778288314441, -0.00148705690281193, -0.014737101366506, 
    -0.0113440298316287, 0.00388816688857755, 0.0106759970332805, 
    0.00588266622754233, -0.00160531953858339, -0.004708423120337, 
    -0.0097202769756186, -0.0220228049953448, -0.0390395160331178, 
    -0.0595847805650665, -0.07697532545736, -0.0854447914632009, 
    -0.11176265278784, -0.151512563210167, -0.173710706336435, 
    -0.178942632692948, -0.158248527645759, -0.134973622361429, 
    -0.143359545164643, -0.16318027680422, -0.179245655800344, 
    -0.17494700423038, -0.186066189722192, -0.189747312581487, 
    -0.191080595952866, -0.193161637137007, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.00629173593875241, 0.0146832037629832, -0.000789290186891054, 
    9.38061505239538e-05, 0.0179361672788966, 0.023300722726872, 
    0.0145683334417158, 0.00566931855298235, -0.00601201397552951, 
    -0.0216347832173339, -0.0423609800379173, -0.0601600859856177, 
    -0.0684592622790695, -0.0725125336902871, -0.0814259210889661, 
    -0.114500526420401, -0.156921423945744, -0.180778422095679, 
    -0.189367018979016, -0.182687047349666, -0.166260857655733, 
    -0.167289188773827, -0.167655671879229, -0.18068743319854, 
    -0.178640284922552, -0.179960666221554, -0.172979911749244, 
    -0.167550999901286, -0.17961166343471, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.00478242423908447, 0.0254706838600644, 0.0264408495028405, 
    0.0311393074037147, 0.0428485520114882, 0.036268432376557, 
    0.0195580336594009, 0.00115468363441185, -0.0169164423705161, 
    -0.0412544235489262, -0.0738120120279181, -0.0896376252557972, 
    -0.0914873605407519, -0.0850986744968654, -0.084937056149135, 
    -0.108689494672492, -0.137412149236035, -0.151775936892123, 
    -0.166550093042148, -0.184328047535008, -0.185990781857041, 
    -0.18135420722535, -0.173740336396727, -0.1699122503477, 
    -0.161391113196915, -0.151589154079601, -0.135789006167606, 
    -0.134472099416099, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.00141896521310437, 0.0217705235732107, 0.048195299513729, 
    0.0588203710945841, 0.0496869658567413, 0.0373566238972158, 
    0.0101954716741399, -0.00533320943994543, -0.0247682738702065, 
    -0.0564218730563905, -0.097943574351063, -0.115203335976391, 
    -0.107898672945007, -0.0969993686201018, -0.0851870810938133, 
    -0.0878171044371905, -0.09688997995647, -0.0990317584642712, 
    -0.114607518477426, -0.147361885563287, -0.165179558595272, 
    -0.164907104460689, -0.163833003880363, -0.147406148297585, 
    -0.132465148921826, -0.123967305466574, -0.124225079015236, 
    -0.12602476379649, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -0.00135825550753611, 0.0153758036040194, 0.0539171578053287, 
    0.0625916639833684, 0.0448537948612845, 0.0173502396431109, 
    -0.00345183278561497, -0.0160029819865104, -0.0267533468503743, 
    -0.0566454164061042, -0.0986499094249244, -0.11098646142308, 
    -0.103465060431259, -0.0914198192050717, -0.0743831405081152, 
    -0.0652954452543518, -0.058053959820162, -0.0501502536157771, 
    -0.0528631689697858, -0.0788527525490811, -0.103708325144139, 
    -0.115732900101007, -0.128510084655789, -0.123560973270487, 
    -0.117137407224507, -0.119582814626209, -0.132332007917903, 
    -0.126854630571831, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.000289937861280725, 0.011574090486473, 0.0457943446802845, 
    0.0523860076244735, 0.0307055375994427, 0.00811088816150917, 
    -0.00632316951247261, -0.0127699018888779, -0.0183180386134198, 
    -0.0409661011743968, -0.0794311141142717, -0.0961758140221216, 
    -0.0838811586681314, -0.0679570729396226, -0.0576023847999752, 
    -0.0527040226085409, -0.0482370135528056, -0.0431490325264242, 
    -0.0424953240310826, -0.0552703146308834, -0.0685821386744628, 
    -0.0880981538875066, -0.109143254041331, -0.120159971517277, 
    -0.115348901361154, -0.118422758650426, -0.13358971837355, 
    -0.11998978935804, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.00324505679602453, 0.0161208901197458, 0.033171663027401, 
    0.027285397788472, 0.0109677050729379, 0.00485257205732607, 
    0.00933304845573103, 0.0100350878917399, 0.00653523461162065, 
    -0.0112841457029932, -0.0485827662779787, -0.0689083544589886, 
    -0.055771920846552, -0.0390716892421104, -0.0396471652094866, 
    -0.0509895971076445, -0.0618068181418859, -0.0659503378118485, 
    -0.066615616461312, -0.0610639235536099, -0.0632841364528643, 
    -0.086042200029382, -0.108155975108101, -0.125969924293441, 
    -0.123801792954275, -0.124043906091211, -0.127456866530051, 
    -0.120377968812702, -0.100264482374892, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.00340606505407028, 0.0113914588395497, 0.0112266378998395, 
    -0.000791997611224926, -0.000511713133044002, 0.022154801304699, 
    0.0362762407445131, 0.0348879737448508, 0.0331655443834845, 
    0.0192627876247282, -0.00736020336556459, -0.0238969651095303, 
    -0.0130298654216751, 0.00104100116710082, -0.0106026934435675, 
    -0.0423484517387582, -0.0701250338785498, -0.0794787649756037, 
    -0.0750644637423839, -0.0693206991183858, -0.0751087567664643, 
    -0.0854331460809947, -0.0992046613587567, -0.116733947416669, 
    -0.125295731922294, -0.126126561331422, -0.124473701444894, 
    -0.126996152106909, -0.110034716532118, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.00247737597535276, 0.000905533762739144, 0.000300709800665529, 
    -0.0081013660926052, -0.00246622065748815, 0.0254218836007998, 
    0.0397524804255429, 0.0454454486348856, 0.0480639490216295, 
    0.0407512653643602, 0.0301210225350058, 0.022511408621176, 
    0.0265147469178052, 0.0282973145787341, 0.00512817103254975, 
    -0.0333356755018063, -0.0655725269419792, -0.082600763311025, 
    -0.0842656674265641, -0.0805973085056745, -0.0744644729207358, 
    -0.0776734611044773, -0.0925364748994739, -0.112780806486203, 
    -0.117762459594303, -0.117987207346515, -0.121672008478914, 
    -0.125390258570053, -0.106699787917406, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.00161369864968152, 0.00354751862046818, 0.00742498141979972, 
    0.00579661624039504, 0.00843585799733833, 0.0159945752814398, 
    0.0262581870743348, 0.0417507340230381, 0.0512909451415485, 
    0.0531033220348709, 0.0523419434600547, 0.0491226580769091, 
    0.042815242398807, 0.0251344860819448, -0.0106974230156285, 
    -0.0464290607270087, -0.0703531404088194, -0.0829696615292754, 
    -0.0879829606723699, -0.0849820044052567, -0.0664676609190502, 
    -0.066816196379815, -0.0912528028655224, -0.112335948877433, 
    -0.117841795872043, -0.112094695851487, -0.112365562938875, 
    -0.117416296937257, -0.101399547712701, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.000549413403575833, 0.0138609343445309, 0.0293051230072199, 
    0.0434423511258199, 0.0492505974095411, 0.0391348334754192, 
    0.0326000669741209, 0.041375724757685, 0.0524933186235031, 
    0.0568264131478829, 0.0586226933710933, 0.0584015138581848, 
    0.0486168514212155, 0.0185333193214535, -0.0208504538091393, 
    -0.0545007944600646, -0.0744995564947189, -0.083042671104751, 
    -0.0884479815844762, -0.0815191512872689, -0.0567439001625589, 
    -0.0464190321529428, -0.0685880556474294, -0.0970878370968973, 
    -0.116470769953759, -0.11125103986204, -0.107146443499163, 
    -0.107734984193917, -0.0900862578823609, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -0.000876824315086877, 0.0184191179063555, 0.0366147834523258, 
    0.0597513339682559, 0.0811154171009781, 0.0824719065443709, 
    0.068219984509954, 0.0667619131238099, 0.0679973826289001, 
    0.0665049594638282, 0.0667066151660691, 0.0728867220861705, 
    0.0648733848833199, 0.0359379160798853, 0.000947824916362721, 
    -0.0290463858603658, -0.0479658190692731, -0.0611186895472386, 
    -0.0759880061222724, -0.0703052832211533, -0.0452347766180581, 
    -0.0308019555296719, -0.0465363580004904, -0.0841875112703651, 
    -0.114736665118155, -0.109855955012029, -0.103130669530014, 
    -0.102590774878042, -0.0901073361978885, -0.0806119540481011, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -0.00118820883482688, 0.0225439225637645, 0.0447624185341323, 
    0.0722294712357344, 0.105443968173031, 0.117350375095603, 
    0.108646575425693, 0.0990660684033909, 0.0922518941050821, 
    0.0831501613870996, 0.0726029202871983, 0.0746793192477183, 
    0.0733496971151509, 0.0579038244643112, 0.0287612117916655, 
    0.00537749880565302, -0.0120282654702272, -0.0287586590129561, 
    -0.0419932308615047, -0.0466667808257572, -0.03766796970701, 
    -0.0340371624202405, -0.0461779106610422, -0.0806263957250813, 
    -0.112904669345683, -0.104043829266395, -0.091294951177527, 
    -0.0926371027537021, -0.0878042506725705, -0.0832726963498247, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0.000629079264515328, 0.0304170494650356, 0.052253864726093, 
    0.0868938127754851, 0.127443801584721, 0.139605598688566, 
    0.130984557944003, 0.113964980822322, 0.108666300340532, 
    0.101119096481942, 0.0814209149961576, 0.0745617747154559, 
    0.0753460507688637, 0.0694149995322673, 0.0544686395616101, 
    0.0435634574557569, 0.0270829353593203, -0.00120682672081296, 
    -0.018243109668247, -0.0342946909183698, -0.0389879251153562, 
    -0.0491828841674305, -0.0593668796594108, -0.0749259681635426, 
    -0.0999079183305026, -0.0973327830276976, -0.0778732025489182, 
    -0.0703591329365266, -0.0660276862757552, -0.0664267582255328, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -0.000562106433904667, 0.0294077816186364, 0.0482965725881777, 
    0.0717816069459196, 0.116707746623828, 0.147141928524773, 
    0.141001724573239, 0.121410086615623, 0.106961411628842, 
    0.100444672598078, 0.0864554329741946, 0.0762903819572552, 
    0.0786219436619214, 0.0781055150509287, 0.073511041964524, 
    0.063027105525086, 0.0363170027048443, 0.00339439424059892, 
    -0.0289992626021552, -0.0562495860640902, -0.0721628661072471, 
    -0.0774491377917552, -0.0759091005612113, -0.0709761772827546, 
    -0.0884615505517034, -0.0917767262085756, -0.0710579697249469, 
    -0.051883503574568, -0.0441515048830867, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -0.00515938828841622, 0.0207802220775177, 0.0313138339946233, 
    0.0376733297524155, 0.0754994411075659, 0.113462471532008, 
    0.117433674746804, 0.0999332287378798, 0.0940530429809903, 
    0.0913371222965744, 0.0805575738013964, 0.080741876746733, 
    0.0824828693182588, 0.074493288795708, 0.0706207492865304, 
    0.0492061712027163, 0.017418618326578, -0.0198245609800642, 
    -0.0620528707414752, -0.0898683339345375, -0.0987112556462041, 
    -0.0916459155503711, -0.081209592565862, -0.0717763152395592, 
    -0.0770350319672291, -0.079790368006404, -0.0655362840804696, 
    -0.0426681852151886, -0.0351647935953923, -0.0319071726111181, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -0.00741108389302793, 0.00936148239752364, 0.0116995657222536, 
    0.0184743056670131, 0.0547803644516232, 0.0810622194187508, 
    0.0785108159469786, 0.0718915477681151, 0.0741893332370187, 
    0.0776152454440016, 0.0754666692177693, 0.0722517190980384, 
    0.0771872469036056, 0.0659442722101405, 0.0417834207252167, 
    0.0152952828654711, -0.00294919290626485, -0.0161478508657198, 
    -0.0410147965141071, -0.0661893091647466, -0.0836431558726858, 
    -0.0772788113771145, -0.0714135154199889, -0.0656840782406646, 
    -0.0652653459610868, -0.0672794224452877, -0.0534949720162833, 
    -0.0334050807146055, -0.0291444289276469, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -0.00903961380076852, 0.00959501453945472, 0.0141885996775922, 
    0.0252057492371473, 0.0483265945898977, 0.0557482848733261, 
    0.0404982701224332, 0.0292341610699337, 0.0458721571847184, 
    0.0687511529242586, 0.062644171807079, 0.0528826462062893, 
    0.0550814473043108, 0.0436319778114815, 0.0079265607792675, 
    -0.0280333325635298, -0.0413364807324819, -0.0324454360795945, 
    -0.0242528018246714, -0.0328580002789255, -0.0502618883310723, 
    -0.0538272354129217, -0.059443926838633, -0.0541937433912064, 
    -0.0600719734132172, -0.0537170660274214, -0.0376546802154042, 
    -0.0247436239978787, -0.0208023087195037, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, -0.0150058031980528, -0.00791455762793496, -0.00744375992627161, 
    -0.00648697130899449, -0.00348564642342225, 0.000585014042302609, 
    -0.00287379197731653, -0.0133566488132648, -0.00662508212875247, 
    0.00751693122207849, 0.00983396005271965, 0.00419750382918283, 
    0.00423149456758387, 0.00502853692378617, -0.00230684182027245, 
    -0.0151533588345881, -0.0208173528202563, -0.0190509312186965, 
    -0.0179400522941304, -0.0187057308728579, -0.0169393832710783, 
    -0.0152147696713086, -0.0199590352510198, -0.0212481737277574, 
    -0.0234737154708985, -0.0203518798740792, -0.01286454294699, 
    -0.00717481671404735, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0 ;

 obs_depth = 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 29.2668575128976, 28.2931106880205, 
    27.4265565482546, 26.5039098414807, 24.423812685455, 23.3385752962144, 
    22.4948155714326, 21.4820027503705, 19.5909409766348, 18.5006832413942, 
    17.5652301596557, 16.5915422979033, 15.5603081578148, 14.5668286869143, 
    13.5724111828824, 12.5531948612262, 11.623666106713, 25.5704522143069, 
    20.66053580274, 29.2668575128976, 28.2931106880205, 27.4265565482546, 
    26.5039098414807, 24.423812685455, 23.3385752962144, 22.4948155714326, 
    21.4820027503705, 19.5909409766348, 18.5006832413942, 17.5652301596557, 
    16.5915422979033, 15.5603081578148, 14.5668286869143, 13.5724111828824, 
    12.5531948612262, 11.623666106713, 25.5704522143069, 20.66053580274, 
    29.1765930075953, 28.2006231286159, 27.3146042719267, 26.3481835357321, 
    25.4044519671984, 24.2381525822845, 23.1385108926005, 22.2941270709058, 
    21.5922015041614, 20.7078648990055, 19.5771362306175, 18.6068110796689, 
    17.6085979442171, 16.5775260280661, 15.4903276058566, 14.4401065754562, 
    13.5199418220692, 12.5752364248567, 11.4483834094807, 10.7162619835978, 
    29.1765930075953, 28.2006231286159, 27.3146042719267, 26.3481835357321, 
    25.4044519671984, 24.2381525822845, 23.1385108926005, 22.2941270709058, 
    21.5922015041614, 20.7078648990055, 19.5771362306175, 18.6068110796689, 
    17.6085979442171, 16.5775260280661, 15.4903276058566, 14.4401065754562, 
    13.5199418220692, 12.5752364248567, 11.4483834094807, 10.7162619835978, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 28.497942925279, 26.8672133975361, 25.7129072256134, 
    24.4366222221351, 23.4392429305181, 22.6538281968931, 21.6140740635757, 
    20.478584858072, 19.4404560056958, 18.4761277049908, 17.452493216506, 
    16.4583249953704, 15.607440036457, 14.7026758073398, 13.5822394262558, 
    12.4266717533476, 11.622671244914, 10.7970234065745, 9.50682217279063, 
    8.223448811319, 7.42083701055481, 6.6473812181214, 5.92611469679479, 
    28.497942925279, 26.8672133975361, 25.7129072256134, 24.4366222221351, 
    23.4392429305181, 22.6538281968931, 21.6140740635757, 20.478584858072, 
    19.4404560056958, 18.4761277049908, 17.452493216506, 16.4583249953704, 
    15.607440036457, 14.7026758073398, 13.5822394262558, 12.4266717533476, 
    11.622671244914, 10.7970234065745, 9.50682217279063, 8.223448811319, 
    7.42083701055481, 6.6473812181214, 5.92611469679479, 29.5194516493063, 
    28.5582946049245, 27.4108598597076, 26.4988476150163, 25.7405626789316, 
    24.7425589011678, 23.542568637073, 22.4113051531266, 21.5287880368751, 
    20.4720596262526, 19.6083439038047, 18.4643809131208, 17.4508813552931, 
    16.5446768113607, 15.5292117520068, 14.5494420567707, 13.5711432106657, 
    12.5626158316309, 11.5145888879628, 10.4180809638348, 9.48128195320091, 
    8.55472553700606, 7.83020373649257, 29.5194516493063, 28.5582946049245, 
    27.4108598597076, 26.4988476150163, 25.7405626789316, 24.7425589011678, 
    23.542568637073, 22.4113051531266, 21.5287880368751, 20.4720596262526, 
    19.6083439038047, 18.4643809131208, 17.4508813552931, 16.5446768113607, 
    15.5292117520068, 14.5494420567707, 13.5711432106657, 12.5626158316309, 
    11.5145888879628, 10.4180809638348, 9.48128195320091, 8.55472553700606, 
    7.83020373649257, 14.2689979780551, 9.80039242473299, 5.43671013393478, 
    27.4934257345086, 25.0633778892587, 23.2306492782743, 21.942642182963, 
    20.959151070739, 19.6070869399149, 18.071523939678, 16.3763420228374, 
    12.1315549015429, 7.45892315102195, 3.79940525580201, 2.5300881915662, 
    1.87581273183135, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 18.4689380153097, 26.8995934164539, 24.2643706312457, 
    22.3152597273092, 20.9584439536121, 19.9255863779856, 16.7701234354496, 
    14.742514807653, 8.82349156434568, 3.73425553800546, 11.9312521281224, 
    5.93909991295722, 2.03862534607762, 12.5203876949826, 6.80019426494749, 
    2.73974882827024, 15.135895876409, 9.64929540266797, 4.50509399197809, 
    1.35111636950138, 27.0242568463261, 24.4545506234755, 22.5262260215658, 
    21.1910920075557, 20.1661447299387, 17.0699949113717, 18.7247264689812, 
    28.7161612298962, 23.6721469892783, 20.9510541403711, 17.9068920995421, 
    15.601300155688, 13.5326890324778, 11.2924797492445, 28.7161612298962, 
    23.6721469892783, 20.9510541403711, 17.9068920995421, 15.601300155688, 
    13.5326890324778, 11.2924797492445, 27.6410529895551, 22.2708069912956, 
    19.3702405519766, 17.3850930789866, 15.7910968375277, 14.2732865119821, 
    11.8926434596387, 7.25410636362123, 2.64189350702765, 27.6410529895551, 
    22.2708069912956, 19.3702405519766, 17.3850930789866, 15.7910968375277, 
    14.2732865119821, 11.8926434596387, 7.25410636362123, 2.64189350702765, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 28.7735790246829, 
    23.0855182855433, 20.506091871842, 18.7392589766159, 17.3460545527911, 
    15.0037141121633, 12.1390236056492, 7.7703533271696, 2.05406206156723, 
    28.7735790246829, 23.0855182855433, 20.506091871842, 18.7392589766159, 
    17.3460545527911, 15.0037141121633, 12.1390236056492, 7.7703533271696, 
    2.05406206156723, 27.5892905279705, 23.8945051304732, 22.4844917818553, 
    21.3376579586492, 20.4633904430287, 19.3777085361571, 17.8264841802613, 
    16.088786419746, 13.8008164291014, 11.8528899502112, 9.97484218427245, 
    7.60465261531815, 5.17551143723144, 3.3097549891584, 1.48774566301297, 
    27.5892905279705, 23.8945051304732, 22.4844917818553, 21.3376579586492, 
    20.4633904430287, 19.3777085361571, 17.8264841802613, 16.088786419746, 
    13.8008164291014, 11.8528899502112, 9.97484218427245, 7.60465261531815, 
    5.17551143723144, 3.3097549891584, 1.48774566301297, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30 ;

 obs_Xgrid = 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.8999938964843, 12.8999938964843, 12.8999938964843, 12.8999938964843, 
    12.8999938964843, 12.8999938964843, 12.8999938964843, 12.8999938964843, 
    12.8999938964843, 12.8999938964843, 12.8999938964843, 12.8999938964843, 
    12.8999938964843, 12.8999938964843, 12.8999938964843, 12.8999938964843, 
    12.8999938964843, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 14.1000061035157, 
    14.1000061035157, 14.1000061035157, 14.1000061035157, 14.1000061035157, 
    14.1000061035157, 14.1000061035157, 14.1000061035157, 14.1000061035157, 
    14.1000061035157, 14.1000061035157, 14.1000061035157, 14.1000061035157, 
    14.1000061035157, 14.1000061035157, 14.1000061035157, 14.1000061035157, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 15, 15, 15, 15, 15, 15, 15, 15, 15, 
    15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 
    15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 
    15, 15, 15, 15, 15, 15, 15.8999938964843, 15.8999938964843, 
    15.8999938964843, 15.8999938964843, 15.8999938964843, 15.8999938964843, 
    15.8999938964843, 15.8999938964843, 15.8999938964843, 15.8999938964843, 
    15.8999938964843, 15.8999938964843, 15.8999938964843, 15.8999938964843, 
    15.8999938964843, 15.8999938964843, 15.8999938964843, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 17.1000061035157, 17.1000061035157, 17.1000061035157, 
    17.1000061035157, 17.1000061035157, 17.1000061035157, 17.1000061035157, 
    17.1000061035157, 17.1000061035157, 17.1000061035157, 17.1000061035157, 
    17.1000061035157, 17.1000061035157, 17.1000061035157, 17.1000061035157, 
    17.1000061035157, 17.1000061035157, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 
    18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 
    18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 
    18.8999938964844, 18.8999938964844, 18.8999938964844, 18.8999938964844, 
    18.8999938964844, 18.8999938964844, 18.8999938964844, 18.8999938964844, 
    18.8999938964844, 18.8999938964844, 18.8999938964844, 18.8999938964844, 
    18.8999938964844, 18.8999938964844, 18.8999938964844, 18.8999938964844, 
    18.8999938964844, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 20.1000061035156, 
    20.1000061035156, 20.1000061035156, 20.1000061035156, 20.1000061035156, 
    20.1000061035156, 20.1000061035156, 20.1000061035156, 20.1000061035156, 
    20.1000061035156, 20.1000061035156, 20.1000061035156, 20.1000061035156, 
    20.1000061035156, 20.1000061035156, 20.1000061035156, 20.1000061035156, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 21, 21, 21, 21, 21, 21, 21, 21, 21, 
    21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 
    21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 
    21, 21, 21, 21, 21, 21, 21.8999938964844, 21.8999938964844, 
    21.8999938964844, 21.8999938964844, 21.8999938964844, 21.8999938964844, 
    21.8999938964844, 21.8999938964844, 21.8999938964844, 21.8999938964844, 
    21.8999938964844, 21.8999938964844, 21.8999938964844, 21.8999938964844, 
    21.8999938964844, 21.8999938964844, 21.8999938964844, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 23.1000061035156, 23.1000061035156, 23.1000061035156, 
    23.1000061035156, 23.1000061035156, 23.1000061035156, 23.1000061035156, 
    23.1000061035156, 23.1000061035156, 23.1000061035156, 23.1000061035156, 
    23.1000061035156, 23.1000061035156, 23.1000061035156, 23.1000061035156, 
    23.1000061035156, 23.1000061035156, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 
    24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 
    24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 
    24.8999938964844, 24.8999938964844, 24.8999938964844, 24.8999938964844, 
    24.8999938964844, 24.8999938964844, 24.8999938964844, 24.8999938964844, 
    24.8999938964844, 24.8999938964844, 24.8999938964844, 24.8999938964844, 
    24.8999938964844, 24.8999938964844, 24.8999938964844, 24.8999938964844, 
    24.8999938964844, 25.0499954223633, 25.0499954223633, 25.0499954223633, 
    25.0499954223633, 25.0499954223633, 25.0499954223633, 25.0499954223633, 
    25.0499954223633, 25.0499954223633, 25.0499954223633, 25.0499954223633, 
    25.0499954223633, 25.0499954223633, 25.0499954223633, 25.0499954223633, 
    25.0499954223633, 25.0499954223633, 25.0363603071733, 25.0499954223633, 
    25.1571350097656, 25.5, 25.1142817905971, 25.1399963378906, 
    25.1624965667725, 25.0499954223633, 24.75, 24.8571428571429, 
    25.0499954223633, 24.9899963378906, 25.0499954223633, 25.0363603071733, 
    25.0363603071733, 25.0090859153054, 25.0499954223633, 26.1000061035156, 
    26.1000061035156, 26.1000061035156, 26.1000061035156, 26.1000061035156, 
    26.1000061035156, 26.1000061035156, 26.1000061035156, 26.1000061035156, 
    26.1000061035156, 26.1000061035156, 26.1000061035156, 26.1000061035156, 
    26.1000061035156, 26.1000061035156, 26.1000061035156, 26.1000061035156, 
    25.9500045776367, 25.9500045776367, 25.9500045776367, 25.9500045776367, 
    25.9500045776367, 25.9500045776367, 25.9500045776367, 25.9500045776367, 
    25.9500045776367, 25.9500045776367, 25.9500045776367, 25.9500045776367, 
    25.9500045776367, 25.9500045776367, 25.9500045776367, 25.9500045776367, 
    25.9636396928267, 25.9500045776367, 25.9500045776367, 25.8600036621094, 
    26.057144165039, 25.9800064086914, 25.6000061035156, 25.7500076293945, 
    25.7625045776367, 25.9500045776367, 25.8000052315848, 26.0100036621094, 
    25.9500045776367, 25.9500045776367, 25.5750045776367, 26.040005493164, 
    27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 
    27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 26.8999938964844, 
    27, 27, 26.9499969482422, 27.0857195172991, 26.9249954223633, 
    26.7999877929688, 27.3000183105469, 27.0500030517578, 26.6999816894531, 
    27.1500091552734, 27.0600036621094, 27.1000061035156, 27, 27, 27, 
    27.0375022888184, 27, 27, 27.8999938964844, 27.8999938964844, 
    27.8999938964844, 27.8999938964844, 27.8999938964844, 27.8999938964844, 
    27.8999938964844, 27.8999938964844, 27.8999938964844, 27.8999938964844, 
    27.8999938964844, 27.8999938964844, 27.8999938964844, 27.8999938964844, 
    27.8999938964844, 27.8999938964844, 27.8999938964844, 28.0499954223633, 
    28.0499954223633, 28.0499954223633, 28.0499954223633, 28.0499954223633, 
    28.0499954223633, 28.0499954223633, 28.0499954223633, 28.0499954223633, 
    28.0499954223633, 28.0499954223633, 28.0499954223633, 28.0499954223633, 
    28.0333302815755, 28.0499954223633, 28.2, 28.0090859153054, 
    28.0333302815755, 28.1142817905971, 27.8571363176618, 27.5999908447266, 
    27.75, 28.1999931335449, 27.999994913737, 28.0999959309896, 
    28.0499954223633, 28.0499954223633, 28.0499954223633, 28.0499954223633, 
    28.0499954223633, 28.0499954223633, 29.1000061035156, 29.1000061035156, 
    29.1000061035156, 29.1000061035156, 29.1000061035156, 29.1000061035156, 
    29.1000061035156, 29.1000061035156, 29.1000061035156, 29.1000061035156, 
    29.1000061035156, 29.1000061035156, 29.1000061035156, 29.1000061035156, 
    29.1000061035156, 29.1000061035156, 29.1000061035156, 28.9500045776367, 
    28.9500045776367, 28.9500045776367, 28.9500045776367, 28.9500045776367, 
    28.9500045776367, 28.9500045776367, 28.9500045776367, 28.9500045776367, 
    28.9500045776367, 28.9500045776367, 28.9500045776367, 28.7400054931641, 
    28.8000030517578, 28.9090950705788, 28.8000052315848, 28.7571454729352, 
    29.0999908447265, 28.6000061035156, 28.8750057220459, 28.9090950705788, 
    28.9500045776367, 28.9500045776367, 28.9500045776367, 28.9500045776367, 
    28.9090950705788, 28.7625045776367, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 29.8799926757813, 29.8499908447266, 29.8499908447266, 
    29.6999816894531, 30.8999938964844, 30.8999938964844, 30.8999938964844, 
    30.8999938964844, 30.8999938964844, 30.8999938964844, 30.8999938964844, 
    30.8999938964844, 30.8999938964844, 30.8999938964844, 30.8999938964844, 
    30.8999938964844, 30.8999938964844, 30.8999938964844, 30.8999938964844, 
    30.8999938964844, 30.8999938964844, 31.0499954223633, 31.0499954223633, 
    31.0499954223633, 31.0499954223633, 31.0499954223633, 31.0499954223633, 
    31.0499954223633, 31.0090859153054, 32.1000061035156, 32.1000061035156, 
    32.1000061035156, 32.1000061035156, 32.1000061035156, 32.1000061035156, 
    32.1000061035156, 32.1000061035156, 32.1000061035156, 32.1000061035156, 
    32.1000061035156, 32.1000061035156, 32.1000061035156, 32.1000061035156, 
    32.1000061035156, 32.1000061035156, 32.1000061035156, 31.9500045776367, 
    31.9500045776367, 31.9500045776367, 31.9500045776367, 31.9500045776367, 
    31.9500045776367, 31.9500045776367, 33, 33, 33, 33, 33, 33, 33, 33, 33, 
    33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33.8999938964844, 
    33.8999938964844, 33.8999938964844, 33.8999938964844, 33.8999938964844, 
    33.8999938964844, 33.8999938964844, 33.8999938964844, 33.8999938964844, 
    33.8999938964844, 33.8999938964844, 33.8999938964844, 33.8999938964844, 
    33.8999938964844, 33.8999938964844, 33.8999938964844, 33.8999938964844, 
    34.0499954223633, 34.0499954223633, 34.0499954223633, 34.0499954223633, 
    33.959994506836, 35.1000061035156, 35.1000061035156, 35.1000061035156, 
    35.1000061035156, 35.1000061035156, 35.1000061035156, 35.1000061035156, 
    35.1000061035156, 35.1000061035156, 35.1000061035156, 35.1000061035156, 
    35.1000061035156, 35.1000061035156, 35.1000061035156, 35.1000061035156, 
    35.1000061035156, 35.1000061035156, 34.9500045776367, 34.9500045776367, 
    34.9090950705788, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 
    36, 36, 36, 35.9624977111816, 35.9624977111816, 36.8999938964844, 
    36.8999938964844, 36.8999938964844, 36.8999938964844, 36.8999938964844, 
    36.8999938964844, 36.8999938964844, 36.8999938964844, 36.8999938964844, 
    36.8999938964844, 36.8999938964844, 36.8999938964844, 36.8999938964844, 
    36.8999938964844, 36.8999938964844, 36.8999938964844, 36.8624954223633, 
    38.1000061035156, 38.1000061035156, 38.1000061035156, 38.1000061035156, 
    38.1000061035156, 38.1000061035156, 38.1000061035156, 38.1000061035156, 
    38.1000061035156, 38.1000061035156, 38.1000061035156, 38.1000061035156, 
    38.1000061035156, 38.1000061035156, 38.1000061035156, 37.9800109863281, 
    39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 
    39.8999938964844, 39.8999938964844, 39.8999938964844, 39.8999938964844, 
    39.8999938964844, 39.8999938964844, 39.8999938964844, 39.8999938964844, 
    39.8999938964844, 39.8999938964844, 39.8999938964844, 39.8999938964844, 
    39.75, 39.75, 41.1000061035156, 41.1000061035156, 41.1000061035156, 
    41.1000061035156, 41.1000061035156, 41.1000061035156, 41.1000061035156, 
    41.1000061035156, 41.1000061035156, 41.1000061035156, 41.0625057220459, 
    41.1000061035156, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 
    42.0375022888184, 42, 42.8999938964844, 42.8999938964844, 
    42.8999938964844, 42.8999938964844, 42.8999938964844, 42.8999938964844, 
    42.8999938964844, 42.8999938964844, 42.8999938964844, 42.8999938964844, 
    42.8999938964844, 42.8999938964844, 44.1000061035156, 44.1000061035156, 
    44.1000061035156, 44.1000061035156, 44.1000061035156, 44.1000061035156, 
    44.1000061035156, 44.1000061035156, 44.1000061035156, 44.1000061035156, 
    44.1000061035156, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 
    45.8999938964844, 45.8999938964844, 45.8999938964844, 45.8999938964844, 
    45.8999938964844, 45.8999938964844, 45.8999938964844, 45.8999938964844, 
    45.8999938964844, 45.8999938964844, 45.8999938964844, 47.1000061035156, 
    47.1000061035156, 47.1000061035156, 47.1000061035156, 47.1000061035156, 
    47.1000061035156, 47.1000061035156, 47.1000061035156, 47.1375045776367, 
    47.1000061035156, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48.8999938964844, 
    48.8999938964844, 48.8999938964844, 48.8999938964844, 48.8999938964844, 
    48.8999938964844, 48.8999938964844, 48.8999938964844, 48.8624954223633, 
    50.1000061035156, 50.1000061035156, 50.1000061035156, 50.1000061035156, 
    50.1000061035156, 50.1000061035156, 50.0142909458706, 49.9200073242188, 
    51, 51, 51, 51, 51, 51.8999938964844, 51.8999938964844, 51.8999938964844, 
    51.75, 17.1239776611328, 17.1239776611328, 17.1239776611328, 
    17.1239776611328, 17.1239776611328, 17.1239776611328, 17.1239776611328, 
    17.1239776611328, 17.1239776611328, 17.1239776611328, 17.1239776611328, 
    17.1239776611328, 17.1239776611328, 17.1239776611328, 17.1239776611328, 
    17.1239776611328, 17.1239776611328, 17.1239776611328, 17.1239776611328, 
    17.1239776611328, 17.1239776611328, 17.1239776611328, 17.1239776611328, 
    17.1239776611328, 17.1239776611328, 17.1239776611328, 17.1239776611328, 
    17.1239776611328, 17.1239776611328, 17.1239776611328, 17.1239776611328, 
    17.1239776611328, 17.1239776611328, 17.1239776611328, 17.1239776611328, 
    17.1239776611328, 17.1239776611328, 17.1239776611328, 20.4299926757812, 
    20.4299926757812, 20.4299926757812, 20.4299926757812, 20.4299926757812, 
    20.4299926757812, 20.4299926757812, 20.4299926757812, 20.4299926757812, 
    20.4299926757812, 20.4299926757812, 20.4299926757812, 20.4299926757812, 
    20.4299926757812, 20.4299926757812, 20.4299926757812, 20.4299926757812, 
    20.4299926757812, 20.4299926757812, 20.4299926757812, 20.4299926757812, 
    20.4299926757812, 20.4299926757812, 20.4299926757812, 20.4299926757812, 
    20.4299926757812, 20.4299926757812, 20.4299926757812, 20.4299926757812, 
    20.4299926757812, 20.4299926757812, 20.4299926757812, 20.4299926757812, 
    20.4299926757812, 20.4299926757812, 20.4299926757812, 20.4299926757812, 
    20.4299926757812, 20.4299926757812, 20.4299926757812, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.8999938964843, 12.8999938964843, 
    12.8999938964843, 12.8999938964843, 12.8999938964843, 12.8999938964843, 
    12.8999938964843, 12.8999938964843, 12.8999938964843, 12.8999938964843, 
    12.8999938964843, 12.8999938964843, 12.8999938964843, 12.8999938964843, 
    12.8999938964843, 12.8999938964843, 12.8999938964843, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 14.1000061035157, 14.1000061035157, 14.1000061035157, 
    14.1000061035157, 14.1000061035157, 14.1000061035157, 14.1000061035157, 
    14.1000061035157, 14.1000061035157, 14.1000061035157, 14.1000061035157, 
    14.1000061035157, 14.1000061035157, 14.1000061035157, 14.1000061035157, 
    14.1000061035157, 14.1000061035157, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 
    15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 
    15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 
    15.8999938964843, 15.8999938964843, 15.8999938964843, 15.8999938964843, 
    15.8999938964843, 15.8999938964843, 15.8999938964843, 15.8999938964843, 
    15.8999938964843, 15.8999938964843, 15.8999938964843, 15.8999938964843, 
    15.8999938964843, 15.8999938964843, 15.8999938964843, 15.8999938964843, 
    15.8999938964843, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 17.1000061035157, 
    17.1000061035157, 17.1000061035157, 17.1000061035157, 17.1000061035157, 
    17.1000061035157, 17.1000061035157, 17.1000061035157, 17.1000061035157, 
    17.1000061035157, 17.1000061035157, 17.1000061035157, 17.1000061035157, 
    17.1000061035157, 17.1000061035157, 17.1000061035157, 17.1000061035157, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 18, 18, 18, 18, 18, 18, 18, 18, 18, 
    18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 
    18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 
    18, 18, 18, 18, 18, 18, 18.8999938964844, 18.8999938964844, 
    18.8999938964844, 18.8999938964844, 18.8999938964844, 18.8999938964844, 
    18.8999938964844, 18.8999938964844, 18.8999938964844, 18.8999938964844, 
    18.8999938964844, 18.8999938964844, 18.8999938964844, 18.8999938964844, 
    18.8999938964844, 18.8999938964844, 18.8999938964844, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 20.1000061035156, 20.1000061035156, 20.1000061035156, 
    20.1000061035156, 20.1000061035156, 20.1000061035156, 20.1000061035156, 
    20.1000061035156, 20.1000061035156, 20.1000061035156, 20.1000061035156, 
    20.1000061035156, 20.1000061035156, 20.1000061035156, 20.1000061035156, 
    20.1000061035156, 20.1000061035156, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 
    21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 
    21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 
    21.8999938964844, 21.8999938964844, 21.8999938964844, 21.8999938964844, 
    21.8999938964844, 21.8999938964844, 21.8999938964844, 21.8999938964844, 
    21.8999938964844, 21.8999938964844, 21.8999938964844, 21.8999938964844, 
    21.8999938964844, 21.8999938964844, 21.8999938964844, 21.8999938964844, 
    21.8999938964844, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 23.1000061035156, 
    23.1000061035156, 23.1000061035156, 23.1000061035156, 23.1000061035156, 
    23.1000061035156, 23.1000061035156, 23.1000061035156, 23.1000061035156, 
    23.1000061035156, 23.1000061035156, 23.1000061035156, 23.1000061035156, 
    23.1000061035156, 23.1000061035156, 23.1000061035156, 23.1000061035156, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 24, 24, 24, 24, 24, 24, 24, 24, 24, 
    24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 
    24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 
    24, 24, 24, 24, 24, 24, 24.8999938964844, 24.8999938964844, 
    24.8999938964844, 24.8999938964844, 24.8999938964844, 24.8999938964844, 
    24.8999938964844, 24.8999938964844, 24.8999938964844, 24.8999938964844, 
    24.8999938964844, 24.8999938964844, 24.8999938964844, 24.8999938964844, 
    24.8999938964844, 24.8999938964844, 24.8999938964844, 25.0499954223633, 
    25.0499954223633, 25.0499954223633, 25.0499954223633, 25.0499954223633, 
    25.0499954223633, 25.0499954223633, 25.0499954223633, 25.0499954223633, 
    25.0499954223633, 25.0499954223633, 25.0499954223633, 25.0499954223633, 
    25.0499954223633, 25.0499954223633, 25.0499954223633, 25.0499954223633, 
    25.0363603071733, 25.0499954223633, 25.1571350097656, 25.5, 25.125, 
    25.1399963378906, 25.1624965667725, 25.0499954223633, 24.75, 
    24.8571428571429, 25.0499954223633, 24.9899963378906, 25.0499954223633, 
    25.0363603071733, 24.9899963378906, 25.0090859153054, 25.0499954223633, 
    26.1000061035156, 26.1000061035156, 26.1000061035156, 26.1000061035156, 
    26.1000061035156, 26.1000061035156, 26.1000061035156, 26.1000061035156, 
    26.1000061035156, 26.1000061035156, 26.1000061035156, 26.1000061035156, 
    26.1000061035156, 26.1000061035156, 26.1000061035156, 26.1000061035156, 
    26.1000061035156, 25.9500045776367, 25.9500045776367, 25.9500045776367, 
    25.9500045776367, 25.9500045776367, 25.9500045776367, 25.9500045776367, 
    25.9500045776367, 25.9500045776367, 25.9500045776367, 25.9500045776367, 
    25.9500045776367, 25.9500045776367, 25.9500045776367, 25.9500045776367, 
    25.9500045776367, 25.9636396928267, 25.9500045776367, 25.9500045776367, 
    25.8600036621094, 26.057144165039, 25.9800064086914, 25.6000061035156, 
    25.7500076293945, 25.7625045776367, 25.9500045776367, 25.8000052315848, 
    26.0100036621094, 25.9500045776367, 25.9500045776367, 25.6000061035156, 
    26.040005493164, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 
    27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 
    26.8799926757813, 27, 27, 26.9499969482422, 27.0857195172991, 
    26.9249954223633, 26.7999877929688, 27.3000183105469, 27.0500030517578, 
    26.6999816894531, 27.1500091552734, 27.0600036621094, 27.1000061035156, 
    27, 27, 27, 27.0375022888184, 27, 27, 27.8999938964844, 27.8999938964844, 
    27.8999938964844, 27.8999938964844, 27.8999938964844, 27.8999938964844, 
    27.8999938964844, 27.8999938964844, 27.8999938964844, 27.8999938964844, 
    27.8999938964844, 27.8999938964844, 27.8999938964844, 27.8999938964844, 
    27.8999938964844, 27.8999938964844, 27.8999938964844, 28.0499954223633, 
    28.0499954223633, 28.0499954223633, 28.0499954223633, 28.0499954223633, 
    28.0499954223633, 28.0499954223633, 28.0499954223633, 28.0499954223633, 
    28.0499954223633, 28.0499954223633, 28.0499954223633, 28.0499954223633, 
    28.0333302815755, 28.0499954223633, 28.2, 28.0090859153054, 
    28.0333302815755, 28.1142817905971, 27.8571363176618, 27.5999908447266, 
    27.75, 28.1999931335449, 27.999994913737, 28.0999959309896, 
    28.0499954223633, 28.0499954223633, 28.0499954223633, 28.0499954223633, 
    28.0499954223633, 28.0499954223633, 29.1000061035156, 29.1000061035156, 
    29.1000061035156, 29.1000061035156, 29.1000061035156, 29.1000061035156, 
    29.1000061035156, 29.1000061035156, 29.1000061035156, 29.1000061035156, 
    29.1000061035156, 29.1000061035156, 29.1000061035156, 29.1000061035156, 
    29.1000061035156, 29.1000061035156, 29.1000061035156, 28.9500045776367, 
    28.9500045776367, 28.9500045776367, 28.9500045776367, 28.9500045776367, 
    28.9500045776367, 28.9500045776367, 28.9500045776367, 28.9500045776367, 
    28.9500045776367, 28.9500045776367, 28.9500045776367, 28.7400054931641, 
    28.8000011444092, 28.9090950705788, 28.8000052315848, 28.7571454729352, 
    29.0999908447265, 28.6000061035156, 28.8750057220459, 28.9090950705788, 
    28.9500045776367, 28.9500045776367, 28.9500045776367, 28.9500045776367, 
    28.9090950705788, 28.7625045776367, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 29.8799926757813, 29.8499908447266, 29.8499908447266, 
    29.6999816894531, 30.8999938964844, 30.8999938964844, 30.8999938964844, 
    30.8999938964844, 30.8999938964844, 30.8999938964844, 30.8999938964844, 
    30.8999938964844, 30.8999938964844, 30.8999938964844, 30.8999938964844, 
    30.8999938964844, 30.8999938964844, 30.8999938964844, 30.8999938964844, 
    30.8999938964844, 30.8999938964844, 31.0499954223633, 31.0499954223633, 
    31.0499954223633, 31.0499954223633, 31.0499954223633, 31.0499954223633, 
    31.0499954223633, 31.0090859153054, 32.1000061035156, 32.1000061035156, 
    32.1000061035156, 32.1000061035156, 32.1000061035156, 32.1000061035156, 
    32.1000061035156, 32.1000061035156, 32.1000061035156, 32.1000061035156, 
    32.1000061035156, 32.1000061035156, 32.1000061035156, 32.1000061035156, 
    32.1000061035156, 32.1000061035156, 32.1000061035156, 31.9500045776367, 
    31.9500045776367, 31.9500045776367, 31.9500045776367, 31.9500045776367, 
    31.9500045776367, 31.9500045776367, 33, 33, 33, 33, 33, 33, 33, 33, 33, 
    33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33.8999938964844, 
    33.8999938964844, 33.8999938964844, 33.8999938964844, 33.8999938964844, 
    33.8999938964844, 33.8999938964844, 33.8999938964844, 33.8999938964844, 
    33.8999938964844, 33.8999938964844, 33.8999938964844, 33.8999938964844, 
    33.8999938964844, 33.8999938964844, 33.8999938964844, 33.8999938964844, 
    34.0499954223633, 34.0499954223633, 34.0499954223633, 34.0499954223633, 
    33.959994506836, 35.1000061035156, 35.1000061035156, 35.1000061035156, 
    35.1000061035156, 35.1000061035156, 35.1000061035156, 35.1000061035156, 
    35.1000061035156, 35.1000061035156, 35.1000061035156, 35.1000061035156, 
    35.1000061035156, 35.1000061035156, 35.1000061035156, 35.1000061035156, 
    35.1000061035156, 35.1000061035156, 34.9500045776367, 34.9500045776367, 
    34.9090950705788, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 
    36, 36, 36, 35.9624977111816, 35.9624977111816, 36.8999938964844, 
    36.8999938964844, 36.8999938964844, 36.8999938964844, 36.8999938964844, 
    36.8999938964844, 36.8999938964844, 36.8999938964844, 36.8999938964844, 
    36.8999938964844, 36.8999938964844, 36.8999938964844, 36.8999938964844, 
    36.8999938964844, 36.8999938964844, 36.8999938964844, 36.8624954223633, 
    38.1000061035156, 38.1000061035156, 38.1000061035156, 38.1000061035156, 
    38.1000061035156, 38.1000061035156, 38.1000061035156, 38.1000061035156, 
    38.1000061035156, 38.1000061035156, 38.1000061035156, 38.1000061035156, 
    38.1000061035156, 38.1000061035156, 38.1000061035156, 37.9800109863281, 
    39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 
    39.8999938964844, 39.8999938964844, 39.8999938964844, 39.8999938964844, 
    39.8999938964844, 39.8999938964844, 39.8999938964844, 39.8999938964844, 
    39.8999938964844, 39.8999938964844, 39.8999938964844, 39.8999938964844, 
    39.75, 39.75, 41.1000061035156, 41.1000061035156, 41.1000061035156, 
    41.1000061035156, 41.1000061035156, 41.1000061035156, 41.1000061035156, 
    41.1000061035156, 41.1000061035156, 41.1000061035156, 41.0625057220459, 
    41.1000061035156, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 
    42.0375022888184, 42, 42.8999938964844, 42.8999938964844, 
    42.8999938964844, 42.8999938964844, 42.8999938964844, 42.8999938964844, 
    42.8999938964844, 42.8999938964844, 42.8999938964844, 42.8999938964844, 
    42.8999938964844, 42.8999938964844, 44.1000061035156, 44.1000061035156, 
    44.1000061035156, 44.1000061035156, 44.1000061035156, 44.1000061035156, 
    44.1000061035156, 44.1000061035156, 44.1000061035156, 44.1000061035156, 
    44.1000061035156, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 
    45.8999938964844, 45.8999938964844, 45.8999938964844, 45.8999938964844, 
    45.8999938964844, 45.8999938964844, 45.8999938964844, 45.8999938964844, 
    45.8999938964844, 45.8999938964844, 45.8999938964844, 47.1000061035156, 
    47.1000061035156, 47.1000061035156, 47.1000061035156, 47.1000061035156, 
    47.1000061035156, 47.1000061035156, 47.1000061035156, 47.1375045776367, 
    47.1000061035156, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48.8999938964844, 
    48.8999938964844, 48.8999938964844, 48.8999938964844, 48.8999938964844, 
    48.8999938964844, 48.8999938964844, 48.8999938964844, 48.8624954223633, 
    50.1000061035156, 50.1000061035156, 50.1000061035156, 50.1000061035156, 
    50.1000061035156, 50.1000061035156, 50.0142909458706, 49.9200073242188, 
    51, 51, 51, 51, 51, 51.8999938964844, 51.8999938964844, 51.8999938964844, 
    51.75, 36.1259994506836, 36.1259994506836, 36.1259994506836, 
    36.1259994506836, 36.1259994506836, 36.1259994506836, 36.1259994506836, 
    36.1259994506836, 36.1259994506836, 36.1259994506836, 36.1259994506836, 
    36.1259994506836, 36.1259994506836, 36.1259994506836, 36.1259994506836, 
    36.1259994506836, 36.1259994506836, 36.1259994506836, 36.1259994506836, 
    36.1259994506836, 36.1259994506836, 36.1259994506836, 36.1259994506836, 
    36.1259994506836, 36.1259994506836, 36.1259994506836, 36.1259994506836, 
    36.1259994506836, 36.1259994506836, 36.1259994506836, 36.1259994506836, 
    36.1259994506836, 36.1259994506836, 36.1259994506836, 36.1259994506836, 
    36.1259994506836, 36.1259994506836, 36.1259994506836, 36.1259994506836, 
    36.1259994506836, 36.1259994506836, 36.1259994506836, 36.1259994506836, 
    36.1259994506836, 36.1259994506836, 36.1259994506836, 5.97898864746094, 
    5.97898864746094, 5.97898864746094, 5.97898864746094, 5.97898864746094, 
    5.97898864746094, 5.97898864746094, 5.97898864746094, 5.97898864746094, 
    5.97898864746094, 5.97898864746094, 5.97898864746094, 5.97898864746094, 
    5.97898864746094, 5.97898864746094, 5.97898864746094, 5.97898864746094, 
    5.97898864746094, 5.97898864746094, 5.97898864746094, 5.97898864746094, 
    5.97898864746094, 5.97898864746094, 5.97898864746094, 5.97898864746094, 
    5.97898864746094, 5.97898864746094, 5.97898864746094, 5.97898864746094, 
    5.97898864746094, 5.97898864746094, 5.97898864746094, 5.97898864746094, 
    5.97898864746094, 5.97898864746094, 5.97898864746094, 5.97898864746094, 
    5.97898864746094, 5.97898864746094, 5.97898864746094, 5.97898864746094, 
    5.97898864746094, 5.97898864746094, 5.97898864746094, 5.97898864746094, 
    5.97898864746094, 26.4090042114258, 26.4090042114258, 26.4090042114258, 
    26.4090042114258, 26.4090042114258, 26.4090042114258, 26.4090042114258, 
    26.4090042114258, 26.4090042114258, 26.4090042114258, 26.4090042114258, 
    26.4090042114258, 26.4090042114258, 26.4090042114258, 26.4090042114258, 
    26.4090042114258, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.8999938964843, 12.8999938964843, 12.8999938964843, 12.8999938964843, 
    12.8999938964843, 12.8999938964843, 12.8999938964843, 12.8999938964843, 
    12.8999938964843, 12.8999938964843, 12.8999938964843, 12.8999938964843, 
    12.8999938964843, 12.8999938964843, 12.8999938964843, 12.8999938964843, 
    12.8999938964843, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 14.1000061035157, 
    14.1000061035157, 14.1000061035157, 14.1000061035157, 14.1000061035157, 
    14.1000061035157, 14.1000061035157, 14.1000061035157, 14.1000061035157, 
    14.1000061035157, 14.1000061035157, 14.1000061035157, 14.1000061035157, 
    14.1000061035157, 14.1000061035157, 14.1000061035157, 14.1000061035157, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 15, 15, 15, 15, 15, 15, 15, 15, 15, 
    15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 
    15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 
    15, 15, 15, 15, 15, 15, 15.8999938964843, 15.8999938964843, 
    15.8999938964843, 15.8999938964843, 15.8999938964843, 15.8999938964843, 
    15.8999938964843, 15.8999938964843, 15.8999938964843, 15.8999938964843, 
    15.8999938964843, 15.8999938964843, 15.8999938964843, 15.8999938964843, 
    15.8999938964843, 15.8999938964843, 15.8999938964843, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 17.1000061035157, 17.1000061035157, 17.1000061035157, 
    17.1000061035157, 17.1000061035157, 17.1000061035157, 17.1000061035157, 
    17.1000061035157, 17.1000061035157, 17.1000061035157, 17.1000061035157, 
    17.1000061035157, 17.1000061035157, 17.1000061035157, 17.1000061035157, 
    17.1000061035157, 17.1000061035157, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 
    18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 
    18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 
    18.8999938964844, 18.8999938964844, 18.8999938964844, 18.8999938964844, 
    18.8999938964844, 18.8999938964844, 18.8999938964844, 18.8999938964844, 
    18.8999938964844, 18.8999938964844, 18.8999938964844, 18.8999938964844, 
    18.8999938964844, 18.8999938964844, 18.8999938964844, 18.8999938964844, 
    18.8999938964844, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 20.1000061035156, 
    20.1000061035156, 20.1000061035156, 20.1000061035156, 20.1000061035156, 
    20.1000061035156, 20.1000061035156, 20.1000061035156, 20.1000061035156, 
    20.1000061035156, 20.1000061035156, 20.1000061035156, 20.1000061035156, 
    20.1000061035156, 20.1000061035156, 20.1000061035156, 20.1000061035156, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 21, 21, 21, 21, 21, 21, 21, 21, 21, 
    21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 
    21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 
    21, 21, 21, 21, 21, 21, 21.8999938964844, 21.8999938964844, 
    21.8999938964844, 21.8999938964844, 21.8999938964844, 21.8999938964844, 
    21.8999938964844, 21.8999938964844, 21.8999938964844, 21.8999938964844, 
    21.8999938964844, 21.8999938964844, 21.8999938964844, 21.8999938964844, 
    21.8999938964844, 21.8999938964844, 21.8999938964844, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 23.1000061035156, 23.1000061035156, 23.1000061035156, 
    23.1000061035156, 23.1000061035156, 23.1000061035156, 23.1000061035156, 
    23.1000061035156, 23.1000061035156, 23.1000061035156, 23.1000061035156, 
    23.1000061035156, 23.1000061035156, 23.1000061035156, 23.1000061035156, 
    23.1000061035156, 23.1000061035156, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 
    24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 
    24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 
    24.8999938964844, 24.8999938964844, 24.8999938964844, 24.8999938964844, 
    24.8999938964844, 24.8999938964844, 24.8999938964844, 24.8999938964844, 
    24.8999938964844, 24.8999938964844, 24.8999938964844, 24.8999938964844, 
    24.8999938964844, 24.8999938964844, 24.8999938964844, 24.8999938964844, 
    24.8999938964844, 25.0499954223633, 25.0499954223633, 25.0499954223633, 
    25.0499954223633, 25.0499954223633, 25.0499954223633, 25.0499954223633, 
    25.0499954223633, 25.0499954223633, 25.0499954223633, 25.0499954223633, 
    25.0499954223633, 25.0499954223633, 25.0499954223633, 25.0499954223633, 
    25.0499954223633, 25.0499954223633, 24.9333292643229, 25.0499954223633, 
    25.1999931335449, 25.125, 25.3499908447266, 25.1142817905971, 
    25.0499954223633, 24.75, 24.8571428571429, 24.9899963378906, 
    25.0090859153054, 25.0499954223633, 25.0363603071733, 24.9899963378906, 
    25.0090859153054, 25.0499954223633, 26.1000061035156, 26.1000061035156, 
    26.1000061035156, 26.1000061035156, 26.1000061035156, 26.1000061035156, 
    26.1000061035156, 26.1000061035156, 26.1000061035156, 26.1000061035156, 
    26.1000061035156, 26.1000061035156, 26.1000061035156, 26.1000061035156, 
    26.1000061035156, 26.1000061035156, 26.1000061035156, 25.9500045776367, 
    25.9500045776367, 25.9500045776367, 25.9500045776367, 25.9500045776367, 
    25.9500045776367, 25.9500045776367, 25.9500045776367, 25.9500045776367, 
    25.9500045776367, 25.9500045776367, 25.9500045776367, 25.9500045776367, 
    25.9500045776367, 25.9500045776367, 25.9500045776367, 25.9636396928267, 
    26.0666707356771, 25.9500045776367, 25.8600036621094, 26.1500015258789, 
    25.9800064086914, 25.5, 25.5, 25.7625045776367, 25.6500091552734, 
    25.8500061035156, 26.0100036621094, 25.9500045776367, 25.9500045776367, 
    25.6000061035156, 26.040005493164, 27, 27, 27, 27, 27, 27, 27, 27, 27, 
    27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 
    27, 27, 27, 27, 27, 26.7749862670898, 26.6999816894531, 26.9499969482422, 
    27.1000061035156, 27.0857195172991, 26.9249954223633, 26.7999877929688, 
    27.3000183105469, 27, 26.6999816894531, 27.1500091552734, 27, 
    27.1000061035156, 27, 27, 27, 27, 27, 27, 27.8999938964844, 
    27.8999938964844, 27.8999938964844, 27.8999938964844, 27.8999938964844, 
    27.8999938964844, 27.8999938964844, 27.8999938964844, 27.8999938964844, 
    27.8999938964844, 27.8999938964844, 27.8999938964844, 27.8999938964844, 
    27.8999938964844, 27.8999938964844, 27.8999938964844, 27.8999938964844, 
    28.0499954223633, 28.0499954223633, 28.0499954223633, 28.0499954223633, 
    28.0499954223633, 28.0499954223633, 28.0499954223633, 28.0499954223633, 
    28.0499954223633, 28.0499954223633, 28.0499954223633, 28.0499954223633, 
    28.0636305375533, 28.0333302815755, 28.079997253418, 28.5, 
    27.959994506836, 27.8999938964844, 27.8249931335449, 27.5999908447266, 
    27.75, 28.0499954223633, 28.0499954223633, 28.0999959309896, 
    28.0499954223633, 28.0499954223633, 28.0499954223633, 28.0499954223633, 
    28.0499954223633, 28.0499954223633, 29.1000061035156, 29.1000061035156, 
    29.1000061035156, 29.1000061035156, 29.1000061035156, 29.1000061035156, 
    29.1000061035156, 29.1000061035156, 29.1000061035156, 29.1000061035156, 
    29.1000061035156, 29.1000061035156, 29.1000061035156, 29.1000061035156, 
    29.1000061035156, 29.1000061035156, 29.1000061035156, 28.9500045776367, 
    28.9500045776367, 28.9500045776367, 28.9500045776367, 28.9500045776367, 
    28.9500045776367, 28.9500045776367, 28.9500045776367, 28.9500045776367, 
    28.9500045776367, 28.9500045776367, 28.9500045776367, 28.7400054931641, 
    28.8000011444092, 29.000005086263, 28.9500045776367, 28.6500091552734, 
    28.8750057220459, 28.9090950705788, 28.9500045776367, 28.9500045776367, 
    28.9500045776367, 28.9500045776367, 28.9090950705788, 28.7625045776367, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 29.8799926757813, 
    29.8499908447266, 29.8499908447266, 29.6999816894531, 30.8999938964844, 
    30.8999938964844, 30.8999938964844, 30.8999938964844, 30.8999938964844, 
    30.8999938964844, 30.8999938964844, 30.8999938964844, 30.8999938964844, 
    30.8999938964844, 30.8999938964844, 30.8999938964844, 30.8999938964844, 
    30.8999938964844, 30.8999938964844, 30.8999938964844, 30.8999938964844, 
    31.0499954223633, 31.0499954223633, 31.0499954223633, 31.0499954223633, 
    31.0499954223633, 31.0499954223633, 31.0499954223633, 31.0090859153054, 
    32.1000061035156, 32.1000061035156, 32.1000061035156, 32.1000061035156, 
    32.1000061035156, 32.1000061035156, 32.1000061035156, 32.1000061035156, 
    32.1000061035156, 32.1000061035156, 32.1000061035156, 32.1000061035156, 
    32.1000061035156, 32.1000061035156, 32.1000061035156, 32.1000061035156, 
    32.1000061035156, 31.9500045776367, 31.9500045776367, 31.9500045776367, 
    31.9500045776367, 31.9500045776367, 31.9500045776367, 31.9500045776367, 
    33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 
    33, 33, 33, 33, 33.8999938964844, 33.8999938964844, 33.8999938964844, 
    33.8999938964844, 33.8999938964844, 33.8999938964844, 33.8999938964844, 
    33.8999938964844, 33.8999938964844, 33.8999938964844, 33.8999938964844, 
    33.8999938964844, 33.8999938964844, 33.8999938964844, 33.8999938964844, 
    33.8999938964844, 33.8999938964844, 34.0499954223633, 34.0499954223633, 
    34.0499954223633, 34.0499954223633, 33.959994506836, 35.1000061035156, 
    35.1000061035156, 35.1000061035156, 35.1000061035156, 35.1000061035156, 
    35.1000061035156, 35.1000061035156, 35.1000061035156, 35.1000061035156, 
    35.1000061035156, 35.1000061035156, 35.1000061035156, 35.1000061035156, 
    35.1000061035156, 35.1000061035156, 35.1000061035156, 35.1000061035156, 
    34.9500045776367, 34.9500045776367, 34.9090950705788, 36, 36, 36, 36, 36, 
    36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 35.9624977111816, 
    35.9624977111816, 36.8999938964844, 36.8999938964844, 36.8999938964844, 
    36.8999938964844, 36.8999938964844, 36.8999938964844, 36.8999938964844, 
    36.8999938964844, 36.8999938964844, 36.8999938964844, 36.8999938964844, 
    36.8999938964844, 36.8999938964844, 36.8999938964844, 36.8999938964844, 
    36.8999938964844, 36.8624954223633, 38.1000061035156, 38.1000061035156, 
    38.1000061035156, 38.1000061035156, 38.1000061035156, 38.1000061035156, 
    38.1000061035156, 38.1000061035156, 38.1000061035156, 38.1000061035156, 
    38.1000061035156, 38.1000061035156, 38.1000061035156, 38.1000061035156, 
    38.1000061035156, 37.9800109863281, 39, 39, 39, 39, 39, 39, 39, 39, 39, 
    39, 39, 39, 39, 39, 39, 39.8999938964844, 39.8999938964844, 
    39.8999938964844, 39.8999938964844, 39.8999938964844, 39.8999938964844, 
    39.8999938964844, 39.8999938964844, 39.8999938964844, 39.8999938964844, 
    39.8999938964844, 39.8999938964844, 39.75, 39.75, 41.1000061035156, 
    41.1000061035156, 41.1000061035156, 41.1000061035156, 41.1000061035156, 
    41.1000061035156, 41.1000061035156, 41.1000061035156, 41.1000061035156, 
    41.1000061035156, 41.0625057220459, 41.1000061035156, 42, 42, 42, 42, 42, 
    42, 42, 42, 42, 42, 42.0375022888184, 42, 42.8999938964844, 
    42.8999938964844, 42.8999938964844, 42.8999938964844, 42.8999938964844, 
    42.8999938964844, 42.8999938964844, 42.8999938964844, 42.8999938964844, 
    42.8999938964844, 42.8999938964844, 42.8999938964844, 44.1000061035156, 
    44.1000061035156, 44.1000061035156, 44.1000061035156, 44.1000061035156, 
    44.1000061035156, 44.1000061035156, 44.1000061035156, 44.1000061035156, 
    44.1000061035156, 44.1000061035156, 45, 45, 45, 45, 45, 45, 45, 45, 45, 
    45, 45, 45.8999938964844, 45.8999938964844, 45.8999938964844, 
    45.8999938964844, 45.8999938964844, 45.8999938964844, 45.8999938964844, 
    45.8999938964844, 45.8999938964844, 45.8999938964844, 45.8999938964844, 
    47.1000061035156, 47.1000061035156, 47.1000061035156, 47.1000061035156, 
    47.1000061035156, 47.1000061035156, 47.1000061035156, 47.1000061035156, 
    47.1375045776367, 47.1000061035156, 48, 48, 48, 48, 48, 48, 48, 48, 48, 
    48.8999938964844, 48.8999938964844, 48.8999938964844, 48.8999938964844, 
    48.8999938964844, 48.8999938964844, 48.8999938964844, 48.8999938964844, 
    48.8624954223633, 50.1000061035156, 50.1000061035156, 50.1000061035156, 
    50.1000061035156, 50.1000061035156, 50.1000061035156, 50.0142909458706, 
    49.9200073242188, 51, 51, 51, 51, 51, 51.8999938964844, 51.8999938964844, 
    51.8999938964844, 51.75, 27.5969924926758, 27.5969924926758, 
    27.5969924926758, 27.5969924926758, 27.5969924926758, 27.5969924926758, 
    27.5969924926758, 27.5969924926758, 27.5969924926758, 27.5969924926758, 
    27.5969924926758, 27.5969924926758, 27.5969924926758, 27.7830047607422, 
    27.7830047607422, 27.7830047607422, 27.7830047607422, 27.7830047607422, 
    27.7830047607422, 27.7830047607422, 27.7830047607422, 27.7830047607422, 
    27.7830047607422, 27.7830047607422, 27.7830047607422, 27.7830047607422, 
    27.7830047607422, 50.0909957885742, 50.0909957885742, 50.0909957885742, 
    50.0909957885742, 50.0909957885742, 50.0909957885742, 50.0909957885742, 
    50.0909957885742, 50.0909957885742, 50.0909957885742, 50.0909957885742, 
    50.0909957885742, 50.0909957885742, 50.0909957885742, 49.754997253418, 
    49.754997253418, 49.754997253418, 49.754997253418, 49.754997253418, 
    49.754997253418, 49.754997253418, 49.754997253418, 49.754997253418, 
    49.754997253418, 49.754997253418, 49.754997253418, 49.754997253418, 
    49.754997253418, 49.754997253418, 49.754997253418, 49.754997253418, 
    49.754997253418, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.1500091552734, 12.1500091552734, 12.1500091552734, 12.1500091552734, 
    12.8999938964843, 12.8999938964843, 12.8999938964843, 12.8999938964843, 
    12.8999938964843, 12.8999938964843, 12.8999938964843, 12.8999938964843, 
    12.8999938964843, 12.8999938964843, 12.8999938964843, 12.8999938964843, 
    12.8999938964843, 12.8999938964843, 12.8999938964843, 12.8999938964843, 
    12.8999938964843, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 13.0499954223633, 
    13.0499954223633, 13.0499954223633, 13.0499954223633, 14.1000061035157, 
    14.1000061035157, 14.1000061035157, 14.1000061035157, 14.1000061035157, 
    14.1000061035157, 14.1000061035157, 14.1000061035157, 14.1000061035157, 
    14.1000061035157, 14.1000061035157, 14.1000061035157, 14.1000061035157, 
    14.1000061035157, 14.1000061035157, 14.1000061035157, 14.1000061035157, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 13.9500045776367, 13.9500045776367, 
    13.9500045776367, 13.9500045776367, 15, 15, 15, 15, 15, 15, 15, 15, 15, 
    15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 
    15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 15, 
    15, 15, 15, 15, 15, 15, 15.8999938964843, 15.8999938964843, 
    15.8999938964843, 15.8999938964843, 15.8999938964843, 15.8999938964843, 
    15.8999938964843, 15.8999938964843, 15.8999938964843, 15.8999938964843, 
    15.8999938964843, 15.8999938964843, 15.8999938964843, 15.8999938964843, 
    15.8999938964843, 15.8999938964843, 15.8999938964843, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 16.0499954223633, 16.0499954223633, 16.0499954223633, 
    16.0499954223633, 17.1000061035157, 17.1000061035157, 17.1000061035157, 
    17.1000061035157, 17.1000061035157, 17.1000061035157, 17.1000061035157, 
    17.1000061035157, 17.1000061035157, 17.1000061035157, 17.1000061035157, 
    17.1000061035157, 17.1000061035157, 17.1000061035157, 17.1000061035157, 
    17.1000061035157, 17.1000061035157, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    16.9500045776367, 16.9500045776367, 16.9500045776367, 16.9500045776367, 
    18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 
    18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 
    18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 18, 
    18.8999938964844, 18.8999938964844, 18.8999938964844, 18.8999938964844, 
    18.8999938964844, 18.8999938964844, 18.8999938964844, 18.8999938964844, 
    18.8999938964844, 18.8999938964844, 18.8999938964844, 18.8999938964844, 
    18.8999938964844, 18.8999938964844, 18.8999938964844, 18.8999938964844, 
    18.8999938964844, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 19.0499954223633, 
    19.0499954223633, 19.0499954223633, 19.0499954223633, 20.1000061035156, 
    20.1000061035156, 20.1000061035156, 20.1000061035156, 20.1000061035156, 
    20.1000061035156, 20.1000061035156, 20.1000061035156, 20.1000061035156, 
    20.1000061035156, 20.1000061035156, 20.1000061035156, 20.1000061035156, 
    20.1000061035156, 20.1000061035156, 20.1000061035156, 20.1000061035156, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 19.9500045776367, 19.9500045776367, 
    19.9500045776367, 19.9500045776367, 21, 21, 21, 21, 21, 21, 21, 21, 21, 
    21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 
    21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 21, 
    21, 21, 21, 21, 21, 21, 21.8999938964844, 21.8999938964844, 
    21.8999938964844, 21.8999938964844, 21.8999938964844, 21.8999938964844, 
    21.8999938964844, 21.8999938964844, 21.8999938964844, 21.8999938964844, 
    21.8999938964844, 21.8999938964844, 21.8999938964844, 21.8999938964844, 
    21.8999938964844, 21.8999938964844, 21.8999938964844, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 22.0499954223633, 22.0499954223633, 22.0499954223633, 
    22.0499954223633, 23.1000061035156, 23.1000061035156, 23.1000061035156, 
    23.1000061035156, 23.1000061035156, 23.1000061035156, 23.1000061035156, 
    23.1000061035156, 23.1000061035156, 23.1000061035156, 23.1000061035156, 
    23.1000061035156, 23.1000061035156, 23.1000061035156, 23.1000061035156, 
    23.1000061035156, 23.1000061035156, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    22.9500045776367, 22.9500045776367, 22.9500045776367, 22.9500045776367, 
    24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 
    24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 
    24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 24, 
    24.8999938964844, 24.8999938964844, 24.8999938964844, 24.8999938964844, 
    24.8999938964844, 24.8999938964844, 24.8999938964844, 24.8999938964844, 
    24.8999938964844, 24.8999938964844, 24.8999938964844, 24.8999938964844, 
    24.8999938964844, 24.8999938964844, 24.8999938964844, 24.8999938964844, 
    24.8999938964844, 25.0499954223633, 25.0499954223633, 25.0499954223633, 
    25.0499954223633, 25.0499954223633, 25.0499954223633, 25.0499954223633, 
    25.0499954223633, 25.0499954223633, 25.0499954223633, 25.0363603071733, 
    25.0499954223633, 25.0363603071733, 25.0499954223633, 25.0090859153054, 
    25.0499954223633, 25.0363603071733, 24.942855834961, 25.0499954223633, 
    25.5, 24.75, 24.959994506836, 24.8999977111817, 24.9333292643229, 
    25.0363603071733, 25.0499954223633, 25.0499954223633, 25.0499954223633, 
    25.0499954223633, 25.0499954223633, 26.1000061035156, 26.1000061035156, 
    26.1000061035156, 26.1000061035156, 26.1000061035156, 26.1000061035156, 
    26.1000061035156, 26.1000061035156, 26.1000061035156, 26.1000061035156, 
    26.1000061035156, 26.1000061035156, 26.1000061035156, 26.1000061035156, 
    26.1000061035156, 26.1000061035156, 26.1000061035156, 25.9500045776367, 
    25.9500045776367, 25.9500045776367, 25.9500045776367, 25.9500045776367, 
    25.9500045776367, 25.9500045776367, 25.9500045776367, 25.9500045776367, 
    25.9500045776367, 25.9090950705788, 25.9500045776367, 25.9500045776367, 
    25.9636396928267, 25.8, 25.8000052315848, 25.9125022888183, 
    25.7000122070312, 25.9666697184245, 25.6500091552734, 25.8000068664551, 
    25.9500045776367, 26.0250091552734, 25.9800018310547, 25.9500045776367, 
    25.9500045776367, 25.9500045776367, 25.9500045776367, 25.9500045776367, 
    27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 27, 
    27, 27, 27, 27, 27, 27, 27, 27, 27, 26.9624977111816, 27, 
    26.9142804827009, 26.8799926757813, 26.6999816894531, 26.6999816894531, 
    27, 27.1000061035156, 27, 27, 27, 27, 27, 26.9624977111816, 
    27.8999938964844, 27.8999938964844, 27.8999938964844, 27.8999938964844, 
    27.8999938964844, 27.8999938964844, 27.8999938964844, 27.8999938964844, 
    27.8999938964844, 27.8999938964844, 27.8999938964844, 27.8999938964844, 
    27.8999938964844, 27.8999938964844, 27.8999938964844, 27.8999938964844, 
    27.8999938964844, 28.0499954223633, 28.0499954223633, 28.0499954223633, 
    28.0499954223633, 28.0499954223633, 28.0499954223633, 28.0499954223633, 
    28.0499954223633, 28.0499954223633, 28.0499954223633, 28.0909049294212, 
    28.0090859153054, 28.0874977111817, 28.079997253418, 28.5, 
    27.5999908447266, 28.0499954223633, 28.109994506836, 28.0499954223633, 
    28.0499954223633, 28.0499954223633, 28.0499954223633, 28.0499954223633, 
    28.0499954223633, 29.1000061035156, 29.1000061035156, 29.1000061035156, 
    29.1000061035156, 29.1000061035156, 29.1000061035156, 29.1000061035156, 
    29.1000061035156, 29.1000061035156, 29.1000061035156, 29.1000061035156, 
    29.1000061035156, 29.1000061035156, 29.1000061035156, 29.1000061035156, 
    29.1000061035156, 29.1000061035156, 28.9500045776367, 28.9500045776367, 
    28.9500045776367, 28.9500045776367, 28.9500045776367, 28.9500045776367, 
    28.9500045776367, 28.9500045776367, 28.9500045776367, 28.9500045776367, 
    28.9500045776367, 28.8857182094029, 28.7400054931641, 28.7000045776367, 
    28.5, 28.8750057220459, 28.9090950705788, 28.9500045776367, 
    28.9500045776367, 28.9500045776367, 28.9500045776367, 28.9090950705788, 
    28.7625045776367, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 29.8799926757813, 
    29.8499908447266, 29.8499908447266, 29.6999816894531, 30.8999938964844, 
    30.8999938964844, 30.8999938964844, 30.8999938964844, 30.8999938964844, 
    30.8999938964844, 30.8999938964844, 30.8999938964844, 30.8999938964844, 
    30.8999938964844, 30.8999938964844, 30.8999938964844, 30.8999938964844, 
    30.8999938964844, 30.8999938964844, 30.8999938964844, 30.8999938964844, 
    31.0499954223633, 31.0499954223633, 31.0499954223633, 31.0499954223633, 
    31.0499954223633, 31.0499954223633, 31.0499954223633, 31.0090859153054, 
    32.1000061035156, 32.1000061035156, 32.1000061035156, 32.1000061035156, 
    32.1000061035156, 32.1000061035156, 32.1000061035156, 32.1000061035156, 
    32.1000061035156, 32.1000061035156, 32.1000061035156, 32.1000061035156, 
    32.1000061035156, 32.1000061035156, 32.1000061035156, 32.1000061035156, 
    32.1000061035156, 31.9500045776367, 31.9500045776367, 31.9500045776367, 
    31.9500045776367, 31.9500045776367, 31.9500045776367, 31.9500045776367, 
    33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 
    33, 33, 33, 33, 33.8999938964844, 33.8999938964844, 33.8999938964844, 
    33.8999938964844, 33.8999938964844, 33.8999938964844, 33.8999938964844, 
    33.8999938964844, 33.8999938964844, 33.8999938964844, 33.8999938964844, 
    33.8999938964844, 33.8999938964844, 33.8999938964844, 33.8999938964844, 
    33.8999938964844, 33.8999938964844, 34.0499954223633, 34.0499954223633, 
    34.0499954223633, 34.0499954223633, 33.8999938964844, 35.1000061035156, 
    35.1000061035156, 35.1000061035156, 35.1000061035156, 35.1000061035156, 
    35.1000061035156, 35.1000061035156, 35.1000061035156, 35.1000061035156, 
    35.1000061035156, 35.1000061035156, 35.1000061035156, 35.1000061035156, 
    35.1000061035156, 35.1000061035156, 35.1000061035156, 35.1000061035156, 
    34.9500045776367, 34.9500045776367, 34.9090950705788, 36, 36, 36, 36, 36, 
    36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 35.9624977111816, 
    35.9624977111816, 36.8999938964844, 36.8999938964844, 36.8999938964844, 
    36.8999938964844, 36.8999938964844, 36.8999938964844, 36.8999938964844, 
    36.8999938964844, 36.8999938964844, 36.8999938964844, 36.8999938964844, 
    36.8999938964844, 36.8999938964844, 36.8999938964844, 36.8999938964844, 
    36.8999938964844, 36.8624954223633, 38.1000061035156, 38.1000061035156, 
    38.1000061035156, 38.1000061035156, 38.1000061035156, 38.1000061035156, 
    38.1000061035156, 38.1000061035156, 38.1000061035156, 38.1000061035156, 
    38.1000061035156, 38.1000061035156, 38.1000061035156, 38.1000061035156, 
    38.1000061035156, 37.9800109863281, 39, 39, 39, 39, 39, 39, 39, 39, 39, 
    39, 39, 39, 39, 39, 39, 39.8999938964844, 39.8999938964844, 
    39.8999938964844, 39.8999938964844, 39.8999938964844, 39.8999938964844, 
    39.8999938964844, 39.8999938964844, 39.8999938964844, 39.8999938964844, 
    39.8999938964844, 39.8999938964844, 39.75, 39.75, 41.1000061035156, 
    41.1000061035156, 41.1000061035156, 41.1000061035156, 41.1000061035156, 
    41.1000061035156, 41.1000061035156, 41.1000061035156, 41.1000061035156, 
    41.1000061035156, 41.0625057220459, 41.1000061035156, 42, 42, 42, 42, 42, 
    42, 42, 42, 42, 42, 42.0375022888184, 42, 42.8999938964844, 
    42.8999938964844, 42.8999938964844, 42.8999938964844, 42.8999938964844, 
    42.8999938964844, 42.8999938964844, 42.8999938964844, 42.8999938964844, 
    42.8999938964844, 42.8999938964844, 42.8999938964844, 44.1000061035156, 
    44.1000061035156, 44.1000061035156, 44.1000061035156, 44.1000061035156, 
    44.1000061035156, 44.1000061035156, 44.1000061035156, 44.1000061035156, 
    44.1000061035156, 44.1000061035156, 45, 45, 45, 45, 45, 45, 45, 45, 45, 
    45, 45, 45.8999938964844, 45.8999938964844, 45.8999938964844, 
    45.8999938964844, 45.8999938964844, 45.8999938964844, 45.8999938964844, 
    45.8999938964844, 45.8999938964844, 45.8999938964844, 45.8999938964844, 
    47.1000061035156, 47.1000061035156, 47.1000061035156, 47.1000061035156, 
    47.1000061035156, 47.1000061035156, 47.1000061035156, 47.1000061035156, 
    47.1375045776367, 47.1000061035156, 48, 48, 48, 48, 48, 48, 48, 48, 48, 
    48.8999938964844, 48.8999938964844, 48.8999938964844, 48.8999938964844, 
    48.8999938964844, 48.8999938964844, 48.8999938964844, 48.8999938964844, 
    48.8624954223633, 50.1000061035156, 50.1000061035156, 50.1000061035156, 
    50.1000061035156, 50.1000061035156, 50.1000061035156, 50.0142909458706, 
    49.9200073242188, 51, 51, 51, 51, 51, 51.8999938964844, 51.8999938964844, 
    51.8999938964844, 51.75, 48.375, 48.375, 48.375, 48.375, 48.375, 48.375, 
    48.375, 48.375, 48.375, 48.375, 48.375, 48.375, 48.375, 48.375, 48.375, 
    48.375, 48.375, 48.375, 46.343994140625, 46.343994140625, 
    46.343994140625, 46.343994140625, 46.343994140625, 46.343994140625, 
    46.343994140625, 46.343994140625, 46.343994140625, 46.343994140625, 
    46.343994140625, 46.343994140625, 46.343994140625, 46.343994140625, 
    46.343994140625, 46.343994140625, 46.343994140625, 46.343994140625, 
    46.343994140625, 46.343994140625, 46.343994140625, 46.343994140625, 
    46.343994140625, 46.343994140625, 46.343994140625, 46.343994140625, 
    46.343994140625, 46.343994140625, 46.343994140625, 46.343994140625, 
    2.99999999993187, 3.99999999993179, 2.99999999993187, 4.9999999999317, 
    3.99999999993179, 5.99999999993162, 4.9999999999317, 6.99999999993145, 
    5.99999999993162, 2.99999999993187, 7.99999999993145, 6.99999999993145, 
    3.99999999993179, 8.99999999993127, 2.99999999993187, 7.99999999993145, 
    4.9999999999317, 9.99999999993119, 3.99999999993179, 8.99999999993128, 
    5.99999999993162, 2.99999999993187, 10.9999999999311, 4.9999999999317, 
    9.99999999993119, 6.99999999993145, 3.99999999993179, 11.999999999931, 
    5.99999999993162, 2.99999999993187, 10.9999999999311, 7.99999999993145, 
    4.9999999999317, 12.9999999999308, 6.99999999993145, 3.99999999993179, 
    11.999999999931, 8.99999999993128, 5.99999999993162, 13.9999999999308, 
    2.99999999993187, 7.99999999993145, 4.9999999999317, 12.9999999999308, 
    9.99999999993119, 6.99999999993145, 14.9999999999307, 3.99999999993179, 
    8.99999999993128, 5.99999999993162, 13.9999999999308, 2.99999999993187, 
    10.9999999999311, 7.99999999993145, 15.9999999999306, 4.9999999999317, 
    9.99999999993119, 6.99999999993145, 14.9999999999307, 3.99999999993179, 
    11.999999999931, 8.99999999993128, 16.9999999999305, 5.99999999993162, 
    2.99999999993187, 10.9999999999311, 7.99999999993145, 15.9999999999306, 
    4.9999999999317, 12.9999999999309, 9.99999999993119, 17.9999999999304, 
    6.99999999993145, 3.99999999993179, 11.999999999931, 8.99999999993128, 
    16.9999999999305, 5.99999999993162, 13.9999999999308, 2.99999999993187, 
    10.9999999999311, 18.9999999999303, 7.99999999993145, 4.9999999999317, 
    12.9999999999308, 9.99999999993119, 17.9999999999304, 6.99999999993145, 
    14.9999999999307, 3.99999999993179, 11.999999999931, 19.9999999999302, 
    8.99999999993128, 5.99999999993162, 13.9999999999308, 2.99999999993187, 
    10.9999999999311, 18.9999999999303, 7.99999999993145, 15.9999999999306, 
    4.9999999999317, 12.9999999999308, 20.9999999999301, 9.99999999993119, 
    6.99999999993145, 14.9999999999307, 3.99999999993179, 11.999999999931, 
    19.9999999999302, 8.99999999993127, 16.9999999999305, 5.99999999993162, 
    13.9999999999308, 21.99999999993, 2.99999999993187, 10.9999999999311, 
    7.99999999993145, 15.9999999999306, 4.9999999999317, 12.9999999999308, 
    20.9999999999301, 9.99999999993119, 17.9999999999304, 6.99999999993145, 
    14.9999999999307, 22.9999999999299, 3.99999999993179, 11.999999999931, 
    8.99999999993128, 16.9999999999305, 5.99999999993162, 13.9999999999308, 
    21.99999999993, 2.99999999993187, 10.9999999999311, 18.9999999999303, 
    7.99999999993145, 15.9999999999306, 23.9999999999298, 4.9999999999317, 
    12.9999999999308, 9.99999999993119, 17.9999999999304, 6.99999999993145, 
    14.9999999999307, 22.9999999999299, 3.99999999993179, 11.999999999931, 
    19.9999999999302, 8.99999999993127, 16.9999999999305, 24.9999999999297, 
    5.99999999993162, 13.9999999999308, 2.99999999993187, 10.9999999999311, 
    18.9999999999303, 7.99999999993145, 15.9999999999306, 23.9999999999298, 
    4.9999999999317, 12.9999999999308, 20.9999999999301, 9.99999999993119, 
    17.9999999999304, 25.9999999999296, 6.99999999993145, 14.9999999999307, 
    3.99999999993179, 11.999999999931, 19.9999999999302, 8.99999999993128, 
    16.9999999999305, 24.9999999999297, 5.99999999993162, 13.9999999999308, 
    21.99999999993, 2.99999999993187, 10.9999999999311, 18.9999999999303, 
    26.9999999999295, 7.99999999993145, 15.9999999999306, 4.9999999999317, 
    12.9999999999308, 20.9999999999301, 9.99999999993119, 17.9999999999304, 
    25.9999999999296, 6.99999999993145, 14.9999999999307, 22.9999999999299, 
    3.99999999993179, 11.999999999931, 19.9999999999302, 27.9999999999294, 
    8.99999999993128, 16.9999999999305, 5.99999999993162, 13.9999999999309, 
    21.99999999993, 2.99999999993187, 10.9999999999311, 18.9999999999303, 
    26.9999999999295, 7.99999999993145, 15.9999999999306, 23.9999999999298, 
    4.9999999999317, 12.9999999999308, 20.9999999999301, 28.9999999999293, 
    9.99999999993119, 17.9999999999304, 6.99999999993145, 14.9999999999307, 
    22.9999999999299, 3.99999999993179, 11.999999999931, 19.9999999999302, 
    27.9999999999294, 8.99999999993128, 16.9999999999305, 24.9999999999297, 
    5.99999999993162, 13.9999999999308, 21.99999999993, 2.99999999993187, 
    29.9999999999292, 10.9999999999311, 18.9999999999303, 7.99999999993145, 
    15.9999999999306, 23.9999999999298, 4.9999999999317, 12.9999999999308, 
    20.9999999999301, 28.9999999999293, 9.99999999993119, 17.9999999999304, 
    25.9999999999296, 6.99999999993145, 14.9999999999307, 22.9999999999299, 
    3.99999999993179, 30.9999999999291, 11.999999999931, 19.9999999999302, 
    8.99999999993128, 16.9999999999305, 24.9999999999297, 5.99999999993162, 
    13.9999999999308, 21.99999999993, 2.99999999993187, 29.9999999999292, 
    10.9999999999311, 18.9999999999303, 26.9999999999295, 7.99999999993145, 
    15.9999999999306, 23.9999999999298, 4.9999999999317, 31.999999999929, 
    12.9999999999308, 20.9999999999301, 9.99999999993119, 17.9999999999304, 
    25.9999999999296, 6.99999999993145, 14.9999999999307, 22.9999999999299, 
    3.99999999993179, 30.9999999999291, 11.999999999931, 19.9999999999302, 
    27.9999999999294, 8.99999999993128, 16.9999999999305, 24.9999999999297, 
    5.99999999993162, 32.9999999999289, 13.9999999999308, 21.99999999993, 
    2.99999999993187, 10.9999999999311, 18.9999999999303, 26.9999999999295, 
    7.99999999993145, 15.9999999999306, 23.9999999999298, 4.9999999999317, 
    31.999999999929, 12.9999999999309, 20.9999999999301, 28.9999999999293, 
    9.99999999993119, 17.9999999999304, 25.9999999999296, 6.99999999993145, 
    33.9999999999288, 14.9999999999307, 22.9999999999299, 3.99999999993179, 
    11.999999999931, 19.9999999999302, 27.9999999999294, 8.99999999993128, 
    16.9999999999305, 24.9999999999297, 5.99999999993162, 32.9999999999289, 
    13.9999999999308, 21.99999999993, 2.99999999993187, 29.9999999999292, 
    10.9999999999311, 18.9999999999303, 26.9999999999295, 7.99999999993145, 
    34.9999999999287, 15.9999999999306, 23.9999999999298, 4.9999999999317, 
    12.9999999999308, 20.9999999999301, 28.9999999999293, 9.99999999993119, 
    17.9999999999304, 25.9999999999296, 6.99999999993145, 33.9999999999288, 
    14.9999999999307, 22.9999999999299, 3.99999999993179, 30.9999999999291, 
    11.999999999931, 19.9999999999302, 27.9999999999294, 8.99999999993128, 
    35.9999999999286, 16.9999999999305, 24.9999999999297, 5.99999999993162, 
    13.9999999999308, 21.99999999993, 2.99999999993187, 29.9999999999292, 
    10.9999999999311, 18.9999999999303, 26.9999999999295, 7.99999999993145, 
    34.9999999999287, 15.9999999999306, 23.9999999999298, 4.9999999999317, 
    31.999999999929, 12.9999999999308, 20.9999999999301, 28.9999999999293, 
    9.99999999993119, 36.9999999999285, 17.9999999999304, 25.9999999999296, 
    6.99999999993145, 14.9999999999307, 22.9999999999299, 3.99999999993179, 
    30.9999999999291, 11.999999999931, 19.9999999999302, 27.9999999999294, 
    8.99999999993127, 35.9999999999286, 16.9999999999305, 24.9999999999297, 
    5.99999999993162, 32.9999999999289, 13.9999999999308, 21.99999999993, 
    2.99999999993187, 29.9999999999292, 10.9999999999311, 37.9999999999284, 
    18.9999999999303, 26.9999999999295, 7.99999999993145, 15.9999999999306, 
    23.9999999999298, 4.9999999999317, 31.999999999929, 12.9999999999308, 
    20.9999999999301, 28.9999999999293, 9.99999999993119, 36.9999999999285, 
    17.9999999999304, 25.9999999999296, 6.99999999993145, 33.9999999999288, 
    14.9999999999307, 22.9999999999299, 3.99999999993179, 30.9999999999291, 
    11.999999999931, 38.9999999999283, 19.9999999999302, 27.9999999999294, 
    8.99999999993128, 16.9999999999305, 24.9999999999297, 5.99999999993162, 
    32.9999999999289, 13.9999999999308, 21.99999999993, 2.99999999993187, 
    29.9999999999292, 10.9999999999311, 37.9999999999284, 18.9999999999303, 
    26.9999999999295, 7.99999999993145, 34.9999999999287, 15.9999999999306, 
    23.9999999999298, 4.9999999999317, 31.999999999929, 12.9999999999309, 
    39.9999999999283, 20.9999999999301, 28.9999999999293, 9.99999999993119, 
    17.9999999999304, 25.9999999999296, 6.99999999993145, 33.9999999999288, 
    14.9999999999307, 22.9999999999299, 3.99999999993179, 30.9999999999291, 
    11.999999999931, 38.9999999999283, 19.9999999999302, 27.9999999999294, 
    8.99999999993128, 35.9999999999286, 16.9999999999305, 24.9999999999297, 
    5.99999999993162, 32.9999999999289, 13.9999999999309, 40.9999999999281, 
    21.99999999993, 2.99999999993187, 29.9999999999292, 10.9999999999311, 
    18.9999999999303, 26.9999999999295, 7.99999999993145, 34.9999999999287, 
    15.9999999999306, 23.9999999999298, 4.9999999999317, 31.999999999929, 
    12.9999999999308, 39.9999999999282, 20.9999999999301, 28.9999999999293, 
    9.99999999993119, 36.9999999999285, 17.9999999999304, 25.9999999999296, 
    6.99999999993145, 33.9999999999288, 14.9999999999307, 41.999999999928, 
    22.9999999999299, 3.99999999993179, 30.9999999999291, 11.999999999931, 
    19.9999999999302, 27.9999999999294, 8.99999999993128, 35.9999999999286, 
    16.9999999999305, 24.9999999999297, 5.99999999993162, 32.9999999999289, 
    13.9999999999309, 40.9999999999281, 21.99999999993, 2.99999999993187, 
    29.9999999999292, 10.9999999999311, 37.9999999999284, 18.9999999999303, 
    26.9999999999295, 7.99999999993145, 34.9999999999287, 15.9999999999306, 
    42.9999999999279, 23.9999999999298, 4.9999999999317, 31.999999999929, 
    12.9999999999308, 20.9999999999301, 28.9999999999293, 9.99999999993119, 
    36.9999999999285, 17.9999999999304, 25.9999999999296, 6.99999999993145, 
    33.9999999999288, 14.9999999999307, 41.999999999928, 22.9999999999299, 
    3.99999999993179, 30.9999999999291, 11.999999999931, 38.9999999999283, 
    19.9999999999302, 27.9999999999294, 8.99999999993128, 35.9999999999286, 
    16.9999999999305, 43.9999999999278, 24.9999999999297, 5.99999999993162, 
    32.9999999999289, 13.9999999999308, 21.99999999993, 2.99999999993187, 
    29.9999999999292, 10.9999999999311, 37.9999999999284, 18.9999999999303, 
    26.9999999999295, 7.99999999993145, 34.9999999999287, 15.9999999999306, 
    42.9999999999279, 23.9999999999298, 4.9999999999317, 31.999999999929, 
    12.9999999999308, 39.9999999999282, 20.9999999999301, 28.9999999999293, 
    9.99999999993119, 36.9999999999285, 17.9999999999304, 44.9999999999277, 
    25.9999999999296, 6.99999999993145, 33.9999999999288, 14.9999999999307, 
    22.9999999999299, 3.99999999993179, 30.9999999999291, 11.999999999931, 
    38.9999999999283, 19.9999999999302, 27.9999999999294, 8.99999999993127, 
    35.9999999999286, 16.9999999999305, 43.9999999999278, 24.9999999999297, 
    5.99999999993162, 32.9999999999289, 13.9999999999308, 40.9999999999281, 
    21.99999999993, 2.99999999993187, 29.9999999999292, 10.9999999999311, 
    37.9999999999284, 18.9999999999303, 45.9999999999277, 26.9999999999295, 
    7.99999999993145, 34.9999999999287, 15.9999999999306, 23.9999999999298, 
    4.9999999999317, 31.999999999929, 12.9999999999308, 39.9999999999282, 
    20.9999999999301, 28.9999999999293, 9.99999999993119, 36.9999999999285, 
    17.9999999999304, 44.9999999999277, 25.9999999999296, 6.99999999993145, 
    33.9999999999288, 14.9999999999307, 41.999999999928, 22.9999999999299, 
    3.99999999993179, 30.9999999999291, 11.999999999931, 38.9999999999283, 
    19.9999999999302, 46.9999999999275, 27.9999999999294, 8.99999999993128, 
    35.9999999999286, 16.9999999999305, 24.9999999999297, 5.99999999993162, 
    32.9999999999289, 13.9999999999308, 40.9999999999281, 21.99999999993, 
    2.99999999993187, 29.9999999999292, 10.9999999999311, 37.9999999999284, 
    18.9999999999303, 45.9999999999277, 26.9999999999295, 7.99999999993145, 
    34.9999999999287, 15.9999999999306, 42.9999999999279, 23.9999999999298, 
    4.9999999999317, 31.999999999929, 12.9999999999308, 39.9999999999282, 
    20.9999999999301, 47.9999999999274, 28.9999999999293, 9.99999999993119, 
    36.9999999999285, 17.9999999999304, 25.9999999999296, 6.99999999993145, 
    33.9999999999288, 14.9999999999307, 41.999999999928, 22.9999999999299, 
    3.99999999993179, 30.9999999999291, 11.999999999931, 38.9999999999283, 
    19.9999999999302, 46.9999999999275, 27.9999999999294, 8.99999999993128, 
    35.9999999999286, 16.9999999999305, 43.9999999999278, 24.9999999999297, 
    5.99999999993162, 32.9999999999289, 13.9999999999308, 40.9999999999281, 
    21.99999999993, 2.99999999993187, 48.9999999999273, 29.9999999999292, 
    10.9999999999311, 37.9999999999284, 18.9999999999303, 26.9999999999295, 
    7.99999999993145, 34.9999999999287, 15.9999999999306, 42.9999999999279, 
    23.9999999999298, 4.9999999999317, 31.999999999929, 12.9999999999308, 
    39.9999999999282, 20.9999999999301, 47.9999999999274, 28.9999999999293, 
    9.99999999993119, 36.9999999999285, 17.9999999999304, 44.9999999999277, 
    25.9999999999296, 6.99999999993145, 33.9999999999288, 14.9999999999307, 
    41.999999999928, 22.9999999999299, 3.99999999993179, 49.9999999999273, 
    30.9999999999291, 11.999999999931, 38.9999999999283, 19.9999999999302, 
    27.9999999999294, 8.99999999993128, 35.9999999999286, 16.9999999999305, 
    43.9999999999278, 24.9999999999297, 5.99999999993162, 32.9999999999289, 
    13.9999999999308, 40.9999999999281, 21.99999999993, 2.99999999993187, 
    48.9999999999273, 29.9999999999292, 10.9999999999311, 37.9999999999284, 
    18.9999999999303, 45.9999999999277, 26.9999999999295, 7.99999999993145, 
    34.9999999999287, 15.9999999999306, 42.9999999999279, 23.9999999999298, 
    4.9999999999317, 50.9999999999271, 31.999999999929, 12.9999999999308, 
    39.9999999999282, 20.9999999999301, 28.9999999999293, 9.99999999993119, 
    36.9999999999285, 17.9999999999304, 44.9999999999277, 25.9999999999296, 
    6.99999999993145, 33.9999999999288, 14.9999999999307, 41.999999999928, 
    22.9999999999299, 3.99999999993179, 49.9999999999273, 30.9999999999291, 
    11.999999999931, 38.9999999999283, 19.9999999999302, 46.9999999999275, 
    27.9999999999294, 8.99999999993128, 35.9999999999286, 16.9999999999305, 
    43.9999999999278, 24.9999999999297, 5.99999999993162, 51.9999999999271, 
    32.9999999999289, 13.9999999999309, 40.9999999999281, 21.99999999993, 
    2.99999999993187, 29.9999999999292, 10.9999999999311, 37.9999999999284, 
    18.9999999999303, 45.9999999999277, 26.9999999999295, 7.99999999993145, 
    34.9999999999287, 15.9999999999306, 42.9999999999279, 23.9999999999298, 
    4.9999999999317, 50.9999999999271, 31.999999999929, 12.9999999999308, 
    39.9999999999282, 20.9999999999301, 47.9999999999274, 28.9999999999293, 
    9.99999999993119, 36.9999999999285, 17.9999999999304, 44.9999999999277, 
    25.9999999999296, 6.99999999993145, 33.9999999999288, 14.9999999999307, 
    41.999999999928, 22.9999999999299, 3.99999999993179, 30.9999999999291, 
    11.999999999931, 38.9999999999283, 19.9999999999302, 46.9999999999275, 
    27.9999999999294, 8.99999999993128, 35.9999999999286, 16.9999999999305, 
    43.9999999999278, 24.9999999999297, 5.99999999993162, 51.9999999999271, 
    32.9999999999289, 13.9999999999309, 40.9999999999281, 21.99999999993, 
    2.99999999993187, 48.9999999999273, 29.9999999999292, 10.9999999999311, 
    37.9999999999284, 18.9999999999303, 45.9999999999277, 26.9999999999295, 
    7.99999999993145, 34.9999999999287, 15.9999999999306, 42.9999999999279, 
    23.9999999999298, 4.9999999999317, 31.999999999929, 12.9999999999308, 
    39.9999999999282, 20.9999999999301, 47.9999999999274, 28.9999999999293, 
    9.99999999993119, 36.9999999999285, 17.9999999999304, 44.9999999999277, 
    25.9999999999296, 6.99999999993145, 33.9999999999288, 14.9999999999307, 
    41.999999999928, 22.9999999999299, 3.99999999993179, 49.9999999999273, 
    30.9999999999291, 11.999999999931, 38.9999999999283, 19.9999999999302, 
    46.9999999999275, 27.9999999999294, 8.99999999993128, 35.9999999999286, 
    16.9999999999305, 43.9999999999278, 24.9999999999297, 5.99999999993162, 
    32.9999999999289, 13.9999999999308, 40.9999999999281, 21.99999999993, 
    2.99999999993187, 48.9999999999273, 29.9999999999292, 10.9999999999311, 
    37.9999999999284, 18.9999999999303, 45.9999999999277, 26.9999999999295, 
    7.99999999993145, 34.9999999999287, 15.9999999999306, 42.9999999999279, 
    23.9999999999298, 4.9999999999317, 50.9999999999271, 31.999999999929, 
    12.9999999999308, 39.9999999999282, 20.9999999999301, 47.9999999999274, 
    28.9999999999293, 9.99999999993119, 36.9999999999285, 17.9999999999304, 
    44.9999999999277, 25.9999999999296, 6.99999999993145, 33.9999999999288, 
    14.9999999999307, 41.999999999928, 22.9999999999299, 3.99999999993179, 
    49.9999999999273, 30.9999999999291, 11.999999999931, 38.9999999999283, 
    19.9999999999302, 46.9999999999275, 27.9999999999294, 8.99999999993128, 
    35.9999999999286, 16.9999999999305, 43.9999999999278, 24.9999999999297, 
    5.99999999993162, 32.9999999999289, 13.9999999999308, 40.9999999999281, 
    21.99999999993, 2.99999999993187, 48.9999999999273, 29.9999999999292, 
    10.9999999999311, 37.9999999999284, 18.9999999999303, 45.9999999999277, 
    26.9999999999295, 7.99999999993145, 34.9999999999287, 15.9999999999306, 
    42.9999999999279, 23.9999999999298, 4.9999999999317, 31.999999999929, 
    12.9999999999308, 39.9999999999282, 20.9999999999301, 28.9999999999293, 
    9.99999999993119, 36.9999999999285, 17.9999999999304, 44.9999999999277, 
    25.9999999999296, 6.99999999993145, 33.9999999999288, 14.9999999999307, 
    41.999999999928, 22.9999999999299, 3.99999999993179, 49.9999999999273, 
    30.9999999999291, 11.999999999931, 38.9999999999283, 19.9999999999302, 
    46.9999999999275, 27.9999999999294, 8.99999999993128, 35.9999999999286, 
    16.9999999999305, 24.9999999999297, 5.99999999993162, 32.9999999999289, 
    13.9999999999308, 21.99999999993, 2.99999999993187, 29.9999999999292, 
    10.9999999999311, 37.9999999999284, 18.9999999999303, 45.9999999999276, 
    26.9999999999295, 7.99999999993145, 34.9999999999287, 15.9999999999306, 
    42.9999999999279, 23.9999999999298, 4.9999999999317, 31.999999999929, 
    12.9999999999309, 39.9999999999282, 20.9999999999301, 28.9999999999293, 
    9.99999999993119, 36.9999999999285, 17.9999999999304, 25.9999999999296, 
    6.99999999993145, 33.9999999999288, 14.9999999999307, 22.9999999999299, 
    3.99999999993179, 30.9999999999291, 11.999999999931, 38.9999999999283, 
    19.9999999999302, 46.9999999999275, 27.9999999999294, 8.99999999993128, 
    35.9999999999286, 16.9999999999305, 24.9999999999297, 5.99999999993162, 
    32.9999999999289, 13.9999999999309, 21.99999999993, 2.99999999993187, 
    29.9999999999292, 10.9999999999311, 37.9999999999284, 18.9999999999303, 
    26.9999999999295, 7.99999999993145, 34.9999999999287, 15.9999999999306, 
    23.9999999999298, 4.9999999999317, 31.999999999929, 12.9999999999308, 
    20.9999999999301, 28.9999999999293, 9.99999999993119, 36.9999999999285, 
    17.9999999999304, 25.9999999999296, 6.99999999993145, 33.9999999999288, 
    14.9999999999307, 22.9999999999299, 3.99999999993179, 30.9999999999291, 
    11.999999999931, 19.9999999999302, 27.9999999999294, 8.99999999993128, 
    35.9999999999286, 16.9999999999305, 24.9999999999297, 5.99999999993162, 
    32.9999999999289, 13.9999999999308, 21.99999999993, 2.99999999993187, 
    29.9999999999292, 10.9999999999311, 18.9999999999303, 26.9999999999295, 
    7.99999999993145, 34.9999999999287, 15.9999999999306, 23.9999999999298, 
    4.9999999999317, 31.999999999929, 12.9999999999308, 20.9999999999301, 
    28.9999999999293, 9.99999999993119, 17.9999999999304, 25.9999999999296, 
    6.99999999993145, 33.9999999999288, 14.9999999999307, 22.9999999999299, 
    3.99999999993179, 30.9999999999291, 11.999999999931, 19.9999999999302, 
    27.9999999999294, 8.99999999993128, 35.9999999999286, 16.9999999999305, 
    24.9999999999297, 5.99999999993162, 32.9999999999289, 13.9999999999309, 
    21.99999999993, 2.99999999993187, 29.9999999999292, 10.9999999999311, 
    18.9999999999303, 26.9999999999295, 7.99999999993145, 34.9999999999287, 
    15.9999999999306, 23.9999999999298, 4.9999999999317, 31.999999999929, 
    12.9999999999308, 20.9999999999301, 28.9999999999293, 9.99999999993119, 
    17.9999999999304, 25.9999999999296, 6.99999999993145, 33.9999999999288, 
    14.9999999999307, 22.9999999999299, 3.99999999993179, 30.9999999999291, 
    11.999999999931, 19.9999999999302, 27.9999999999294, 8.99999999993128, 
    16.9999999999305, 24.9999999999297, 5.99999999993162, 32.9999999999289, 
    13.9999999999308, 21.99999999993, 2.99999999993187, 29.9999999999292, 
    10.9999999999311, 18.9999999999303, 26.9999999999295, 7.99999999993145, 
    15.9999999999306, 23.9999999999298, 4.9999999999317, 31.999999999929, 
    12.9999999999308, 20.9999999999301, 28.9999999999293, 9.99999999993119, 
    17.9999999999304, 25.9999999999296, 6.99999999993145, 33.9999999999288, 
    14.9999999999307, 22.9999999999299, 3.99999999993179, 30.9999999999291, 
    11.999999999931, 19.9999999999302, 27.9999999999294, 8.99999999993128, 
    16.9999999999305, 24.9999999999297, 5.99999999993162, 13.9999999999308, 
    21.99999999993, 2.99999999993187, 29.9999999999292, 10.9999999999311, 
    18.9999999999303, 26.9999999999295, 7.99999999993145, 15.9999999999306, 
    23.9999999999298, 4.9999999999317, 12.9999999999308, 20.9999999999301, 
    28.9999999999293, 9.99999999993119, 17.9999999999304, 25.9999999999296, 
    6.99999999993145, 14.9999999999307, 22.9999999999299, 3.99999999993179, 
    30.9999999999291, 11.999999999931, 19.9999999999302, 27.9999999999294, 
    8.99999999993128, 16.9999999999305, 24.9999999999297, 5.99999999993162, 
    13.9999999999308, 21.99999999993, 2.99999999993187, 29.9999999999292, 
    10.9999999999311, 18.9999999999303, 26.9999999999295, 7.99999999993145, 
    15.9999999999306, 23.9999999999298, 4.9999999999317, 12.9999999999308, 
    20.9999999999301, 28.9999999999293, 9.99999999993119, 17.9999999999304, 
    25.9999999999296, 6.99999999993145, 14.9999999999307, 22.9999999999299, 
    3.99999999993179, 11.999999999931, 19.9999999999302, 27.9999999999294, 
    8.99999999993128, 16.9999999999305, 24.9999999999297, 5.99999999993162, 
    13.9999999999308, 21.99999999993, 2.99999999993187, 29.9999999999292, 
    10.9999999999311, 18.9999999999303, 26.9999999999295, 7.99999999993145, 
    15.9999999999306, 23.9999999999298, 4.9999999999317, 12.9999999999308, 
    20.9999999999301, 28.9999999999293, 9.99999999993119, 17.9999999999304, 
    25.9999999999296, 6.99999999993145, 14.9999999999307, 22.9999999999299, 
    3.99999999993179, 11.999999999931, 19.9999999999302, 27.9999999999294, 
    8.99999999993127, 16.9999999999305, 24.9999999999297, 5.99999999993162, 
    13.9999999999308, 21.99999999993, 2.99999999993187, 29.9999999999292, 
    10.9999999999311, 18.9999999999303, 26.9999999999295, 7.99999999993145, 
    15.9999999999306, 23.9999999999298, 4.9999999999317, 12.9999999999308, 
    20.9999999999301, 28.9999999999293, 9.99999999993119, 17.9999999999304, 
    25.9999999999296, 6.99999999993145, 14.9999999999307, 22.9999999999299, 
    3.99999999993179, 11.999999999931, 19.9999999999302, 27.9999999999294, 
    8.99999999993128, 16.9999999999305, 24.9999999999297, 5.99999999993162, 
    13.9999999999309, 21.99999999993, 2.99999999993187, 10.9999999999311, 
    18.9999999999303, 26.9999999999295, 7.99999999993145, 15.9999999999306, 
    23.9999999999298, 4.9999999999317, 12.9999999999308, 20.9999999999301, 
    9.99999999993119, 17.9999999999304, 25.9999999999296, 6.99999999993145, 
    14.9999999999307, 22.9999999999299, 3.99999999993179, 11.999999999931, 
    19.9999999999302, 27.9999999999294, 8.99999999993128, 16.9999999999305, 
    24.9999999999297, 5.99999999993162, 13.9999999999308, 21.99999999993, 
    2.99999999993187, 10.9999999999311, 18.9999999999303, 26.9999999999295, 
    7.99999999993145, 15.9999999999306, 23.9999999999298, 4.9999999999317, 
    12.9999999999308, 20.9999999999301, 28.9999999999293, 9.99999999993119, 
    17.9999999999304, 25.9999999999296, 6.99999999993145, 14.9999999999307, 
    22.9999999999299, 3.99999999993179, 11.999999999931, 19.9999999999302, 
    27.9999999999294, 8.99999999993128, 16.9999999999305, 24.9999999999297, 
    5.99999999993162, 13.9999999999308, 21.99999999993, 2.99999999993187, 
    10.9999999999311, 18.9999999999303, 26.9999999999295, 7.99999999993145, 
    15.9999999999306, 23.9999999999298, 4.9999999999317, 12.9999999999308, 
    20.9999999999301, 28.9999999999293, 9.99999999993119, 17.9999999999304, 
    25.9999999999296, 6.99999999993145, 14.9999999999307, 22.9999999999299, 
    3.99999999993179, 11.999999999931, 19.9999999999302, 8.99999999993128, 
    16.9999999999305, 24.9999999999297, 5.99999999993162, 13.9999999999308, 
    21.99999999993, 2.99999999993187, 10.9999999999311, 18.9999999999303, 
    26.9999999999295, 7.99999999993145, 15.9999999999306, 23.9999999999298, 
    4.9999999999317, 12.9999999999308, 20.9999999999301, 9.99999999993119, 
    17.9999999999304, 25.9999999999296, 6.99999999993145, 14.9999999999307, 
    22.9999999999299, 3.99999999993179, 11.999999999931, 19.9999999999302, 
    8.99999999993128, 16.9999999999305, 24.9999999999297, 5.99999999993162, 
    13.9999999999308, 21.99999999993, 2.99999999993187, 10.9999999999311, 
    18.9999999999303, 26.9999999999295, 7.99999999993145, 15.9999999999306, 
    23.9999999999298, 4.9999999999317, 12.9999999999308, 20.9999999999301, 
    9.99999999993119, 17.9999999999304, 25.9999999999296, 6.99999999993145, 
    14.9999999999307, 22.9999999999299, 3.99999999993179, 11.999999999931, 
    19.9999999999302, 8.99999999993128, 16.9999999999305, 24.9999999999297, 
    5.99999999993162, 13.9999999999308, 21.99999999993, 10.9999999999311, 
    18.9999999999303, 26.9999999999295, 7.99999999993145, 15.9999999999306, 
    23.9999999999298, 4.9999999999317, 12.9999999999308, 20.9999999999301, 
    9.99999999993119, 17.9999999999304, 25.9999999999296, 6.99999999993145, 
    14.9999999999307, 22.9999999999299, 11.999999999931, 19.9999999999302, 
    27.9999999999294, 8.99999999993127, 16.9999999999305, 24.9999999999297, 
    5.99999999993162, 13.9999999999309, 21.99999999993, 10.9999999999311, 
    18.9999999999303, 26.9999999999295, 7.99999999993145, 15.9999999999306, 
    23.9999999999298, 12.9999999999308, 20.9999999999301, 9.99999999993119, 
    17.9999999999304, 25.9999999999296, 6.99999999993145, 14.9999999999307, 
    22.9999999999299, 11.999999999931, 19.9999999999302, 27.9999999999294, 
    8.99999999993128, 16.9999999999305, 24.9999999999297, 13.9999999999308, 
    21.99999999993, 10.9999999999311, 18.9999999999303, 26.9999999999295, 
    7.99999999993145, 15.9999999999306, 23.9999999999298, 12.9999999999309, 
    20.9999999999301, 9.99999999993119, 17.9999999999304, 25.9999999999296, 
    14.9999999999307, 22.9999999999299, 11.999999999931, 19.9999999999302, 
    27.9999999999294, 8.99999999993128, 16.9999999999305, 24.9999999999297, 
    13.9999999999308, 21.99999999993, 10.9999999999311, 18.9999999999303, 
    26.9999999999295, 15.9999999999306, 23.9999999999298, 12.9999999999308, 
    20.9999999999301, 9.99999999993119, 17.9999999999304, 25.9999999999296, 
    14.9999999999307, 22.9999999999299, 11.999999999931, 19.9999999999302, 
    27.9999999999294, 16.9999999999305, 24.9999999999297, 13.9999999999309, 
    21.99999999993, 10.9999999999311, 18.9999999999303, 26.9999999999295, 
    15.9999999999306, 23.9999999999298, 12.9999999999309, 20.9999999999301, 
    17.9999999999304, 25.9999999999296, 14.9999999999307, 22.9999999999299, 
    11.999999999931, 19.9999999999302, 27.9999999999294, 16.9999999999305, 
    24.9999999999297, 13.9999999999308, 21.99999999993, 18.9999999999303, 
    26.9999999999295, 15.9999999999306, 23.9999999999298, 12.9999999999308, 
    20.9999999999301, 28.9999999999293, 17.9999999999304, 25.9999999999296, 
    14.9999999999307, 22.9999999999299, 19.9999999999302, 27.9999999999294, 
    16.9999999999305, 24.9999999999297, 13.9999999999308, 21.99999999993, 
    18.9999999999303, 26.9999999999295, 15.9999999999306, 23.9999999999298, 
    20.9999999999301, 28.9999999999293, 17.9999999999304, 25.9999999999296, 
    14.9999999999307, 22.9999999999299, 19.9999999999302, 27.9999999999294, 
    16.9999999999305, 24.9999999999297, 21.99999999993, 18.9999999999303, 
    26.9999999999295, 15.9999999999306, 23.9999999999298, 20.9999999999301, 
    28.9999999999293, 17.9999999999304, 25.9999999999296, 22.9999999999299, 
    19.9999999999302, 27.9999999999294, 16.9999999999305, 24.9999999999297, 
    21.99999999993, 18.9999999999303, 26.9999999999295, 23.9999999999298, 
    20.9999999999301, 28.9999999999293, 17.9999999999304, 25.9999999999296, 
    22.9999999999299, 19.9999999999302, 27.9999999999294, 24.9999999999297, 
    21.99999999993, 18.9999999999303, 26.9999999999295, 23.9999999999298, 
    20.9999999999301, 28.9999999999293, 25.9999999999296, 22.9999999999299, 
    19.9999999999302, 27.9999999999294, 24.9999999999297, 21.99999999993, 
    26.9999999999295, 23.9999999999298, 20.9999999999301, 28.9999999999293, 
    25.9999999999296, 22.9999999999299, 27.9999999999294, 24.9999999999297, 
    21.99999999993, 29.9999999999292, 26.9999999999295, 23.9999999999298, 
    28.9999999999293, 25.9999999999296, 22.9999999999299, 27.9999999999294, 
    24.9999999999297, 29.9999999999292, 26.9999999999295, 23.9999999999298, 
    28.9999999999293, 25.9999999999296, 27.9999999999294, 24.9999999999297, 
    29.9999999999292, 26.9999999999295, 28.9999999999293, 25.9999999999296, 
    27.9999999999294, 26.9999999999295, 28.9999999999293, 27.9999999999294, 
    29.9999999999292, 28.9999999999293 ;

 obs_Ygrid = 2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36.0272723111239, 36.9000015258789, 38.0571408952985, 
    38.7000045776367, 39.9857155936105, 41.0999977111816, 41.8875017166138, 
    42.9000015258789, 44.0999984741211, 45.042856488909, 45.9000015258789, 
    47.0699981689453, 48, 48.9000018726696, 50.1272714788263, 51, 
    51.9000015258789, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0727258162065, 36, 
    36.9000015258789, 38.0999977111816, 38.9142870221819, 39.9000011444092, 
    41.1999969482422, 42.0999984741211, 42.8625011444092, 45.2999954223633, 
    45.9000026157924, 47.0999977111816, 48, 48.9000015258789, 
    50.0999994277954, 51, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.8000011444092, 38.1428555079869, 38.7750034332275, 40.1000022888183, 
    40.9499988555908, 42.0999984741211, 42.75, 43.7999954223633, 
    45.0599990844727, 46.0000038146972, 47.0999984741211, 48, 
    48.9000015258789, 50.1374988555908, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.1666653951009, 33, 34.020002746582, 35.0727258162065, 
    35.9333343505859, 36.9857155936105, 38.1857136317662, 38.7000045776367, 
    40.9499988555908, 41.9250011444092, 45.0999984741211, 45.9000027974446, 
    47.0999984741211, 48, 48.9000015258789, 50.0999984741211, 51, 
    51.9000015258789, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 32.2799995422363, 33, 
    33.9272741837935, 35.0142844063895, 35.9142870221819, 40.9499988555908, 
    42, 45.1124982833862, 45.9272741837935, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 50.9727276888761, 51.8625011444092, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 45.960001373291, 47.0999984741211, 
    48, 50.0999984741211, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0727258162065, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.1299983978271, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 
    20.9727276888761, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.8625011444092, 20.1374988555908, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 17.9625005722046, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    16.979997253418, 2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 
    11.8500022888184, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 11.8500022888184, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.86250114440917, 10.9499988555908, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.86250114440917, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.05714089529856, 8.94000091552734, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 2.10000038146972, 
    3, 3.89999961853028, 5.10000038146972, 23.7539978027344, 
    23.7539978027344, 23.7539978027344, 23.7539978027344, 23.7539978027344, 
    23.7539978027344, 23.7539978027344, 23.7539978027344, 23.7539978027344, 
    23.7539978027344, 23.7539978027344, 23.7539978027344, 23.7539978027344, 
    23.7539978027344, 23.7539978027344, 23.7539978027344, 23.7539978027344, 
    23.7539978027344, 23.7539978027344, 23.7539978027344, 23.7539978027344, 
    23.7539978027344, 23.7539978027344, 23.7539978027344, 23.7539978027344, 
    23.7539978027344, 23.7539978027344, 23.7539978027344, 23.7539978027344, 
    23.7539978027344, 23.7539978027344, 23.7539978027344, 23.7539978027344, 
    23.7539978027344, 23.7539978027344, 23.7539978027344, 23.7539978027344, 
    23.7539978027344, 26.3579978942871, 26.3579978942871, 26.3579978942871, 
    26.3579978942871, 26.3579978942871, 26.3579978942871, 26.3579978942871, 
    26.3579978942871, 26.3579978942871, 26.3579978942871, 26.3579978942871, 
    26.3579978942871, 26.3579978942871, 26.3579978942871, 26.3579978942871, 
    26.3579978942871, 26.3579978942871, 26.3579978942871, 26.3579978942871, 
    26.3579978942871, 26.3579978942871, 26.3579978942871, 26.3579978942871, 
    26.3579978942871, 26.3579978942871, 26.3579978942871, 26.3579978942871, 
    26.3579978942871, 26.3579978942871, 26.3579978942871, 26.3579978942871, 
    26.3579978942871, 26.3579978942871, 26.3579978942871, 26.3579978942871, 
    26.3579978942871, 26.3579978942871, 26.3579978942871, 26.3579978942871, 
    26.3579978942871, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36.0272723111239, 36.9000015258789, 38.0571408952985, 
    38.7000045776367, 39.9000005722046, 41.0999977111816, 41.8875017166138, 
    42.9000015258789, 44.0999984741211, 45.042856488909, 45.9000015258789, 
    47.0699981689453, 48, 48.9000018726696, 50.1599990844726, 51, 
    51.9000015258789, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0727258162065, 36, 
    36.9000015258789, 38.0999977111816, 38.9142870221819, 39.9000011444092, 
    41.1999969482422, 42.0999984741211, 42.8625011444092, 45.2999954223633, 
    45.9000026157924, 47.0999977111816, 48, 48.9000015258789, 
    50.2000007629394, 51, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000022888184, 35.0999984741211, 36, 
    36.8000011444092, 38.1428555079869, 38.7750034332275, 40.1000022888183, 
    40.9499988555908, 42.0999984741211, 42.75, 43.7999954223633, 
    45.0599990844727, 46.0000038146972, 47.0999984741211, 48, 
    48.9000015258789, 50.1374988555908, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.1666653951009, 33, 34.020002746582, 35.0727258162065, 
    35.9333343505859, 36.9857155936105, 38.1857136317662, 38.7000045776367, 
    40.9499988555908, 41.9250011444092, 45.0999984741211, 45.9000027974446, 
    47.0999984741211, 48, 48.9000015258789, 50.0999984741211, 51, 
    51.9000015258789, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 32.2799995422363, 
    33.0374994277954, 33.9272741837935, 35.0142844063895, 35.9142870221819, 
    40.9499988555908, 42, 45.1124982833862, 45.9272741837935, 
    47.0999984741211, 48, 48.9000015258789, 50.0999984741211, 
    50.9727276888761, 51.8625011444092, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 
    45.960001373291, 47.0999984741211, 48, 50.0999984741211, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0727258162065, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.1299983978271, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 
    20.9727276888761, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.8625011444092, 20.1374988555908, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 17.9625005722046, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    16.979997253418, 2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 
    11.8500022888184, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 11.8500022888184, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.86250114440917, 10.9499988555908, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.86250114440917, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.05714089529856, 8.94000091552734, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 2.10000038146972, 
    3, 3.89999961853028, 5.10000038146972, 13.3680038452148, 
    13.3680038452148, 13.3680038452148, 13.3680038452148, 13.3680038452148, 
    13.3680038452148, 13.3680038452148, 13.3680038452148, 13.3680038452148, 
    13.3680038452148, 13.3680038452148, 13.3680038452148, 13.3680038452148, 
    13.3680038452148, 13.3680038452148, 13.3680038452148, 13.3680038452148, 
    13.3680038452148, 13.3680038452148, 13.3680038452148, 13.3680038452148, 
    13.3680038452148, 13.3680038452148, 13.3680038452148, 13.3680038452148, 
    13.3680038452148, 13.3680038452148, 13.3680038452148, 13.3680038452148, 
    13.3680038452148, 13.3680038452148, 13.3680038452148, 13.3680038452148, 
    13.3680038452148, 13.3680038452148, 13.3680038452148, 13.3680038452148, 
    13.3680038452148, 13.3680038452148, 13.3680038452148, 13.3680038452148, 
    13.3680038452148, 13.3680038452148, 13.3680038452148, 13.3680038452148, 
    13.3680038452148, 37.7250022888184, 37.7250022888184, 37.7250022888184, 
    37.7250022888184, 37.7250022888184, 37.7250022888184, 37.7250022888184, 
    37.7250022888184, 37.7250022888184, 37.7250022888184, 37.7250022888184, 
    37.7250022888184, 37.7250022888184, 37.7250022888184, 37.7250022888184, 
    37.7250022888184, 37.7250022888184, 37.7250022888184, 37.7250022888184, 
    37.7250022888184, 37.7250022888184, 37.7250022888184, 37.7250022888184, 
    37.7250022888184, 37.7250022888184, 37.7250022888184, 37.7250022888184, 
    37.7250022888184, 37.7250022888184, 37.7250022888184, 37.7250022888184, 
    37.7250022888184, 37.7250022888184, 37.7250022888184, 37.7250022888184, 
    37.7250022888184, 37.7250022888184, 37.7250022888184, 37.7250022888184, 
    37.7250022888184, 37.7250022888184, 37.7250022888184, 37.7250022888184, 
    37.7250022888184, 37.7250022888184, 37.7250022888184, 45.6870002746582, 
    45.6870002746582, 45.6870002746582, 45.6870002746582, 45.6870002746582, 
    45.6870002746582, 45.6870002746582, 45.6870002746582, 45.6870002746582, 
    45.6870002746582, 45.6870002746582, 45.6870002746582, 45.6870002746582, 
    45.6870002746582, 45.6870002746582, 45.6870002746582, 2.10000038146972, 
    3, 3.89999961853028, 5.10000038146972, 5.99999809265136, 
    6.90000152587891, 8.09999847412109, 9, 9.90000152587891, 
    11.0999984741211, 12, 12.9000015258789, 14.0999984741211, 15, 
    15.9000015258789, 17.0999984741211, 18, 18.9000015258789, 
    20.0999984741211, 21, 21.9000015258789, 23.0999984741211, 24, 
    24.9000015258789, 26.0999984741211, 27, 27.9000015258789, 
    29.0999984741211, 30, 30.9000015258789, 32.0999984741211, 33, 
    33.9000015258789, 35.0999984741211, 36, 36.9000015258789, 
    38.0999984741211, 39, 39.9000015258789, 41.0999984741211, 42, 
    42.9000015258789, 44.0999984741211, 45, 45.9000015258789, 
    47.0999984741211, 48, 48.9000015258789, 50.0999984741211, 51, 
    51.9000015258789, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 
    36.0666656494141, 36.9000015258789, 37.874997138977, 39.9000005722046, 
    40.7999954223633, 41.8285740443638, 42.9000015258789, 44.0999984741211, 
    45.042856488909, 45.9000022888184, 47.0999981273304, 48, 
    48.9000018726696, 50.1599990844726, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0727258162065, 
    36.033332824707, 36.9000015258789, 38.0999977111816, 38.9500007629395, 
    39.9000011444092, 40.7999954223633, 41.8500022888184, 42.8625011444092, 
    45.2999954223633, 45.9000034332275, 47.0999977111816, 48, 
    48.9000015258789, 50.2000007629394, 51, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.8250017166138, 
    35.0999965667724, 36.0999984741211, 36.7000007629395, 38.1428555079869, 
    38.7750034332275, 40.1000022888183, 41.1000022888183, 42.0599990844727, 
    42.75, 43.7999954223633, 45.2999954223633, 46.0000038146972, 
    47.0999984741211, 48, 48.9000015258789, 50.0999984741211, 51, 
    51.9000015258789, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.8727285211736, 
    32.1666653951009, 32.9700004577637, 33.6000022888184, 35.0399963378906, 
    35.7000045776367, 38.1750011444092, 38.7000045776367, 40.9499988555908, 
    42.1499977111816, 45.1499977111816, 45.9000027974446, 47.0999984741211, 
    48, 48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 32.2799995422363, 
    33.0374994277954, 33.9000015258789, 36, 42.1499977111816, 
    45.1124982833862, 45.9272741837935, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 50.9727276888761, 51.8625011444092, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 45.960001373291, 47.0999984741211, 
    48, 50.0999984741211, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0727258162065, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.1299983978271, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 
    20.9727276888761, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.8625011444092, 20.1374988555908, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 17.9625005722046, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    16.979997253418, 2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 
    11.8500022888184, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 11.8500022888184, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.86250114440917, 10.9499988555908, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.86250114440917, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.05714089529856, 8.94000091552734, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 2.10000038146972, 
    3, 3.89999961853028, 5.10000038146972, 34.7880020141601, 
    34.7880020141601, 34.7880020141601, 34.7880020141601, 34.7880020141601, 
    34.7880020141601, 34.7880020141601, 34.7880020141601, 34.7880020141601, 
    34.7880020141601, 34.7880020141601, 34.7880020141601, 34.7880020141601, 
    33.6509971618652, 33.6509971618652, 33.6509971618652, 33.6509971618652, 
    33.6509971618652, 33.6509971618652, 33.6509971618652, 33.6509971618652, 
    33.6509971618652, 33.6509971618652, 33.6509971618652, 33.6509971618652, 
    33.6509971618652, 33.6509971618652, 8.8440055847168, 8.8440055847168, 
    8.8440055847168, 8.8440055847168, 8.8440055847168, 8.8440055847168, 
    8.8440055847168, 8.8440055847168, 8.8440055847168, 8.8440055847168, 
    8.8440055847168, 8.8440055847168, 8.8440055847168, 8.8440055847168, 
    8.7509994506836, 8.7509994506836, 8.7509994506836, 8.7509994506836, 
    8.7509994506836, 8.7509994506836, 8.7509994506836, 8.7509994506836, 
    8.7509994506836, 8.7509994506836, 8.7509994506836, 8.7509994506836, 
    8.7509994506836, 8.7509994506836, 8.7509994506836, 8.7509994506836, 
    8.7509994506836, 8.7509994506836, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 30, 
    30.9000015258789, 32.0999984741211, 33, 33.9000015258789, 
    35.0999984741211, 36, 36.9000015258789, 38.0999984741211, 39, 
    39.9000015258789, 41.0999984741211, 42, 42.9000015258789, 
    44.0999984741211, 45, 45.9000015258789, 47.0999984741211, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 30, 30.9000015258789, 
    32.0999984741211, 33, 33.9000015258789, 35.0999984741211, 36, 
    36.9000015258789, 38.0999984741211, 39, 39.9000015258789, 
    41.0999984741211, 42, 42.9000015258789, 44.0999984741211, 45, 
    45.9000015258789, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999981273304, 30, 
    30.8727285211736, 32.0999984741211, 33, 33.9000015258789, 
    35.0727258162065, 36.042856488909, 36.8625011444092, 38.1000022888183, 
    42.9000015258789, 44.0999988555908, 45.0374994277954, 45.8666687011719, 
    47.0999981273304, 48, 48.9000015258789, 50.0999984741211, 51, 
    51.9000015258789, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999981273304, 30, 30.9000015258789, 
    32.0999981273304, 32.8800018310547, 34.0285737173898, 34.9874982833862, 
    36.0999984741211, 36.8000005086263, 37.9499988555908, 44.1750011444092, 
    45.1499977111816, 45.7500028610229, 47.1299983978271, 48, 
    48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.8625011444092, 29.0624985694885, 30, 30.8571444920131, 
    31.979997253418, 34.7999954223633, 36.2999954223633, 45.1499977111816, 
    46.0000019073486, 47.0999984741211, 48, 48.9000015258789, 
    50.0999984741211, 51, 51.8625011444092, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0727258162065, 
    29.9727276888761, 32.2124991416931, 32.9700004577637, 33.6000022888184, 
    38.7000045776367, 45.1499977111816, 45.9000022888184, 47.0999984741211, 
    48, 48.9000015258789, 50.0999984741211, 51, 51.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0999984741211, 27, 
    27.9000015258789, 29.0999984741211, 29.9142870221819, 32.2799995422363, 
    33, 33.6000022888184, 45.1124982833862, 45.9272741837935, 
    47.0999984741211, 48, 48.9000015258789, 50.0999984741211, 
    50.9727276888761, 51.8625011444092, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 24, 24.9000015258789, 
    26.0999984741211, 27, 27.9000015258789, 29.0999984741211, 
    45.960001373291, 47.0999984741211, 48, 50.0999984741211, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 26.0727258162065, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.9000015258789, 20.0999984741211, 21, 21.9000015258789, 
    23.0999984741211, 24, 24.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 21, 
    21.9000015258789, 23.0999984741211, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 18, 18.9000015258789, 20.0999984741211, 
    20.9727276888761, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 17.0999984741211, 18, 
    18.8625011444092, 20.1374988555908, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    17.0999984741211, 17.9625005722046, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 15.9000015258789, 
    16.979997253418, 2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    14.0999984741211, 15, 15.9000015258789, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 14.0999984741211, 15, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 12, 
    12.9000015258789, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 12.9000015258789, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.90000152587891, 11.0999984741211, 12, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 11.0999984741211, 
    11.8500022888184, 2.10000038146972, 3, 3.89999961853028, 
    5.10000038146972, 5.99999809265136, 6.90000152587891, 8.09999847412109, 
    9, 9.90000152587891, 11.0999984741211, 11.8500022888184, 
    2.10000038146972, 3, 3.89999961853028, 5.10000038146972, 
    5.99999809265136, 6.90000152587891, 8.09999847412109, 9, 
    9.86250114440917, 10.9499988555908, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.90000152587891, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.09999847412109, 9, 9.86250114440917, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 6.90000152587891, 
    8.05714089529856, 8.94000091552734, 2.10000038146972, 3, 
    3.89999961853028, 5.10000038146972, 5.99999809265136, 2.10000038146972, 
    3, 3.89999961853028, 5.10000038146972, 8.04899597167969, 
    8.04899597167969, 8.04899597167969, 8.04899597167969, 8.04899597167969, 
    8.04899597167969, 8.04899597167969, 8.04899597167969, 8.04899597167969, 
    8.04899597167969, 8.04899597167969, 8.04899597167969, 8.04899597167969, 
    8.04899597167969, 8.04899597167969, 8.04899597167969, 8.04899597167969, 
    8.04899597167969, 7.04100036621093, 7.04100036621093, 7.04100036621093, 
    7.04100036621093, 7.04100036621093, 7.04100036621093, 7.04100036621093, 
    7.04100036621093, 7.04100036621093, 7.04100036621093, 7.04100036621093, 
    7.04100036621093, 7.04100036621093, 7.04100036621093, 7.04100036621093, 
    7.04100036621093, 7.04100036621093, 7.04100036621093, 7.04100036621093, 
    7.04100036621093, 7.04100036621093, 7.04100036621093, 7.04100036621093, 
    7.04100036621093, 7.04100036621093, 7.04100036621093, 7.04100036621093, 
    7.04100036621093, 7.04100036621093, 7.04100036621093, 2.8511893712683, 
    2.8511893712683, 3.70751696511747, 2.8511893712683, 3.70751696511747, 
    2.8511893712683, 3.70751696511747, 2.8511893712683, 3.70751696511747, 
    6.26097000315193, 2.8511893712683, 3.70751696511747, 6.26097000315193, 
    2.8511893712683, 7.10690132310917, 3.70751696511747, 6.26097000315193, 
    2.8511893712683, 7.10690132310917, 3.70751696511747, 6.26097000315193, 
    7.95020197539848, 2.8511893712683, 7.10690132310917, 3.70751696511747, 
    6.26097000315193, 7.95020197539848, 2.8511893712683, 7.10690132310917, 
    8.79085990591997, 3.70751696511747, 6.26097000315193, 7.95020197539848, 
    2.8511893712683, 7.10690132310917, 8.79085990591997, 3.70751696511747, 
    6.26097000315193, 7.95020197539848, 2.8511893712683, 9.62886335158985, 
    7.10690132310916, 8.79085990591997, 3.70751696511747, 6.26097000315193, 
    7.95020197539848, 2.8511893712683, 9.62886335158985, 7.10690132310917, 
    8.79085990591997, 3.70751696511747, 11.296861184434, 6.26097000315193, 
    7.95020197539848, 2.8511893712683, 9.62886335158985, 7.10690132310917, 
    8.79085990591997, 3.70751696511747, 11.296861184434, 6.26097000315193, 
    7.95020197539848, 2.8511893712683, 9.62886335158985, 12.126833490299, 
    7.10690132310916, 8.79085990591997, 3.70751696511747, 11.296861184434, 
    6.26097000315193, 7.95020197539848, 2.8511893712683, 9.62886335158985, 
    12.126833490299, 7.10690132310917, 8.79085990591997, 3.70751696511747, 
    11.296861184434, 6.26097000315193, 12.9541071462105, 7.95020197539848, 
    2.8511893712683, 9.62886335158985, 12.126833490299, 7.10690132310916, 
    8.79085990591997, 3.70751696511747, 11.296861184434, 6.26097000315193, 
    12.9541071462105, 7.95020197539848, 2.8511893712683, 9.62886335158985, 
    12.126833490299, 7.10690132310916, 13.7786718264961, 8.79085990591997, 
    3.70751696511747, 11.296861184434, 6.26097000315193, 12.9541071462105, 
    7.95020197539848, 2.8511893712683, 9.62886335158985, 12.126833490299, 
    7.10690132310917, 13.7786718264961, 8.79085990591997, 3.70751696511747, 
    11.296861184434, 6.26097000315193, 12.9541071462105, 7.95020197539848, 
    2.8511893712683, 14.60051748906, 9.62886335158985, 12.126833490299, 
    7.10690132310916, 13.7786718264961, 8.79085990591997, 3.70751696511747, 
    11.296861184434, 6.26097000315193, 12.9541071462105, 7.95020197539848, 
    2.8511893712683, 14.60051748906, 9.62886335158985, 12.126833490299, 
    7.10690132310916, 13.7786718264961, 8.79085990591997, 3.70751696511747, 
    16.2360130019538, 11.296861184434, 6.26097000315193, 12.9541071462105, 
    7.95020197539848, 2.8511893712683, 14.60051748906, 9.62886335158985, 
    12.126833490299, 7.10690132310917, 13.7786718264961, 8.79085990591997, 
    3.70751696511747, 16.2360130019538, 11.296861184434, 6.26097000315193, 
    12.9541071462105, 7.95020197539848, 2.8511893712683, 14.60051748906, 
    9.62886335158985, 17.0496441729557, 12.126833490299, 7.10690132310917, 
    13.7786718264961, 8.79085990591997, 3.70751696511747, 16.2360130019538, 
    11.296861184434, 6.26097000315193, 12.9541071462105, 7.95020197539848, 
    2.8511893712683, 14.60051748906, 9.62886335158985, 17.0496441729557, 
    12.126833490299, 7.10690132310917, 13.7786718264961, 8.79085990591997, 
    3.70751696511747, 16.2360130019538, 11.296861184434, 6.26097000315193, 
    17.860518964504, 12.9541071462105, 7.95020197539848, 2.8511893712683, 
    14.60051748906, 9.62886335158985, 17.0496441729557, 12.126833490299, 
    7.10690132310916, 13.7786718264961, 8.79085990591997, 3.70751696511747, 
    16.2360130019538, 11.296861184434, 6.26097000315193, 17.860518964504, 
    12.9541071462105, 7.95020197539848, 2.8511893712683, 14.60051748906, 
    9.62886335158985, 17.0496441729557, 12.126833490299, 7.10690132310916, 
    18.6686287301423, 13.7786718264961, 8.79085990591997, 3.70751696511747, 
    16.2360130019538, 11.296861184434, 6.26097000315193, 17.860518964504, 
    12.9541071462105, 7.95020197539848, 2.8511893712683, 14.60051748906, 
    9.62886335158985, 17.0496441729557, 12.126833490299, 7.10690132310917, 
    18.6686287301423, 13.7786718264961, 8.79085990591997, 3.70751696511747, 
    16.2360130019538, 11.296861184434, 6.26097000315193, 17.860518964504, 
    12.9541071462105, 7.95020197539848, 20.2765199679718, 2.8511893712683, 
    14.60051748906, 9.62886335158985, 17.0496441729557, 12.126833490299, 
    7.10690132310916, 18.6686287301423, 13.7786718264961, 8.79085990591997, 
    3.70751696511747, 16.2360130019538, 11.296861184434, 6.26097000315193, 
    17.860518964504, 12.9541071462105, 7.95020197539848, 20.2765199679718, 
    2.8511893712683, 14.60051748906, 9.62886335158985, 17.0496441729557, 
    12.126833490299, 7.10690132310917, 18.6686287301423, 13.7786718264961, 
    8.79085990591997, 21.0762855122492, 3.70751696511747, 16.2360130019538, 
    11.296861184434, 6.26097000315193, 17.860518964504, 12.9541071462105, 
    7.95020197539848, 20.2765199679718, 2.8511893712683, 14.60051748906, 
    9.62886335158985, 17.0496441729557, 12.126833490299, 7.10690132310917, 
    18.6686287301423, 13.7786718264961, 8.79085990591997, 21.0762855122492, 
    3.70751696511747, 16.2360130019538, 11.296861184434, 6.26097000315193, 
    17.860518964504, 12.9541071462105, 7.95020197539848, 20.2765199679718, 
    2.8511893712683, 14.60051748906, 9.62886335158985, 21.8732541712884, 
    17.0496441729557, 12.126833490299, 7.10690132310916, 18.6686287301423, 
    13.7786718264961, 8.79085990591997, 21.0762855122492, 3.70751696511747, 
    16.2360130019538, 11.296861184434, 6.26097000315193, 17.860518964504, 
    12.9541071462105, 7.95020197539848, 20.2765199679718, 2.8511893712683, 
    14.60051748906, 9.62886335158985, 21.8732541712884, 17.0496441729557, 
    12.126833490299, 7.10690132310917, 18.6686287301423, 13.7786718264961, 
    8.79085990591997, 21.0762855122492, 3.70751696511747, 16.2360130019538, 
    11.296861184434, 22.6674186531335, 6.26097000315193, 17.860518964504, 
    12.9541071462105, 7.95020197539848, 20.2765199679718, 2.8511893712683, 
    14.60051748906, 9.62886335158985, 21.8732541712884, 17.0496441729557, 
    12.126833490299, 7.10690132310917, 18.6686287301423, 13.7786718264961, 
    8.79085990591997, 21.0762855122492, 3.70751696511747, 16.2360130019538, 
    11.296861184434, 22.6674186531335, 6.26097000315193, 17.860518964504, 
    12.9541071462105, 7.95020197539848, 20.2765199679718, 2.8511893712683, 
    14.60051748906, 9.62886335158985, 21.8732541712884, 17.0496441729557, 
    12.126833490299, 24.2473072431218, 7.10690132310916, 18.6686287301423, 
    13.7786718264961, 8.79085990591997, 21.0762855122492, 3.70751696511747, 
    16.2360130019538, 11.296861184434, 22.6674186531335, 6.26097000315193, 
    17.860518964504, 12.9541071462105, 7.95020197539848, 20.2765199679718, 
    2.8511893712683, 14.60051748906, 9.62886335158985, 21.8732541712884, 
    17.0496441729557, 12.126833490299, 24.2473072431218, 7.10690132310916, 
    18.6686287301423, 13.7786718264961, 8.79085990591997, 21.0762855122492, 
    3.70751696511747, 16.2360130019538, 11.296861184434, 22.6674186531335, 
    6.26097000315193, 17.860518964504, 12.9541071462105, 25.0330180873813, 
    7.95020197539848, 20.2765199679718, 2.8511893712683, 14.60051748906, 
    9.62886335158985, 21.8732541712884, 17.0496441729557, 12.126833490299, 
    24.2473072431218, 7.10690132310917, 18.6686287301423, 13.7786718264961, 
    8.79085990591997, 21.0762855122492, 3.70751696511747, 16.2360130019538, 
    11.296861184434, 22.6674186531335, 6.26097000315193, 17.860518964504, 
    12.9541071462105, 25.0330180873813, 7.95020197539848, 20.2765199679718, 
    2.8511893712683, 14.60051748906, 9.62886335158985, 21.8732541712884, 
    17.0496441729557, 12.126833490299, 24.2473072431218, 7.10690132310916, 
    18.6686287301423, 13.7786718264961, 25.8158982228162, 8.79085990591997, 
    21.0762855122492, 3.70751696511747, 16.2360130019538, 11.296861184434, 
    22.6674186531335, 6.26097000315193, 17.860518964504, 12.9541071462105, 
    25.0330180873813, 7.95020197539848, 20.2765199679718, 2.8511893712683, 
    14.60051748906, 9.62886335158985, 21.8732541712884, 17.0496441729557, 
    12.126833490299, 24.2473072431218, 7.10690132310916, 18.6686287301423, 
    13.7786718264961, 25.8158982228162, 8.79085990591997, 21.0762855122492, 
    3.70751696511747, 16.2360130019538, 11.296861184434, 22.6674186531335, 
    6.26097000315193, 17.860518964504, 12.9541071462105, 25.0330180873813, 
    7.95020197539848, 20.2765199679718, 2.8511893712683, 14.60051748906, 
    26.9845421774241, 9.62886335158985, 21.8732541712884, 17.0496441729557, 
    12.126833490299, 24.2473072431218, 7.10690132310916, 18.6686287301423, 
    13.7786718264961, 25.8158982228162, 8.79085990591997, 21.0762855122492, 
    3.70751696511747, 16.2360130019538, 11.296861184434, 22.6674186531335, 
    6.26097000315193, 17.860518964504, 12.9541071462105, 25.0330180873813, 
    7.95020197539848, 20.2765199679718, 2.8511893712683, 14.60051748906, 
    26.9845421774241, 9.62886335158985, 21.8732541712884, 17.0496441729557, 
    12.126833490299, 24.2473072431218, 7.10690132310916, 18.6686287301423, 
    13.7786718264961, 25.8158982228162, 8.79085990591997, 21.0762855122492, 
    3.70751696511747, 16.2360130019538, 28.147495817899, 11.296861184434, 
    22.6674186531335, 6.26097000315193, 17.860518964504, 12.9541071462105, 
    25.0330180873813, 7.95020197539848, 20.2765199679718, 2.8511893712683, 
    14.60051748906, 26.9845421774241, 9.62886335158985, 21.8732541712884, 
    17.0496441729557, 12.126833490299, 24.2473072431218, 7.10690132310916, 
    18.6686287301423, 13.7786718264961, 25.8158982228162, 8.79085990591997, 
    21.0762855122492, 3.70751696511747, 16.2360130019538, 28.147495817899, 
    11.296861184434, 22.6674186531335, 6.26097000315193, 17.860518964504, 
    12.9541071462105, 25.0330180873813, 7.95020197539848, 20.2765199679718, 
    2.8511893712683, 14.60051748906, 26.9845421774241, 9.62886335158985, 
    21.8732541712884, 17.0496441729557, 28.9189958304827, 12.126833490299, 
    24.2473072431218, 7.10690132310916, 18.6686287301423, 13.7786718264961, 
    25.8158982228162, 8.79085990591997, 21.0762855122492, 3.70751696511747, 
    16.2360130019538, 28.147495817899, 11.296861184434, 22.6674186531335, 
    6.26097000315193, 17.860518964504, 12.9541071462105, 25.0330180873813, 
    7.95020197539848, 20.2765199679718, 2.8511893712683, 14.60051748906, 
    26.9845421774241, 9.62886335158985, 21.8732541712884, 17.0496441729557, 
    28.9189958304827, 12.126833490299, 24.2473072431218, 7.10690132310917, 
    18.6686287301423, 13.7786718264961, 25.8158982228162, 8.79085990591997, 
    21.0762855122492, 3.70751696511747, 16.2360130019538, 28.147495817899, 
    11.296861184434, 22.6674186531335, 6.26097000315193, 17.860518964504, 
    29.6876377539464, 12.9541071462105, 25.0330180873813, 7.95020197539848, 
    20.2765199679718, 2.8511893712683, 14.60051748906, 26.9845421774241, 
    9.62886335158985, 21.8732541712884, 17.0496441729557, 28.9189958304827, 
    12.126833490299, 24.2473072431218, 7.10690132310916, 18.6686287301423, 
    13.7786718264961, 25.8158982228162, 8.79085990591997, 21.0762855122492, 
    3.70751696511747, 16.2360130019538, 28.147495817899, 11.296861184434, 
    22.6674186531335, 6.26097000315193, 17.860518964504, 29.6876377539464, 
    12.9541071462105, 25.0330180873813, 7.95020197539848, 20.2765199679718, 
    2.8511893712683, 14.60051748906, 26.9845421774241, 9.62886335158985, 
    21.8732541712884, 17.0496441729557, 28.9189958304827, 12.126833490299, 
    24.2473072431218, 7.10690132310916, 18.6686287301423, 31.2163286776756, 
    13.7786718264961, 25.8158982228162, 8.79085990591997, 21.0762855122492, 
    3.70751696511747, 16.2360130019538, 28.147495817899, 11.296861184434, 
    22.6674186531335, 6.26097000315193, 17.860518964504, 29.6876377539464, 
    12.9541071462105, 25.0330180873813, 7.95020197539848, 20.2765199679718, 
    2.8511893712683, 14.60051748906, 26.9845421774241, 9.62886335158985, 
    21.8732541712884, 17.0496441729557, 28.9189958304827, 12.126833490299, 
    24.2473072431218, 7.10690132310917, 18.6686287301423, 31.2163286776756, 
    13.7786718264961, 25.8158982228162, 8.79085990591997, 21.0762855122492, 
    3.70751696511747, 16.2360130019538, 28.147495817899, 11.296861184434, 
    22.6674186531335, 6.26097000315193, 17.860518964504, 29.6876377539464, 
    12.9541071462105, 25.0330180873813, 7.95020197539848, 20.2765199679718, 
    31.9763689611184, 2.8511893712683, 14.60051748906, 26.9845421774241, 
    9.62886335158985, 21.8732541712884, 17.0496441729557, 28.9189958304827, 
    12.126833490299, 24.2473072431218, 7.10690132310916, 18.6686287301423, 
    31.2163286776756, 13.7786718264961, 25.8158982228162, 8.79085990591997, 
    21.0762855122492, 3.70751696511747, 16.2360130019538, 28.147495817899, 
    11.296861184434, 22.6674186531335, 6.26097000315193, 17.860518964504, 
    29.6876377539464, 12.9541071462105, 25.0330180873813, 7.95020197539848, 
    20.2765199679718, 31.9763689611184, 2.8511893712683, 14.60051748906, 
    26.9845421774241, 9.62886335158985, 21.8732541712884, 17.0496441729557, 
    28.9189958304827, 12.126833490299, 24.2473072431218, 7.10690132310916, 
    18.6686287301423, 31.2163286776756, 13.7786718264961, 25.8158982228162, 
    8.79085990591997, 21.0762855122492, 32.7335337174312, 3.70751696511747, 
    16.2360130019538, 28.147495817899, 11.296861184434, 22.6674186531335, 
    6.26097000315193, 17.860518964504, 29.6876377539464, 12.9541071462105, 
    25.0330180873813, 7.95020197539848, 20.2765199679718, 31.9763689611184, 
    2.8511893712683, 14.60051748906, 26.9845421774241, 9.62886335158985, 
    21.8732541712884, 17.0496441729557, 28.9189958304827, 12.126833490299, 
    24.2473072431218, 7.10690132310916, 18.6686287301423, 31.2163286776756, 
    13.7786718264961, 25.8158982228162, 8.79085990591997, 21.0762855122492, 
    32.7335337174312, 3.70751696511747, 16.2360130019538, 28.147495817899, 
    11.296861184434, 22.6674186531335, 6.26097000315193, 17.860518964504, 
    29.6876377539464, 12.9541071462105, 25.0330180873813, 7.95020197539848, 
    20.2765199679718, 31.9763689611184, 2.8511893712683, 14.60051748906, 
    26.9845421774241, 9.62886335158985, 21.8732541712884, 34.2392218564619, 
    17.0496441729557, 28.9189958304827, 12.126833490299, 24.2473072431218, 
    7.10690132310916, 18.6686287301423, 31.2163286776756, 13.7786718264961, 
    25.8158982228162, 8.79085990591997, 21.0762855122492, 32.7335337174312, 
    3.70751696511747, 16.2360130019538, 28.147495817899, 11.296861184434, 
    22.6674186531335, 6.26097000315193, 17.860518964504, 29.6876377539464, 
    12.9541071462105, 25.0330180873813, 7.95020197539848, 20.2765199679718, 
    31.9763689611184, 14.60051748906, 26.9845421774241, 9.62886335158985, 
    21.8732541712884, 34.2392218564619, 17.0496441729557, 28.9189958304827, 
    12.126833490299, 24.2473072431218, 7.10690132310917, 18.6686287301423, 
    31.2163286776756, 13.7786718264961, 25.8158982228162, 8.79085990591997, 
    21.0762855122492, 32.7335337174312, 3.70751696511747, 16.2360130019538, 
    28.147495817899, 11.296861184434, 22.6674186531335, 34.9877384320501, 
    6.26097000315193, 17.860518964504, 29.6876377539464, 12.9541071462105, 
    25.0330180873813, 7.95020197539848, 20.2765199679718, 31.9763689611184, 
    14.60051748906, 26.9845421774241, 9.62886335158985, 21.8732541712884, 
    34.2392218564619, 17.0496441729557, 28.9189958304827, 12.126833490299, 
    24.2473072431218, 7.10690132310917, 18.6686287301423, 31.2163286776756, 
    13.7786718264961, 25.8158982228162, 8.79085990591997, 21.0762855122492, 
    32.7335337174312, 16.2360130019538, 28.147495817899, 11.296861184434, 
    22.6674186531335, 34.9877384320501, 6.26097000315193, 17.860518964504, 
    29.6876377539464, 12.9541071462105, 25.0330180873813, 7.95020197539848, 
    20.2765199679718, 31.9763689611184, 14.60051748906, 26.9845421774241, 
    9.62886335158985, 21.8732541712884, 34.2392218564619, 17.0496441729557, 
    28.9189958304827, 12.126833490299, 24.2473072431218, 35.7333658617202, 
    7.10690132310916, 18.6686287301423, 31.2163286776756, 13.7786718264961, 
    25.8158982228162, 8.79085990591997, 21.0762855122492, 32.7335337174312, 
    16.2360130019538, 28.147495817899, 11.296861184434, 22.6674186531335, 
    34.9877384320501, 6.26097000315193, 17.860518964504, 29.6876377539464, 
    12.9541071462105, 25.0330180873813, 7.95020197539848, 20.2765199679718, 
    31.9763689611184, 14.60051748906, 26.9845421774241, 9.62886335158985, 
    21.8732541712884, 34.2392218564619, 17.0496441729557, 28.9189958304827, 
    12.126833490299, 24.2473072431218, 35.7333658617202, 7.10690132310917, 
    18.6686287301423, 31.2163286776756, 13.7786718264961, 25.8158982228162, 
    8.79085990591997, 21.0762855122492, 32.7335337174312, 16.2360130019538, 
    28.147495817899, 11.296861184434, 22.6674186531335, 34.9877384320501, 
    17.860518964504, 29.6876377539464, 12.9541071462105, 25.0330180873813, 
    37.2159422114215, 7.95020197539848, 20.2765199679718, 31.9763689611184, 
    14.60051748906, 26.9845421774241, 9.62886335158985, 21.8732541712884, 
    34.2392218564619, 17.0496441729557, 28.9189958304827, 12.126833490299, 
    24.2473072431218, 35.7333658617202, 18.6686287301423, 31.2163286776756, 
    13.7786718264961, 25.8158982228162, 21.0762855122492, 32.7335337174312, 
    16.2360130019538, 28.147495817899, 11.296861184434, 22.6674186531335, 
    34.9877384320501, 17.860518964504, 29.6876377539464, 12.9541071462105, 
    25.0330180873813, 37.2159422114215, 7.95020197539848, 20.2765199679718, 
    31.9763689611184, 14.60051748906, 26.9845421774241, 9.62886335158985, 
    21.8732541712884, 34.2392218564619, 17.0496441729557, 28.9189958304827, 
    24.2473072431218, 35.7333658617202, 18.6686287301423, 31.2163286776756, 
    25.8158982228162, 37.9528861616004, 21.0762855122492, 32.7335337174312, 
    16.2360130019538, 28.147495817899, 11.296861184434, 22.6674186531335, 
    34.9877384320501, 17.860518964504, 29.6876377539464, 12.9541071462105, 
    25.0330180873813, 37.2159422114215, 20.2765199679718, 31.9763689611184, 
    14.60051748906, 26.9845421774241, 21.8732541712884, 34.2392218564619, 
    17.0496441729557, 28.9189958304827, 24.2473072431218, 35.7333658617202, 
    18.6686287301423, 31.2163286776756, 25.8158982228162, 37.9528861616004, 
    21.0762855122492, 32.7335337174312, 16.2360130019538, 28.147495817899, 
    11.296861184434, 22.6674186531335, 34.9877384320501, 17.860518964504, 
    29.6876377539464, 25.0330180873813, 37.2159422114215, 20.2765199679718, 
    31.9763689611184, 26.9845421774241, 38.6869310214985, 21.8732541712884, 
    34.2392218564619, 17.0496441729557, 28.9189958304827, 24.2473072431218, 
    35.7333658617202, 18.6686287301423, 31.2163286776756, 25.8158982228162, 
    37.9528861616004, 21.0762855122492, 32.7335337174312, 28.147495817899, 
    22.6674186531335, 34.9877384320501, 17.860518964504, 29.6876377539464, 
    25.0330180873813, 37.2159422114215, 20.2765199679718, 31.9763689611184, 
    26.9845421774241, 38.6869310214985, 21.8732541712884, 34.2392218564619, 
    28.9189958304827, 24.2473072431218, 35.7333658617202, 18.6686287301423, 
    31.2163286776756, 25.8158982228162, 37.9528861616004, 21.0762855122492, 
    32.7335337174312, 28.147495817899, 40.146315971085, 22.6674186531335, 
    34.9877384320501, 29.6876377539464, 25.0330180873813, 37.2159422114215, 
    20.2765199679718, 31.9763689611184, 26.9845421774241, 38.6869310214985, 
    21.8732541712884, 34.2392218564619, 28.9189958304827, 24.2473072431218, 
    35.7333658617202, 31.2163286776756, 25.8158982228162, 37.9528861616004, 
    21.0762855122492, 32.7335337174312, 28.147495817899, 40.146315971085, 
    22.6674186531335, 34.9877384320501, 29.6876377539464, 25.0330180873813, 
    37.2159422114215, 20.2765199679718, 31.9763689611184, 26.9845421774241, 
    38.6869310214985, 21.8732541712884, 34.2392218564619, 28.9189958304827, 
    40.8716528537064, 24.2473072431218, 35.7333658617202, 31.2163286776756, 
    25.8158982228162, 37.9528861616004, 21.0762855122492, 32.7335337174312, 
    28.147495817899, 40.146315971085, 22.6674186531335, 34.9877384320501, 
    29.6876377539464, 25.0330180873813, 37.2159422114215, 31.9763689611184, 
    26.9845421774241, 38.6869310214985, 21.8732541712884, 34.2392218564619, 
    28.9189958304827, 40.8716528537064, 24.2473072431218, 35.7333658617202, 
    31.2163286776756, 25.8158982228162, 37.9528861616004, 32.7335337174312, 
    28.147495817899, 40.146315971085, 22.6674186531335, 34.9877384320501, 
    29.6876377539464, 42.313609019804, 25.0330180873813, 37.2159422114215, 
    31.9763689611184, 26.9845421774241, 38.6869310214985, 34.2392218564619, 
    28.9189958304827, 40.8716528537064, 24.2473072431218, 35.7333658617202, 
    31.2163286776756, 25.8158982228162, 37.9528861616004, 32.7335337174312, 
    28.147495817899, 40.146315971085, 22.6674186531335, 34.9877384320501, 
    29.6876377539464, 42.313609019804, 25.0330180873813, 37.2159422114215, 
    31.9763689611184, 26.9845421774241, 38.6869310214985, 34.2392218564619, 
    28.9189958304827, 40.8716528537064, 35.7333658617202, 31.2163286776756, 
    43.0302263684599, 25.8158982228162, 37.9528861616004, 32.7335337174312, 
    28.147495817899, 40.146315971085, 34.9877384320501, 29.6876377539464, 
    42.313609019804, 37.2159422114215, 31.9763689611184, 26.9845421774241, 
    38.6869310214985, 34.2392218564619, 28.9189958304827, 40.8716528537064, 
    35.7333658617202, 31.2163286776756, 43.0302263684599, 25.8158982228162, 
    37.9528861616004, 32.7335337174312, 28.147495817899, 40.146315971085, 
    34.9877384320501, 29.6876377539464, 42.313609019804, 37.2159422114215, 
    31.9763689611184, 43.743935615978, 26.9845421774241, 38.6869310214985, 
    34.2392218564619, 28.9189958304827, 40.8716528537064, 35.7333658617202, 
    31.2163286776756, 43.0302263684599, 37.9528861616004, 32.7335337174312, 
    28.147495817899, 40.146315971085, 34.9877384320501, 29.6876377539464, 
    42.313609019804, 37.2159422114215, 31.9763689611184, 43.7439356159779, 
    38.6869310214985, 34.2392218564619, 28.9189958304827, 40.8716528537064, 
    35.7333658617202, 31.2163286776756, 43.0302263684599, 37.9528861616004, 
    32.7335337174312, 45.1626281947156, 28.147495817899, 40.146315971085, 
    34.9877384320501, 29.6876377539464, 42.313609019804, 37.2159422114215, 
    31.9763689611184, 43.7439356159779, 38.6869310214985, 34.2392218564619, 
    28.9189958304827, 40.8716528537064, 35.7333658617202, 31.2163286776756, 
    43.0302263684599, 37.9528861616004, 32.7335337174312, 45.1626281947156, 
    40.146315971085, 34.9877384320501, 29.6876377539464, 42.313609019804, 
    37.2159422114215, 31.9763689611184, 43.7439356159779, 38.6869310214985, 
    34.2392218564619, 45.8676112200792, 28.9189958304827, 40.8716528537064, 
    35.7333658617202, 31.2163286776756, 43.0302263684599, 37.9528861616004, 
    32.7335337174312, 45.1626281947156, 40.146315971085, 34.9877384320501, 
    29.6876377539464, 42.313609019804, 37.2159422114215, 31.9763689611184, 
    43.7439356159779, 38.6869310214985, 34.2392218564619, 45.8676112200792, 
    40.8716528537064, 35.7333658617202, 31.2163286776756, 43.0302263684599, 
    37.9528861616004, 32.7335337174312, 45.1626281947156, 40.146315971085, 
    34.9877384320501, 47.268851454425, 42.313609019804, 37.2159422114215, 
    31.9763689611184, 43.7439356159779, 38.6869310214985, 34.2392218564619, 
    45.8676112200792, 40.8716528537064, 35.7333658617202, 43.0302263684599, 
    37.9528861616004, 32.7335337174312, 45.1626281947156, 40.146315971085, 
    34.9877384320501, 47.268851454425, 42.313609019804, 37.2159422114215, 
    31.9763689611184, 43.7439356159779, 38.6869310214985, 34.2392218564619, 
    45.8676112200792, 40.8716528537064, 35.7333658617202, 47.965109528352, 
    43.0302263684599, 37.9528861616004, 32.7335337174312, 45.1626281947156, 
    40.146315971085, 34.9877384320501, 47.268851454425, 42.313609019804, 
    37.2159422114215, 31.9763689611184, 43.7439356159779, 38.6869310214985, 
    34.2392218564619, 45.8676112200792, 40.8716528537064, 35.7333658617202, 
    47.965109528352, 43.0302263684599, 37.9528861616004, 32.7335337174312, 
    45.1626281947156, 40.146315971085, 34.9877384320501, 47.268851454425, 
    42.313609019804, 37.2159422114215, 49.0036828201845, 43.7439356159779, 
    38.6869310214985, 34.2392218564619, 45.8676112200792, 40.8716528537064, 
    35.7333658617202, 47.965109528352, 43.0302263684599, 37.9528861616004, 
    32.7335337174312, 45.1626281947156, 40.146315971085, 34.9877384320501, 
    47.268851454425, 42.313609019804, 37.2159422114215, 49.0036828201845, 
    43.7439356159779, 38.6869310214985, 45.8676112200792, 40.8716528537064, 
    35.7333658617202, 47.965109528352, 43.0302263684599, 37.9528861616004, 
    50.0364447368152, 45.1626281947156, 40.146315971085, 34.9877384320501, 
    47.268851454425, 42.313609019804, 37.2159422114215, 49.0036828201845, 
    43.7439356159779, 38.6869310214985, 45.8676112200792, 40.8716528537064, 
    35.7333658617202, 47.965109528352, 43.0302263684599, 37.9528861616004, 
    50.0364447368153, 45.1626281947156, 40.146315971085, 47.268851454425, 
    42.313609019804, 37.2159422114215, 49.0036828201845, 43.7439356159779, 
    38.6869310214985, 51.0619470586162, 45.8676112200792, 40.8716528537064, 
    35.7333658617202, 47.965109528352, 43.0302263684599, 37.9528861616004, 
    50.0364447368152, 45.1626281947156, 40.146315971085, 47.268851454425, 
    42.313609019804, 37.2159422114215, 49.0036828201845, 43.7439356159779, 
    38.6869310214985, 51.0619470586162, 45.8676112200792, 40.8716528537064, 
    47.965109528352, 43.0302263684599, 37.9528861616004, 50.0364447368153, 
    45.1626281947156, 40.146315971085, 47.268851454425, 42.313609019804, 
    37.2159422114215, 49.0036828201845, 43.7439356159779, 38.6869310214985, 
    51.0619470586162, 45.8676112200792, 40.8716528537064, 47.965109528352, 
    43.0302263684599, 37.9528861616004, 50.0364447368152, 45.1626281947156, 
    40.146315971085, 47.268851454425, 42.313609019804, 37.2159422114215, 
    49.0036828201845, 43.743935615978, 38.6869310214985, 51.0619470586162, 
    45.8676112200792, 40.8716528537064, 47.965109528352, 43.0302263684599, 
    37.9528861616004, 50.0364447368152, 45.1626281947156, 40.146315971085, 
    47.268851454425, 42.313609019804, 49.0036828201845, 43.7439356159779, 
    38.6869310214985, 51.0619470586162, 45.8676112200792, 40.8716528537064, 
    47.965109528352, 43.0302263684599, 37.9528861616004, 50.0364447368152, 
    45.1626281947156, 40.1463159710849, 47.268851454425, 42.313609019804, 
    49.0036828201845, 43.7439356159779, 38.6869310214985, 51.0619470586162, 
    45.8676112200792, 40.8716528537064, 47.965109528352, 43.0302263684599, 
    50.0364447368152, 45.1626281947156, 40.146315971085, 47.268851454425, 
    42.313609019804, 49.0036828201845, 43.743935615978, 38.6869310214985, 
    51.0619470586162, 45.8676112200792, 40.8716528537064, 47.965109528352, 
    43.0302263684599, 50.0364447368152, 45.1626281947156, 40.1463159710849, 
    47.268851454425, 42.313609019804, 49.0036828201845, 43.743935615978, 
    51.0619470586162, 45.8676112200792, 40.8716528537064, 47.965109528352, 
    43.0302263684599, 50.0364447368153, 45.1626281947156, 40.146315971085, 
    47.268851454425, 42.313609019804, 49.0036828201845, 43.7439356159779, 
    51.0619470586162, 45.8676112200792, 40.8716528537064, 47.965109528352, 
    43.0302263684599, 50.0364447368153, 45.1626281947156, 47.268851454425, 
    42.313609019804, 49.0036828201845, 43.7439356159779, 51.0619470586162, 
    45.8676112200792, 40.8716528537064, 47.965109528352, 43.0302263684599, 
    50.0364447368152, 45.1626281947156, 47.268851454425, 42.313609019804, 
    49.0036828201845, 43.7439356159779, 51.0619470586162, 45.8676112200792, 
    40.8716528537064, 47.965109528352, 43.0302263684599, 50.0364447368152, 
    45.1626281947156, 47.268851454425, 42.313609019804, 49.0036828201845, 
    43.7439356159779, 51.0619470586162, 45.8676112200792, 47.965109528352, 
    43.0302263684599, 50.0364447368153, 45.1626281947156, 47.268851454425, 
    42.313609019804, 49.0036828201845, 43.7439356159779, 51.0619470586162, 
    45.8676112200792, 47.965109528352, 43.0302263684599, 50.0364447368152, 
    45.1626281947156, 47.268851454425, 49.0036828201845, 43.7439356159779, 
    51.0619470586162, 45.8676112200792, 47.965109528352, 43.0302263684599, 
    50.0364447368152, 45.1626281947156, 47.268851454425, 49.0036828201845, 
    43.743935615978, 51.0619470586162, 45.8676112200792, 47.965109528352, 
    50.0364447368152, 45.1626281947156, 47.268851454425, 49.0036828201845, 
    43.7439356159779, 51.0619470586162, 45.8676112200792, 47.965109528352, 
    50.0364447368153, 45.1626281947156, 47.268851454425, 49.0036828201845, 
    51.0619470586162, 45.8676112200792, 47.965109528352, 50.0364447368152, 
    45.1626281947156, 47.268851454425, 49.0036828201845, 51.0619470586162, 
    45.8676112200792, 47.965109528352, 50.0364447368152, 47.268851454425, 
    49.0036828201845, 51.0619470586162, 45.8676112200792, 47.965109528352, 
    50.0364447368152, 47.268851454425, 49.0036828201845, 51.0619470586162, 
    45.8676112200792, 47.965109528352, 50.0364447368153, 47.268851454425, 
    49.0036828201845, 51.0619470586162, 47.965109528352, 50.0364447368152, 
    47.268851454425, 49.0036828201845, 51.0619470586162, 47.965109528352, 
    50.0364447368152, 49.0036828201845, 51.0619470586162, 47.965109528352, 
    50.0364447368152, 49.0036828201845, 51.0619470586162, 50.0364447368153, 
    51.0619470586162, 50.0364447368152, 51.0619470586162, 50.0364447368152, 
    51.0619470586162 ;

 obs_Zgrid = 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0 ;

 obs_lon = -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -125.983334859212, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.987879897609, -125.983334859212, 
    -125.947621663411, -125.833333333333, -125.961906069801, 
    -125.953334554036, -125.945834477743, -125.983334859212, 
    -126.083333333333, -126.047619047619, -125.983334859212, 
    -126.003334554036, -125.983334859212, -125.987879897609, 
    -125.987879897609, -125.996971361565, -125.983334859212, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.678786769058, -125.683331807454, -125.683331807454, 
    -125.71333211263, -125.647618611654, -125.673331197103, 
    -125.799997965495, -125.749997456868, -125.745831807454, 
    -125.683331807454, -125.733331589472, -125.66333211263, 
    -125.683331807454, -125.683331807454, -125.808331807454, 
    -125.653331502279, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.366668701172, -125.333333333333, -125.333333333333, 
    -125.350001017253, -125.3047601609, -125.358334859212, -125.40000406901, 
    -125.233327229818, -125.316665649414, -125.433339436849, 
    -125.283330281576, -125.31333211263, -125.299997965495, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.320832570394, -125.333333333333, -125.333333333333, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.988889906141, -124.983334859212, -124.933333333333, 
    -124.996971361565, -124.988889906142, -124.961906069801, 
    -125.047621227446, -125.133336385091, -125.083333333333, 
    -124.933335622152, -125.000001695421, -124.966668023003, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.683331807454, 
    -124.683331807454, -124.683331807454, -124.683331807454, 
    -124.683331807454, -124.683331807454, -124.683331807454, 
    -124.683331807454, -124.683331807454, -124.683331807454, 
    -124.683331807454, -124.683331807454, -124.753331502279, 
    -124.733332316081, -124.696968309807, -124.733331589472, 
    -124.747618175688, -124.633336385091, -124.799997965495, 
    -124.708331425985, -124.696968309807, -124.683331807454, 
    -124.683331807454, -124.683331807454, -124.683331807454, 
    -124.696968309807, -124.745831807454, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.37333577474, -124.383336385091, -124.383336385091, 
    -124.433339436849, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -123.983334859212, -123.983334859212, -123.983334859212, 
    -123.983334859212, -123.983334859212, -123.983334859212, 
    -123.983334859212, -123.996971361565, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.683331807454, -123.683331807454, 
    -123.683331807454, -123.683331807454, -123.683331807454, 
    -123.683331807454, -123.683331807454, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -122.983334859212, 
    -122.983334859212, -122.983334859212, -122.983334859212, 
    -123.013335164388, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.683331807454, -122.683331807454, -122.696968309807, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.345834096273, 
    -122.345834096273, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.045834859212, 
    -121.633331298828, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.633331298828, -121.633331298828, 
    -121.673329671224, -121.333333333333, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.333333333333, 
    -121.333333333333, -121.033335367839, -121.033335367839, 
    -121.033335367839, -121.033335367839, -121.033335367839, 
    -121.033335367839, -121.033335367839, -121.033335367839, 
    -121.033335367839, -121.033335367839, -121.033335367839, 
    -121.033335367839, -121.083333333333, -121.083333333333, 
    -120.633331298828, -120.633331298828, -120.633331298828, 
    -120.633331298828, -120.633331298828, -120.633331298828, 
    -120.633331298828, -120.633331298828, -120.633331298828, 
    -120.633331298828, -120.645831425985, -120.633331298828, 
    -120.333333333333, -120.333333333333, -120.333333333333, 
    -120.333333333333, -120.333333333333, -120.333333333333, 
    -120.333333333333, -120.333333333333, -120.333333333333, 
    -120.333333333333, -120.320832570394, -120.333333333333, 
    -120.033335367839, -120.033335367839, -120.033335367839, 
    -120.033335367839, -120.033335367839, -120.033335367839, 
    -120.033335367839, -120.033335367839, -120.033335367839, 
    -120.033335367839, -120.033335367839, -120.033335367839, 
    -119.633331298828, -119.633331298828, -119.633331298828, 
    -119.633331298828, -119.633331298828, -119.633331298828, 
    -119.633331298828, -119.633331298828, -119.633331298828, 
    -119.633331298828, -119.633331298828, -119.333333333333, 
    -119.333333333333, -119.333333333333, -119.333333333333, 
    -119.333333333333, -119.333333333333, -119.333333333333, 
    -119.333333333333, -119.333333333333, -119.333333333333, 
    -119.333333333333, -119.033335367839, -119.033335367839, 
    -119.033335367839, -119.033335367839, -119.033335367839, 
    -119.033335367839, -119.033335367839, -119.033335367839, 
    -119.033335367839, -119.033335367839, -119.033335367839, 
    -118.633331298828, -118.633331298828, -118.633331298828, 
    -118.633331298828, -118.633331298828, -118.633331298828, 
    -118.633331298828, -118.633331298828, -118.620831807454, 
    -118.633331298828, -118.333333333333, -118.333333333333, 
    -118.333333333333, -118.333333333333, -118.333333333333, 
    -118.333333333333, -118.333333333333, -118.333333333333, 
    -118.333333333333, -118.033335367839, -118.033335367839, 
    -118.033335367839, -118.033335367839, -118.033335367839, 
    -118.033335367839, -118.033335367839, -118.033335367839, 
    -118.045834859212, -117.633331298828, -117.633331298828, 
    -117.633331298828, -117.633331298828, -117.633331298828, 
    -117.633331298828, -117.661903018043, -117.693330891927, 
    -117.333333333333, -117.333333333333, -117.333333333333, 
    -117.333333333333, -117.333333333333, -117.033335367839, 
    -117.033335367839, -117.033335367839, -117.083333333333, 
    -128.625340779622, -128.625340779622, -128.625340779622, 
    -128.625340779622, -128.625340779622, -128.625340779622, 
    -128.625340779622, -128.625340779622, -128.625340779622, 
    -128.625340779622, -128.625340779622, -128.625340779622, 
    -128.625340779622, -128.625340779622, -128.625340779622, 
    -128.625340779622, -128.625340779622, -128.625340779622, 
    -128.625340779622, -128.625340779622, -128.625340779622, 
    -128.625340779622, -128.625340779622, -128.625340779622, 
    -128.625340779622, -128.625340779622, -128.625340779622, 
    -128.625340779622, -128.625340779622, -128.625340779622, 
    -128.625340779622, -128.625340779622, -128.625340779622, 
    -128.625340779622, -128.625340779622, -128.625340779622, 
    -128.625340779622, -128.625340779622, -127.52333577474, -127.52333577474, 
    -127.52333577474, -127.52333577474, -127.52333577474, -127.52333577474, 
    -127.52333577474, -127.52333577474, -127.52333577474, -127.52333577474, 
    -127.52333577474, -127.52333577474, -127.52333577474, -127.52333577474, 
    -127.52333577474, -127.52333577474, -127.52333577474, -127.52333577474, 
    -127.52333577474, -127.52333577474, -127.52333577474, -127.52333577474, 
    -127.52333577474, -127.52333577474, -127.52333577474, -127.52333577474, 
    -127.52333577474, -127.52333577474, -127.52333577474, -127.52333577474, 
    -127.52333577474, -127.52333577474, -127.52333577474, -127.52333577474, 
    -127.52333577474, -127.52333577474, -127.52333577474, -127.52333577474, 
    -127.52333577474, -127.52333577474, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.983334859212, -125.987879897609, 
    -125.983334859212, -125.947621663411, -125.833333333333, 
    -125.958333333333, -125.953334554036, -125.945834477743, 
    -125.983334859212, -126.083333333333, -126.047619047619, 
    -125.983334859212, -126.003334554036, -125.983334859212, 
    -125.987879897609, -126.003334554036, -125.996971361565, 
    -125.983334859212, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.683331807454, -125.678786769058, -125.683331807454, 
    -125.683331807454, -125.71333211263, -125.647618611654, 
    -125.673331197103, -125.799997965495, -125.749997456868, 
    -125.745831807454, -125.683331807454, -125.733331589472, 
    -125.66333211263, -125.683331807454, -125.683331807454, 
    -125.799997965495, -125.653331502279, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.37333577474, -125.333333333333, 
    -125.333333333333, -125.350001017253, -125.3047601609, -125.358334859212, 
    -125.40000406901, -125.233327229818, -125.316665649414, 
    -125.433339436849, -125.283330281576, -125.31333211263, 
    -125.299997965495, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.320832570394, -125.333333333333, 
    -125.333333333333, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.988889906141, -124.983334859212, 
    -124.933333333333, -124.996971361565, -124.988889906142, 
    -124.961906069801, -125.047621227446, -125.133336385091, 
    -125.083333333333, -124.933335622152, -125.000001695421, 
    -124.966668023003, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.683331807454, -124.683331807454, -124.683331807454, 
    -124.683331807454, -124.683331807454, -124.683331807454, 
    -124.683331807454, -124.683331807454, -124.683331807454, 
    -124.683331807454, -124.683331807454, -124.683331807454, 
    -124.753331502279, -124.733332951864, -124.696968309807, 
    -124.733331589472, -124.747618175688, -124.633336385091, 
    -124.799997965495, -124.708331425985, -124.696968309807, 
    -124.683331807454, -124.683331807454, -124.683331807454, 
    -124.683331807454, -124.696968309807, -124.745831807454, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.37333577474, -124.383336385091, 
    -124.383336385091, -124.433339436849, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -123.983334859212, -123.983334859212, 
    -123.983334859212, -123.983334859212, -123.983334859212, 
    -123.983334859212, -123.983334859212, -123.996971361565, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.683331807454, 
    -123.683331807454, -123.683331807454, -123.683331807454, 
    -123.683331807454, -123.683331807454, -123.683331807454, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -122.983334859212, -122.983334859212, -122.983334859212, 
    -122.983334859212, -123.013335164388, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.683331807454, -122.683331807454, 
    -122.696968309807, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.345834096273, -122.345834096273, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.045834859212, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.673329671224, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.033335367839, 
    -121.033335367839, -121.033335367839, -121.033335367839, 
    -121.033335367839, -121.033335367839, -121.033335367839, 
    -121.033335367839, -121.033335367839, -121.033335367839, 
    -121.033335367839, -121.033335367839, -121.083333333333, 
    -121.083333333333, -120.633331298828, -120.633331298828, 
    -120.633331298828, -120.633331298828, -120.633331298828, 
    -120.633331298828, -120.633331298828, -120.633331298828, 
    -120.633331298828, -120.633331298828, -120.645831425985, 
    -120.633331298828, -120.333333333333, -120.333333333333, 
    -120.333333333333, -120.333333333333, -120.333333333333, 
    -120.333333333333, -120.333333333333, -120.333333333333, 
    -120.333333333333, -120.333333333333, -120.320832570394, 
    -120.333333333333, -120.033335367839, -120.033335367839, 
    -120.033335367839, -120.033335367839, -120.033335367839, 
    -120.033335367839, -120.033335367839, -120.033335367839, 
    -120.033335367839, -120.033335367839, -120.033335367839, 
    -120.033335367839, -119.633331298828, -119.633331298828, 
    -119.633331298828, -119.633331298828, -119.633331298828, 
    -119.633331298828, -119.633331298828, -119.633331298828, 
    -119.633331298828, -119.633331298828, -119.633331298828, 
    -119.333333333333, -119.333333333333, -119.333333333333, 
    -119.333333333333, -119.333333333333, -119.333333333333, 
    -119.333333333333, -119.333333333333, -119.333333333333, 
    -119.333333333333, -119.333333333333, -119.033335367839, 
    -119.033335367839, -119.033335367839, -119.033335367839, 
    -119.033335367839, -119.033335367839, -119.033335367839, 
    -119.033335367839, -119.033335367839, -119.033335367839, 
    -119.033335367839, -118.633331298828, -118.633331298828, 
    -118.633331298828, -118.633331298828, -118.633331298828, 
    -118.633331298828, -118.633331298828, -118.633331298828, 
    -118.620831807454, -118.633331298828, -118.333333333333, 
    -118.333333333333, -118.333333333333, -118.333333333333, 
    -118.333333333333, -118.333333333333, -118.333333333333, 
    -118.333333333333, -118.333333333333, -118.033335367839, 
    -118.033335367839, -118.033335367839, -118.033335367839, 
    -118.033335367839, -118.033335367839, -118.033335367839, 
    -118.033335367839, -118.045834859212, -117.633331298828, 
    -117.633331298828, -117.633331298828, -117.633331298828, 
    -117.633331298828, -117.633331298828, -117.661903018043, 
    -117.693330891927, -117.333333333333, -117.333333333333, 
    -117.333333333333, -117.333333333333, -117.333333333333, 
    -117.033335367839, -117.033335367839, -117.033335367839, 
    -117.083333333333, -122.291333516439, -122.291333516439, 
    -122.291333516439, -122.291333516439, -122.291333516439, 
    -122.291333516439, -122.291333516439, -122.291333516439, 
    -122.291333516439, -122.291333516439, -122.291333516439, 
    -122.291333516439, -122.291333516439, -122.291333516439, 
    -122.291333516439, -122.291333516439, -122.291333516439, 
    -122.291333516439, -122.291333516439, -122.291333516439, 
    -122.291333516439, -122.291333516439, -122.291333516439, 
    -122.291333516439, -122.291333516439, -122.291333516439, 
    -122.291333516439, -122.291333516439, -122.291333516439, 
    -122.291333516439, -122.291333516439, -122.291333516439, 
    -122.291333516439, -122.291333516439, -122.291333516439, 
    -122.291333516439, -122.291333516439, -122.291333516439, 
    -122.291333516439, -122.291333516439, -122.291333516439, 
    -122.291333516439, -122.291333516439, -122.291333516439, 
    -122.291333516439, -122.291333516439, -132.340337117513, 
    -132.340337117513, -132.340337117513, -132.340337117513, 
    -132.340337117513, -132.340337117513, -132.340337117513, 
    -132.340337117513, -132.340337117513, -132.340337117513, 
    -132.340337117513, -132.340337117513, -132.340337117513, 
    -132.340337117513, -132.340337117513, -132.340337117513, 
    -132.340337117513, -132.340337117513, -132.340337117513, 
    -132.340337117513, -132.340337117513, -132.340337117513, 
    -132.340337117513, -132.340337117513, -132.340337117513, 
    -132.340337117513, -132.340337117513, -132.340337117513, 
    -132.340337117513, -132.340337117513, -132.340337117513, 
    -132.340337117513, -132.340337117513, -132.340337117513, 
    -132.340337117513, -132.340337117513, -132.340337117513, 
    -132.340337117513, -132.340337117513, -132.340337117513, 
    -132.340337117513, -132.340337117513, -132.340337117513, 
    -132.340337117513, -132.340337117513, -132.340337117513, 
    -125.530331929525, -125.530331929525, -125.530331929525, 
    -125.530331929525, -125.530331929525, -125.530331929525, 
    -125.530331929525, -125.530331929525, -125.530331929525, 
    -125.530331929525, -125.530331929525, -125.530331929525, 
    -125.530331929525, -125.530331929525, -125.530331929525, 
    -125.530331929525, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.983334859212, -126.022223578559, 
    -125.983334859212, -125.933335622152, -125.958333333333, 
    -125.883336385091, -125.961906069801, -125.983334859212, 
    -126.083333333333, -126.047619047619, -126.003334554036, 
    -125.996971361565, -125.983334859212, -125.987879897609, 
    -126.003334554036, -125.996971361565, -125.983334859212, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.678786769058, -125.644443088108, -125.683331807454, 
    -125.71333211263, -125.61666615804, -125.673331197103, -125.833333333333, 
    -125.833333333333, -125.745831807454, -125.783330281576, 
    -125.716664632161, -125.66333211263, -125.683331807454, 
    -125.683331807454, -125.799997965495, -125.653331502279, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.40833791097, 
    -125.433339436849, -125.350001017253, -125.299997965495, -125.3047601609, 
    -125.358334859212, -125.40000406901, -125.233327229818, 
    -125.333333333333, -125.433339436849, -125.283330281576, 
    -125.333333333333, -125.299997965495, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.978789820816, -124.988889906141, 
    -124.973334248861, -124.833333333333, -125.013335164388, 
    -125.033335367839, -125.058335622152, -125.133336385091, 
    -125.083333333333, -124.983334859212, -124.983334859212, 
    -124.966668023003, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.683331807454, -124.683331807454, -124.683331807454, 
    -124.683331807454, -124.683331807454, -124.683331807454, 
    -124.683331807454, -124.683331807454, -124.683331807454, 
    -124.683331807454, -124.683331807454, -124.683331807454, 
    -124.753331502279, -124.733332951864, -124.666664971246, 
    -124.683331807454, -124.783330281576, -124.708331425985, 
    -124.696968309807, -124.683331807454, -124.683331807454, 
    -124.683331807454, -124.683331807454, -124.696968309807, 
    -124.745831807454, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.37333577474, 
    -124.383336385091, -124.383336385091, -124.433339436849, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -123.983334859212, 
    -123.983334859212, -123.983334859212, -123.983334859212, 
    -123.983334859212, -123.983334859212, -123.983334859212, 
    -123.996971361565, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.683331807454, -123.683331807454, -123.683331807454, 
    -123.683331807454, -123.683331807454, -123.683331807454, 
    -123.683331807454, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -122.983334859212, -122.983334859212, 
    -122.983334859212, -122.983334859212, -123.013335164388, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.683331807454, 
    -122.683331807454, -122.696968309807, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.345834096273, -122.345834096273, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.045834859212, -121.633331298828, 
    -121.633331298828, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.633331298828, -121.673329671224, 
    -121.333333333333, -121.333333333333, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.333333333333, 
    -121.033335367839, -121.033335367839, -121.033335367839, 
    -121.033335367839, -121.033335367839, -121.033335367839, 
    -121.033335367839, -121.033335367839, -121.033335367839, 
    -121.033335367839, -121.033335367839, -121.033335367839, 
    -121.083333333333, -121.083333333333, -120.633331298828, 
    -120.633331298828, -120.633331298828, -120.633331298828, 
    -120.633331298828, -120.633331298828, -120.633331298828, 
    -120.633331298828, -120.633331298828, -120.633331298828, 
    -120.645831425985, -120.633331298828, -120.333333333333, 
    -120.333333333333, -120.333333333333, -120.333333333333, 
    -120.333333333333, -120.333333333333, -120.333333333333, 
    -120.333333333333, -120.333333333333, -120.333333333333, 
    -120.320832570394, -120.333333333333, -120.033335367839, 
    -120.033335367839, -120.033335367839, -120.033335367839, 
    -120.033335367839, -120.033335367839, -120.033335367839, 
    -120.033335367839, -120.033335367839, -120.033335367839, 
    -120.033335367839, -120.033335367839, -119.633331298828, 
    -119.633331298828, -119.633331298828, -119.633331298828, 
    -119.633331298828, -119.633331298828, -119.633331298828, 
    -119.633331298828, -119.633331298828, -119.633331298828, 
    -119.633331298828, -119.333333333333, -119.333333333333, 
    -119.333333333333, -119.333333333333, -119.333333333333, 
    -119.333333333333, -119.333333333333, -119.333333333333, 
    -119.333333333333, -119.333333333333, -119.333333333333, 
    -119.033335367839, -119.033335367839, -119.033335367839, 
    -119.033335367839, -119.033335367839, -119.033335367839, 
    -119.033335367839, -119.033335367839, -119.033335367839, 
    -119.033335367839, -119.033335367839, -118.633331298828, 
    -118.633331298828, -118.633331298828, -118.633331298828, 
    -118.633331298828, -118.633331298828, -118.633331298828, 
    -118.633331298828, -118.620831807454, -118.633331298828, 
    -118.333333333333, -118.333333333333, -118.333333333333, 
    -118.333333333333, -118.333333333333, -118.333333333333, 
    -118.333333333333, -118.333333333333, -118.333333333333, 
    -118.033335367839, -118.033335367839, -118.033335367839, 
    -118.033335367839, -118.033335367839, -118.033335367839, 
    -118.033335367839, -118.033335367839, -118.045834859212, 
    -117.633331298828, -117.633331298828, -117.633331298828, 
    -117.633331298828, -117.633331298828, -117.633331298828, 
    -117.661903018043, -117.693330891927, -117.333333333333, 
    -117.333333333333, -117.333333333333, -117.333333333333, 
    -117.333333333333, -117.033335367839, -117.033335367839, 
    -117.033335367839, -117.083333333333, -125.134335835775, 
    -125.134335835775, -125.134335835775, -125.134335835775, 
    -125.134335835775, -125.134335835775, -125.134335835775, 
    -125.134335835775, -125.134335835775, -125.134335835775, 
    -125.134335835775, -125.134335835775, -125.134335835775, 
    -125.072331746419, -125.072331746419, -125.072331746419, 
    -125.072331746419, -125.072331746419, -125.072331746419, 
    -125.072331746419, -125.072331746419, -125.072331746419, 
    -125.072331746419, -125.072331746419, -125.072331746419, 
    -125.072331746419, -125.072331746419, -117.636334737142, 
    -117.636334737142, -117.636334737142, -117.636334737142, 
    -117.636334737142, -117.636334737142, -117.636334737142, 
    -117.636334737142, -117.636334737142, -117.636334737142, 
    -117.636334737142, -117.636334737142, -117.636334737142, 
    -117.636334737142, -117.748334248861, -117.748334248861, 
    -117.748334248861, -117.748334248861, -117.748334248861, 
    -117.748334248861, -117.748334248861, -117.748334248861, 
    -117.748334248861, -117.748334248861, -117.748334248861, 
    -117.748334248861, -117.748334248861, -117.748334248861, 
    -117.748334248861, -117.748334248861, -117.748334248861, 
    -117.748334248861, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.283330281576, -130.283330281576, 
    -130.283330281576, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -130.033335367839, -130.033335367839, -130.033335367839, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.983334859212, -129.983334859212, 
    -129.983334859212, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.633331298828, -129.633331298828, -129.633331298828, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.683331807454, -129.683331807454, 
    -129.683331807454, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.333333333333, -129.333333333333, 
    -129.333333333333, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -129.033335367839, -129.033335367839, -129.033335367839, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.983334859212, -128.983334859212, 
    -128.983334859212, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.633331298828, -128.633331298828, -128.633331298828, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.683331807454, -128.683331807454, 
    -128.683331807454, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.333333333333, -128.333333333333, 
    -128.333333333333, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -128.033335367839, -128.033335367839, -128.033335367839, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.983334859212, -127.983334859212, 
    -127.983334859212, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.633331298828, -127.633331298828, -127.633331298828, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.683331807454, -127.683331807454, 
    -127.683331807454, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.333333333333, -127.333333333333, 
    -127.333333333333, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -127.033335367839, -127.033335367839, -127.033335367839, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.983334859212, -126.983334859212, 
    -126.983334859212, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.633331298828, -126.633331298828, -126.633331298828, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.683331807454, -126.683331807454, 
    -126.683331807454, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.333333333333, -126.333333333333, 
    -126.333333333333, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -126.033335367839, -126.033335367839, -126.033335367839, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.987879897609, -125.983334859212, 
    -125.987879897609, -125.983334859212, -125.996971361565, 
    -125.983334859212, -125.987879897609, -126.019048055013, 
    -125.983334859212, -125.833333333333, -126.083333333333, 
    -126.013335164388, -126.033334096273, -126.022223578559, 
    -125.987879897609, -125.983334859212, -125.983334859212, 
    -125.983334859212, -125.983334859212, -125.983334859212, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.633331298828, 
    -125.633331298828, -125.633331298828, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.696968309807, -125.683331807454, -125.683331807454, 
    -125.678786769058, -125.733333333333, -125.733331589472, 
    -125.695832570394, -125.766662597656, -125.677776760525, 
    -125.783330281576, -125.733331044515, -125.683331807454, 
    -125.658330281576, -125.673332722982, -125.683331807454, 
    -125.683331807454, -125.683331807454, -125.683331807454, 
    -125.683331807454, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.345834096273, -125.333333333333, 
    -125.361906505766, -125.37333577474, -125.433339436849, 
    -125.433339436849, -125.333333333333, -125.299997965495, 
    -125.333333333333, -125.333333333333, -125.333333333333, 
    -125.333333333333, -125.333333333333, -125.345834096273, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -125.033335367839, 
    -125.033335367839, -125.033335367839, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.96969835686, -124.996971361565, -124.970834096273, 
    -124.973334248861, -124.833333333333, -125.133336385091, 
    -124.983334859212, -124.963335164388, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.983334859212, 
    -124.983334859212, -124.983334859212, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.633331298828, -124.633331298828, 
    -124.633331298828, -124.683331807454, -124.683331807454, 
    -124.683331807454, -124.683331807454, -124.683331807454, 
    -124.683331807454, -124.683331807454, -124.683331807454, 
    -124.683331807454, -124.683331807454, -124.683331807454, 
    -124.704760596866, -124.753331502279, -124.766665140788, 
    -124.833333333333, -124.708331425985, -124.696968309807, 
    -124.683331807454, -124.683331807454, -124.683331807454, 
    -124.683331807454, -124.696968309807, -124.745831807454, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.333333333333, -124.333333333333, 
    -124.333333333333, -124.37333577474, -124.383336385091, 
    -124.383336385091, -124.433339436849, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -124.033335367839, -124.033335367839, 
    -124.033335367839, -123.983334859212, -123.983334859212, 
    -123.983334859212, -123.983334859212, -123.983334859212, 
    -123.983334859212, -123.983334859212, -123.996971361565, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.633331298828, 
    -123.633331298828, -123.633331298828, -123.683331807454, 
    -123.683331807454, -123.683331807454, -123.683331807454, 
    -123.683331807454, -123.683331807454, -123.683331807454, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.333333333333, -123.333333333333, 
    -123.333333333333, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -123.033335367839, -123.033335367839, -123.033335367839, 
    -122.983334859212, -122.983334859212, -122.983334859212, 
    -122.983334859212, -123.033335367839, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.633331298828, -122.633331298828, 
    -122.633331298828, -122.683331807454, -122.683331807454, 
    -122.696968309807, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.333333333333, -122.333333333333, -122.333333333333, 
    -122.345834096273, -122.345834096273, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.033335367839, -122.033335367839, -122.033335367839, 
    -122.045834859212, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.633331298828, -121.633331298828, 
    -121.633331298828, -121.673329671224, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.333333333333, 
    -121.333333333333, -121.333333333333, -121.033335367839, 
    -121.033335367839, -121.033335367839, -121.033335367839, 
    -121.033335367839, -121.033335367839, -121.033335367839, 
    -121.033335367839, -121.033335367839, -121.033335367839, 
    -121.033335367839, -121.033335367839, -121.083333333333, 
    -121.083333333333, -120.633331298828, -120.633331298828, 
    -120.633331298828, -120.633331298828, -120.633331298828, 
    -120.633331298828, -120.633331298828, -120.633331298828, 
    -120.633331298828, -120.633331298828, -120.645831425985, 
    -120.633331298828, -120.333333333333, -120.333333333333, 
    -120.333333333333, -120.333333333333, -120.333333333333, 
    -120.333333333333, -120.333333333333, -120.333333333333, 
    -120.333333333333, -120.333333333333, -120.320832570394, 
    -120.333333333333, -120.033335367839, -120.033335367839, 
    -120.033335367839, -120.033335367839, -120.033335367839, 
    -120.033335367839, -120.033335367839, -120.033335367839, 
    -120.033335367839, -120.033335367839, -120.033335367839, 
    -120.033335367839, -119.633331298828, -119.633331298828, 
    -119.633331298828, -119.633331298828, -119.633331298828, 
    -119.633331298828, -119.633331298828, -119.633331298828, 
    -119.633331298828, -119.633331298828, -119.633331298828, 
    -119.333333333333, -119.333333333333, -119.333333333333, 
    -119.333333333333, -119.333333333333, -119.333333333333, 
    -119.333333333333, -119.333333333333, -119.333333333333, 
    -119.333333333333, -119.333333333333, -119.033335367839, 
    -119.033335367839, -119.033335367839, -119.033335367839, 
    -119.033335367839, -119.033335367839, -119.033335367839, 
    -119.033335367839, -119.033335367839, -119.033335367839, 
    -119.033335367839, -118.633331298828, -118.633331298828, 
    -118.633331298828, -118.633331298828, -118.633331298828, 
    -118.633331298828, -118.633331298828, -118.633331298828, 
    -118.620831807454, -118.633331298828, -118.333333333333, 
    -118.333333333333, -118.333333333333, -118.333333333333, 
    -118.333333333333, -118.333333333333, -118.333333333333, 
    -118.333333333333, -118.333333333333, -118.033335367839, 
    -118.033335367839, -118.033335367839, -118.033335367839, 
    -118.033335367839, -118.033335367839, -118.033335367839, 
    -118.033335367839, -118.045834859212, -117.633331298828, 
    -117.633331298828, -117.633331298828, -117.633331298828, 
    -117.633331298828, -117.633331298828, -117.661903018043, 
    -117.693330891927, -117.333333333333, -117.333333333333, 
    -117.333333333333, -117.333333333333, -117.333333333333, 
    -117.033335367839, -117.033335367839, -117.033335367839, 
    -117.083333333333, -118.208333333333, -118.208333333333, 
    -118.208333333333, -118.208333333333, -118.208333333333, 
    -118.208333333333, -118.208333333333, -118.208333333333, 
    -118.208333333333, -118.208333333333, -118.208333333333, 
    -118.208333333333, -118.208333333333, -118.208333333333, 
    -118.208333333333, -118.208333333333, -118.208333333333, 
    -118.208333333333, -118.885335286458, -118.885335286458, 
    -118.885335286458, -118.885335286458, -118.885335286458, 
    -118.885335286458, -118.885335286458, -118.885335286458, 
    -118.885335286458, -118.885335286458, -118.885335286458, 
    -118.885335286458, -118.885335286458, -118.885335286458, 
    -118.885335286458, -118.885335286458, -118.885335286458, 
    -118.885335286458, -118.885335286458, -118.885335286458, 
    -118.885335286458, -118.885335286458, -118.885335286458, 
    -118.885335286458, -118.885335286458, -118.885335286458, 
    -118.885335286458, -118.885335286458, -118.885335286458, 
    -118.885335286458, -133.333333333356, -133.000000000023, 
    -133.333333333356, -132.666666666689, -133.000000000023, 
    -132.333333333356, -132.666666666689, -132.000000000023, 
    -132.333333333356, -133.333333333356, -131.66666666669, 
    -132.000000000023, -133.000000000023, -131.333333333356, 
    -133.333333333356, -131.66666666669, -132.666666666689, 
    -131.000000000023, -133.000000000023, -131.333333333356, 
    -132.333333333356, -133.333333333356, -130.66666666669, 
    -132.666666666689, -131.000000000023, -132.000000000023, 
    -133.000000000023, -130.333333333356, -132.333333333356, 
    -133.333333333356, -130.66666666669, -131.66666666669, -132.666666666689, 
    -130.000000000023, -132.000000000023, -133.000000000023, 
    -130.333333333356, -131.333333333356, -132.333333333356, 
    -129.66666666669, -133.333333333356, -131.66666666669, -132.666666666689, 
    -130.000000000023, -131.000000000023, -132.000000000023, 
    -129.333333333356, -133.000000000023, -131.333333333356, 
    -132.333333333356, -129.66666666669, -133.333333333356, -130.66666666669, 
    -131.66666666669, -129.000000000023, -132.666666666689, 
    -131.000000000023, -132.000000000023, -129.333333333356, 
    -133.000000000023, -130.333333333356, -131.333333333356, 
    -128.66666666669, -132.333333333356, -133.333333333356, -130.66666666669, 
    -131.66666666669, -129.000000000023, -132.666666666689, 
    -130.000000000023, -131.000000000023, -128.333333333357, 
    -132.000000000023, -133.000000000023, -130.333333333356, 
    -131.333333333356, -128.66666666669, -132.333333333356, -129.66666666669, 
    -133.333333333356, -130.66666666669, -128.000000000023, -131.66666666669, 
    -132.666666666689, -130.000000000023, -131.000000000023, 
    -128.333333333357, -132.000000000023, -129.333333333356, 
    -133.000000000023, -130.333333333356, -127.66666666669, 
    -131.333333333356, -132.333333333356, -129.66666666669, 
    -133.333333333356, -130.66666666669, -128.000000000023, -131.66666666669, 
    -129.000000000023, -132.666666666689, -130.000000000023, 
    -127.333333333357, -131.000000000023, -132.000000000023, 
    -129.333333333356, -133.000000000023, -130.333333333356, 
    -127.66666666669, -131.333333333356, -128.66666666669, -132.333333333356, 
    -129.66666666669, -127.000000000023, -133.333333333356, -130.66666666669, 
    -131.66666666669, -129.000000000023, -132.666666666689, 
    -130.000000000023, -127.333333333357, -131.000000000023, 
    -128.333333333357, -132.000000000023, -129.333333333356, 
    -126.66666666669, -133.000000000023, -130.333333333356, 
    -131.333333333356, -128.66666666669, -132.333333333356, -129.66666666669, 
    -127.000000000023, -133.333333333356, -130.66666666669, 
    -128.000000000023, -131.66666666669, -129.000000000023, 
    -126.333333333357, -132.666666666689, -130.000000000023, 
    -131.000000000023, -128.333333333357, -132.000000000023, 
    -129.333333333356, -126.66666666669, -133.000000000023, 
    -130.333333333356, -127.66666666669, -131.333333333356, -128.66666666669, 
    -126.000000000023, -132.333333333356, -129.66666666669, 
    -133.333333333356, -130.66666666669, -128.000000000023, -131.66666666669, 
    -129.000000000023, -126.333333333357, -132.666666666689, 
    -130.000000000023, -127.333333333357, -131.000000000023, 
    -128.333333333357, -125.66666666669, -132.000000000023, 
    -129.333333333356, -133.000000000023, -130.333333333356, 
    -127.66666666669, -131.333333333356, -128.66666666669, -126.000000000023, 
    -132.333333333356, -129.66666666669, -127.000000000023, 
    -133.333333333356, -130.66666666669, -128.000000000023, 
    -125.333333333357, -131.66666666669, -129.000000000023, 
    -132.666666666689, -130.000000000023, -127.333333333357, 
    -131.000000000023, -128.333333333357, -125.66666666669, 
    -132.000000000023, -129.333333333356, -126.66666666669, 
    -133.000000000023, -130.333333333356, -127.66666666669, 
    -125.000000000024, -131.333333333356, -128.66666666669, 
    -132.333333333356, -129.66666666669, -127.000000000023, 
    -133.333333333356, -130.66666666669, -128.000000000023, 
    -125.333333333357, -131.66666666669, -129.000000000023, 
    -126.333333333357, -132.666666666689, -130.000000000023, 
    -127.333333333357, -124.66666666669, -131.000000000023, 
    -128.333333333357, -132.000000000023, -129.333333333356, 
    -126.66666666669, -133.000000000023, -130.333333333356, -127.66666666669, 
    -125.000000000024, -131.333333333356, -128.66666666669, 
    -126.000000000023, -132.333333333356, -129.66666666669, 
    -127.000000000023, -133.333333333356, -124.333333333357, 
    -130.66666666669, -128.000000000023, -131.66666666669, -129.000000000023, 
    -126.333333333357, -132.666666666689, -130.000000000023, 
    -127.333333333357, -124.66666666669, -131.000000000023, 
    -128.333333333357, -125.66666666669, -132.000000000023, 
    -129.333333333356, -126.66666666669, -133.000000000023, 
    -124.000000000024, -130.333333333356, -127.66666666669, 
    -131.333333333356, -128.66666666669, -126.000000000023, 
    -132.333333333356, -129.66666666669, -127.000000000023, 
    -133.333333333356, -124.333333333357, -130.66666666669, 
    -128.000000000023, -125.333333333357, -131.66666666669, 
    -129.000000000023, -126.333333333357, -132.666666666689, 
    -123.66666666669, -130.000000000023, -127.333333333357, 
    -131.000000000023, -128.333333333357, -125.66666666669, 
    -132.000000000023, -129.333333333356, -126.66666666669, 
    -133.000000000023, -124.000000000024, -130.333333333356, 
    -127.66666666669, -125.000000000024, -131.333333333356, -128.66666666669, 
    -126.000000000023, -132.333333333356, -123.333333333357, 
    -129.66666666669, -127.000000000023, -133.333333333356, -130.66666666669, 
    -128.000000000023, -125.333333333357, -131.66666666669, 
    -129.000000000023, -126.333333333357, -132.666666666689, 
    -123.66666666669, -130.000000000023, -127.333333333357, -124.66666666669, 
    -131.000000000023, -128.333333333357, -125.66666666669, 
    -132.000000000023, -123.000000000024, -129.333333333356, 
    -126.66666666669, -133.000000000023, -130.333333333356, -127.66666666669, 
    -125.000000000024, -131.333333333356, -128.66666666669, 
    -126.000000000023, -132.333333333356, -123.333333333357, 
    -129.66666666669, -127.000000000023, -133.333333333356, 
    -124.333333333357, -130.66666666669, -128.000000000023, 
    -125.333333333357, -131.66666666669, -122.66666666669, -129.000000000023, 
    -126.333333333357, -132.666666666689, -130.000000000023, 
    -127.333333333357, -124.66666666669, -131.000000000023, 
    -128.333333333357, -125.66666666669, -132.000000000023, 
    -123.000000000024, -129.333333333356, -126.66666666669, 
    -133.000000000023, -124.000000000024, -130.333333333356, 
    -127.66666666669, -125.000000000024, -131.333333333356, 
    -122.333333333357, -128.66666666669, -126.000000000023, 
    -132.333333333356, -129.66666666669, -127.000000000023, 
    -133.333333333356, -124.333333333357, -130.66666666669, 
    -128.000000000023, -125.333333333357, -131.66666666669, -122.66666666669, 
    -129.000000000023, -126.333333333357, -132.666666666689, 
    -123.66666666669, -130.000000000023, -127.333333333357, -124.66666666669, 
    -131.000000000023, -122.000000000024, -128.333333333357, 
    -125.66666666669, -132.000000000023, -129.333333333356, -126.66666666669, 
    -133.000000000023, -124.000000000024, -130.333333333356, 
    -127.66666666669, -125.000000000024, -131.333333333356, 
    -122.333333333357, -128.66666666669, -126.000000000023, 
    -132.333333333356, -123.333333333357, -129.66666666669, 
    -127.000000000023, -133.333333333356, -124.333333333357, 
    -130.66666666669, -121.666666666691, -128.000000000023, 
    -125.333333333357, -131.66666666669, -129.000000000023, 
    -126.333333333357, -132.666666666689, -123.66666666669, 
    -130.000000000023, -127.333333333357, -124.66666666669, 
    -131.000000000023, -122.000000000024, -128.333333333357, 
    -125.66666666669, -132.000000000023, -123.000000000024, 
    -129.333333333356, -126.66666666669, -133.000000000023, 
    -124.000000000024, -130.333333333356, -121.333333333357, 
    -127.66666666669, -125.000000000024, -131.333333333356, -128.66666666669, 
    -126.000000000023, -132.333333333356, -123.333333333357, 
    -129.66666666669, -127.000000000023, -133.333333333356, 
    -124.333333333357, -130.66666666669, -121.666666666691, 
    -128.000000000023, -125.333333333357, -131.66666666669, -122.66666666669, 
    -129.000000000023, -126.333333333357, -132.666666666689, 
    -123.66666666669, -130.000000000023, -121.000000000024, 
    -127.333333333357, -124.66666666669, -131.000000000023, 
    -128.333333333357, -125.66666666669, -132.000000000023, 
    -123.000000000024, -129.333333333356, -126.66666666669, 
    -133.000000000023, -124.000000000024, -130.333333333356, 
    -121.333333333357, -127.66666666669, -125.000000000024, 
    -131.333333333356, -122.333333333357, -128.66666666669, 
    -126.000000000023, -132.333333333356, -123.333333333357, 
    -129.66666666669, -120.666666666691, -127.000000000023, 
    -133.333333333356, -124.333333333357, -130.66666666669, 
    -128.000000000023, -125.333333333357, -131.66666666669, -122.66666666669, 
    -129.000000000023, -126.333333333357, -132.666666666689, 
    -123.66666666669, -130.000000000023, -121.000000000024, 
    -127.333333333357, -124.66666666669, -131.000000000023, 
    -122.000000000024, -128.333333333357, -125.66666666669, 
    -132.000000000023, -123.000000000024, -129.333333333356, 
    -120.333333333357, -126.66666666669, -133.000000000023, 
    -124.000000000024, -130.333333333356, -127.66666666669, 
    -125.000000000024, -131.333333333356, -122.333333333357, 
    -128.66666666669, -126.000000000023, -132.333333333356, 
    -123.333333333357, -129.66666666669, -120.666666666691, 
    -127.000000000023, -133.333333333356, -124.333333333357, 
    -130.66666666669, -121.666666666691, -128.000000000023, 
    -125.333333333357, -131.666666666689, -122.66666666669, 
    -129.000000000023, -120.000000000024, -126.333333333357, 
    -132.666666666689, -123.66666666669, -130.000000000023, 
    -127.333333333357, -124.66666666669, -131.000000000023, 
    -122.000000000024, -128.333333333357, -125.66666666669, 
    -132.000000000023, -123.000000000024, -129.333333333356, 
    -120.333333333357, -126.66666666669, -133.000000000023, 
    -124.000000000024, -130.333333333356, -121.333333333357, 
    -127.66666666669, -125.000000000024, -131.333333333356, 
    -122.333333333357, -128.66666666669, -119.666666666691, 
    -126.000000000023, -132.333333333356, -123.333333333357, 
    -129.66666666669, -127.000000000023, -133.333333333356, 
    -124.333333333357, -130.66666666669, -121.666666666691, 
    -128.000000000023, -125.333333333357, -131.66666666669, -122.66666666669, 
    -129.000000000023, -120.000000000024, -126.333333333357, 
    -132.666666666689, -123.66666666669, -130.000000000023, 
    -121.000000000024, -127.333333333357, -124.66666666669, 
    -131.000000000023, -122.000000000024, -128.333333333357, 
    -119.333333333357, -125.66666666669, -132.000000000023, 
    -123.000000000024, -129.333333333356, -126.66666666669, 
    -133.000000000023, -124.000000000024, -130.333333333356, 
    -121.333333333357, -127.66666666669, -125.000000000024, 
    -131.333333333356, -122.333333333357, -128.66666666669, 
    -119.666666666691, -126.000000000023, -132.333333333356, 
    -123.333333333357, -129.66666666669, -120.666666666691, 
    -127.000000000023, -133.333333333356, -124.333333333357, 
    -130.66666666669, -121.666666666691, -128.000000000023, 
    -119.000000000024, -125.333333333357, -131.666666666689, 
    -122.66666666669, -129.000000000023, -126.333333333357, 
    -132.666666666689, -123.66666666669, -130.000000000023, 
    -121.000000000024, -127.333333333357, -124.66666666669, 
    -131.000000000023, -122.000000000024, -128.333333333357, 
    -119.333333333357, -125.66666666669, -132.000000000023, 
    -123.000000000024, -129.333333333356, -120.333333333357, 
    -126.66666666669, -133.000000000023, -124.000000000024, 
    -130.333333333356, -121.333333333357, -127.66666666669, 
    -118.666666666691, -125.000000000024, -131.333333333356, 
    -122.333333333357, -128.66666666669, -126.000000000023, 
    -132.333333333356, -123.333333333357, -129.66666666669, 
    -120.666666666691, -127.000000000023, -133.333333333356, 
    -124.333333333357, -130.66666666669, -121.666666666691, 
    -128.000000000023, -119.000000000024, -125.333333333357, 
    -131.66666666669, -122.66666666669, -129.000000000023, -120.000000000024, 
    -126.333333333357, -132.666666666689, -123.66666666669, 
    -130.000000000023, -121.000000000024, -127.333333333357, 
    -118.333333333358, -124.66666666669, -131.000000000023, 
    -122.000000000024, -128.333333333357, -125.66666666669, 
    -132.000000000023, -123.000000000024, -129.333333333356, 
    -120.333333333357, -126.66666666669, -133.000000000023, 
    -124.000000000024, -130.333333333356, -121.333333333357, 
    -127.66666666669, -118.666666666691, -125.000000000024, 
    -131.333333333356, -122.333333333357, -128.66666666669, 
    -119.666666666691, -126.000000000023, -132.333333333356, 
    -123.333333333357, -129.66666666669, -120.666666666691, 
    -127.000000000023, -133.333333333356, -118.000000000024, 
    -124.333333333357, -130.66666666669, -121.666666666691, 
    -128.000000000023, -125.333333333357, -131.66666666669, -122.66666666669, 
    -129.000000000023, -120.000000000024, -126.333333333357, 
    -132.666666666689, -123.66666666669, -130.000000000023, 
    -121.000000000024, -127.333333333357, -118.333333333358, 
    -124.66666666669, -131.000000000023, -122.000000000024, 
    -128.333333333357, -119.333333333357, -125.66666666669, 
    -132.000000000023, -123.000000000024, -129.333333333356, 
    -120.333333333357, -126.66666666669, -133.000000000023, 
    -117.666666666691, -124.000000000024, -130.333333333356, 
    -121.333333333357, -127.66666666669, -125.000000000024, 
    -131.333333333356, -122.333333333357, -128.66666666669, 
    -119.666666666691, -126.000000000023, -132.333333333356, 
    -123.333333333357, -129.66666666669, -120.666666666691, 
    -127.000000000023, -133.333333333356, -118.000000000024, 
    -124.333333333357, -130.66666666669, -121.666666666691, 
    -128.000000000023, -119.000000000024, -125.333333333357, 
    -131.66666666669, -122.66666666669, -129.000000000023, -120.000000000024, 
    -126.333333333357, -132.666666666689, -117.333333333358, 
    -123.66666666669, -130.000000000023, -121.000000000024, 
    -127.333333333357, -124.66666666669, -131.000000000023, 
    -122.000000000024, -128.333333333357, -119.333333333357, 
    -125.66666666669, -132.000000000023, -123.000000000024, 
    -129.333333333356, -120.333333333357, -126.66666666669, 
    -133.000000000023, -117.666666666691, -124.000000000024, 
    -130.333333333356, -121.333333333357, -127.66666666669, 
    -118.666666666691, -125.000000000024, -131.333333333356, 
    -122.333333333357, -128.66666666669, -119.666666666691, 
    -126.000000000023, -132.333333333356, -117.000000000024, 
    -123.333333333357, -129.66666666669, -120.666666666691, 
    -127.000000000023, -133.333333333356, -124.333333333357, 
    -130.66666666669, -121.666666666691, -128.000000000023, 
    -119.000000000024, -125.333333333357, -131.66666666669, -122.66666666669, 
    -129.000000000023, -120.000000000024, -126.333333333357, 
    -132.666666666689, -117.333333333358, -123.66666666669, 
    -130.000000000023, -121.000000000024, -127.333333333357, 
    -118.333333333358, -124.66666666669, -131.000000000023, 
    -122.000000000024, -128.333333333357, -119.333333333357, 
    -125.66666666669, -132.000000000023, -123.000000000024, 
    -129.333333333356, -120.333333333357, -126.66666666669, 
    -133.000000000023, -124.000000000024, -130.333333333356, 
    -121.333333333357, -127.66666666669, -118.666666666691, 
    -125.000000000024, -131.333333333356, -122.333333333357, 
    -128.66666666669, -119.666666666691, -126.000000000023, 
    -132.333333333356, -117.000000000024, -123.333333333357, 
    -129.66666666669, -120.666666666691, -127.000000000023, 
    -133.333333333356, -118.000000000024, -124.333333333357, 
    -130.66666666669, -121.666666666691, -128.000000000023, 
    -119.000000000024, -125.333333333357, -131.66666666669, -122.66666666669, 
    -129.000000000023, -120.000000000024, -126.333333333357, 
    -132.666666666689, -123.66666666669, -130.000000000023, 
    -121.000000000024, -127.333333333357, -118.333333333358, 
    -124.66666666669, -131.000000000023, -122.000000000024, 
    -128.333333333357, -119.333333333357, -125.66666666669, 
    -132.000000000023, -123.000000000024, -129.333333333356, 
    -120.333333333357, -126.66666666669, -133.000000000023, 
    -117.666666666691, -124.000000000024, -130.333333333356, 
    -121.333333333357, -127.66666666669, -118.666666666691, 
    -125.000000000024, -131.333333333356, -122.333333333357, 
    -128.66666666669, -119.666666666691, -126.000000000023, 
    -132.333333333356, -123.333333333357, -129.66666666669, 
    -120.666666666691, -127.000000000023, -133.333333333356, 
    -118.000000000024, -124.333333333357, -130.66666666669, 
    -121.666666666691, -128.000000000023, -119.000000000024, 
    -125.333333333357, -131.66666666669, -122.66666666669, -129.000000000023, 
    -120.000000000024, -126.333333333357, -132.666666666689, 
    -117.333333333358, -123.66666666669, -130.000000000023, 
    -121.000000000024, -127.333333333357, -118.333333333358, 
    -124.66666666669, -131.000000000023, -122.000000000024, 
    -128.333333333357, -119.333333333357, -125.66666666669, 
    -132.000000000023, -123.000000000024, -129.333333333356, 
    -120.333333333357, -126.66666666669, -133.000000000023, 
    -117.666666666691, -124.000000000024, -130.333333333356, 
    -121.333333333357, -127.66666666669, -118.666666666691, 
    -125.000000000024, -131.333333333356, -122.333333333357, 
    -128.66666666669, -119.666666666691, -126.000000000023, 
    -132.333333333356, -123.333333333357, -129.66666666669, 
    -120.666666666691, -127.000000000023, -133.333333333356, 
    -118.000000000024, -124.333333333357, -130.66666666669, 
    -121.666666666691, -128.000000000023, -119.000000000024, 
    -125.333333333357, -131.66666666669, -122.66666666669, -129.000000000023, 
    -120.000000000024, -126.333333333357, -132.666666666689, 
    -123.66666666669, -130.000000000023, -121.000000000024, 
    -127.333333333357, -124.66666666669, -131.000000000023, 
    -122.000000000024, -128.333333333357, -119.333333333357, 
    -125.66666666669, -132.000000000023, -123.000000000024, 
    -129.333333333356, -120.333333333357, -126.66666666669, 
    -133.000000000023, -117.666666666691, -124.000000000024, 
    -130.333333333356, -121.333333333357, -127.66666666669, 
    -118.666666666691, -125.000000000024, -131.333333333356, 
    -122.333333333357, -128.66666666669, -126.000000000023, 
    -132.333333333356, -123.333333333357, -129.66666666669, 
    -127.000000000023, -133.333333333356, -124.333333333357, 
    -130.66666666669, -121.666666666691, -128.000000000023, 
    -119.000000000024, -125.333333333357, -131.66666666669, -122.66666666669, 
    -129.000000000023, -120.000000000024, -126.333333333357, 
    -132.666666666689, -123.66666666669, -130.000000000023, 
    -121.000000000024, -127.333333333357, -124.66666666669, 
    -131.000000000023, -122.000000000024, -128.333333333357, 
    -125.66666666669, -132.000000000023, -123.000000000024, 
    -129.333333333356, -126.66666666669, -133.000000000023, 
    -124.000000000024, -130.333333333356, -121.333333333357, 
    -127.66666666669, -118.666666666691, -125.000000000024, 
    -131.333333333356, -122.333333333357, -128.66666666669, 
    -126.000000000023, -132.333333333356, -123.333333333357, 
    -129.66666666669, -127.000000000023, -133.333333333356, 
    -124.333333333357, -130.66666666669, -121.666666666691, 
    -128.000000000023, -125.333333333357, -131.66666666669, -122.66666666669, 
    -129.000000000023, -126.333333333357, -132.666666666689, 
    -123.66666666669, -130.000000000023, -127.333333333357, -124.66666666669, 
    -131.000000000023, -122.000000000024, -128.333333333357, 
    -125.66666666669, -132.000000000023, -123.000000000024, 
    -129.333333333356, -126.66666666669, -133.000000000023, 
    -124.000000000024, -130.333333333356, -127.66666666669, 
    -125.000000000024, -131.333333333356, -122.333333333357, 
    -128.66666666669, -126.000000000023, -132.333333333356, 
    -123.333333333357, -129.66666666669, -127.000000000023, 
    -133.333333333356, -124.333333333357, -130.66666666669, 
    -128.000000000023, -125.333333333357, -131.66666666669, -122.66666666669, 
    -129.000000000023, -126.333333333357, -132.666666666689, 
    -123.66666666669, -130.000000000023, -127.333333333357, -124.66666666669, 
    -131.000000000023, -128.333333333357, -125.66666666669, 
    -132.000000000023, -123.000000000024, -129.333333333356, 
    -126.66666666669, -133.000000000023, -124.000000000024, 
    -130.333333333356, -127.66666666669, -125.000000000024, 
    -131.333333333356, -122.333333333357, -128.66666666669, 
    -126.000000000023, -132.333333333356, -123.333333333357, 
    -129.66666666669, -127.000000000023, -133.333333333356, 
    -124.333333333357, -130.66666666669, -128.000000000023, 
    -125.333333333357, -131.66666666669, -122.66666666669, -129.000000000023, 
    -126.333333333357, -132.666666666689, -123.66666666669, 
    -130.000000000023, -127.333333333357, -124.66666666669, 
    -131.000000000023, -128.333333333357, -125.66666666669, 
    -132.000000000023, -123.000000000024, -129.333333333356, 
    -126.66666666669, -133.000000000023, -124.000000000024, 
    -130.333333333356, -127.66666666669, -125.000000000024, 
    -131.333333333356, -128.66666666669, -126.000000000023, 
    -132.333333333356, -123.333333333357, -129.66666666669, 
    -127.000000000023, -133.333333333356, -124.333333333357, 
    -130.66666666669, -128.000000000023, -125.333333333357, -131.66666666669, 
    -129.000000000023, -126.333333333357, -132.666666666689, 
    -123.66666666669, -130.000000000023, -127.333333333357, -124.66666666669, 
    -131.000000000023, -128.333333333357, -125.66666666669, 
    -132.000000000023, -123.000000000024, -129.333333333356, 
    -126.66666666669, -133.000000000023, -124.000000000024, 
    -130.333333333356, -127.66666666669, -125.000000000024, 
    -131.333333333356, -128.66666666669, -126.000000000023, 
    -132.333333333356, -129.66666666669, -127.000000000023, 
    -133.333333333356, -124.333333333357, -130.66666666669, 
    -128.000000000023, -125.333333333357, -131.66666666669, 
    -129.000000000023, -126.333333333357, -132.666666666689, 
    -130.000000000023, -127.333333333357, -124.66666666669, 
    -131.000000000023, -128.333333333357, -125.66666666669, 
    -132.000000000023, -129.333333333356, -126.66666666669, 
    -133.000000000023, -124.000000000024, -130.333333333356, 
    -127.66666666669, -125.000000000024, -131.333333333356, -128.66666666669, 
    -126.000000000023, -132.333333333356, -129.66666666669, 
    -127.000000000023, -133.333333333356, -124.333333333357, 
    -130.66666666669, -128.000000000023, -125.333333333357, -131.66666666669, 
    -129.000000000023, -126.333333333357, -132.666666666689, 
    -130.000000000023, -127.333333333357, -124.66666666669, 
    -131.000000000023, -128.333333333357, -125.66666666669, 
    -132.000000000023, -129.333333333356, -126.66666666669, 
    -133.000000000023, -130.333333333356, -127.66666666669, 
    -125.000000000024, -131.333333333356, -128.66666666669, 
    -126.000000000023, -132.333333333356, -129.66666666669, 
    -127.000000000023, -133.333333333356, -124.333333333357, 
    -130.66666666669, -128.000000000023, -125.333333333357, -131.66666666669, 
    -129.000000000023, -126.333333333357, -132.666666666689, 
    -130.000000000023, -127.333333333357, -124.66666666669, 
    -131.000000000023, -128.333333333357, -125.66666666669, 
    -132.000000000023, -129.333333333356, -126.66666666669, 
    -133.000000000023, -130.333333333356, -127.66666666669, 
    -125.000000000024, -131.333333333356, -128.66666666669, 
    -126.000000000023, -132.333333333356, -129.66666666669, 
    -127.000000000023, -133.333333333356, -124.333333333357, 
    -130.66666666669, -128.000000000023, -125.333333333357, -131.66666666669, 
    -129.000000000023, -126.333333333357, -132.666666666689, 
    -130.000000000023, -127.333333333357, -124.66666666669, 
    -131.000000000023, -128.333333333357, -125.66666666669, 
    -132.000000000023, -129.333333333356, -126.66666666669, 
    -133.000000000023, -130.333333333356, -127.66666666669, 
    -125.000000000024, -131.333333333356, -128.66666666669, 
    -126.000000000023, -132.333333333356, -129.66666666669, 
    -127.000000000023, -133.333333333356, -130.66666666669, 
    -128.000000000023, -125.333333333357, -131.66666666669, 
    -129.000000000023, -126.333333333357, -132.666666666689, 
    -130.000000000023, -127.333333333357, -131.000000000023, 
    -128.333333333357, -125.66666666669, -132.000000000023, 
    -129.333333333356, -126.66666666669, -133.000000000023, 
    -130.333333333356, -127.66666666669, -125.000000000024, 
    -131.333333333356, -128.66666666669, -126.000000000023, 
    -132.333333333356, -129.66666666669, -127.000000000023, 
    -133.333333333356, -130.66666666669, -128.000000000023, 
    -125.333333333357, -131.66666666669, -129.000000000023, 
    -126.333333333357, -132.666666666689, -130.000000000023, 
    -127.333333333357, -124.66666666669, -131.000000000023, 
    -128.333333333357, -125.66666666669, -132.000000000023, 
    -129.333333333356, -126.66666666669, -133.000000000023, 
    -130.333333333356, -127.66666666669, -125.000000000024, 
    -131.333333333356, -128.66666666669, -126.000000000023, 
    -132.333333333356, -129.66666666669, -127.000000000023, 
    -133.333333333356, -130.66666666669, -128.000000000023, 
    -125.333333333357, -131.66666666669, -129.000000000023, 
    -126.333333333357, -132.666666666689, -130.000000000023, 
    -127.333333333357, -124.66666666669, -131.000000000023, 
    -128.333333333357, -125.66666666669, -132.000000000023, 
    -129.333333333356, -126.66666666669, -133.000000000023, 
    -130.333333333356, -127.66666666669, -131.333333333356, -128.66666666669, 
    -126.000000000023, -132.333333333356, -129.66666666669, 
    -127.000000000023, -133.333333333356, -130.66666666669, 
    -128.000000000023, -125.333333333357, -131.66666666669, 
    -129.000000000023, -126.333333333357, -132.666666666689, 
    -130.000000000023, -127.333333333357, -131.000000000023, 
    -128.333333333357, -125.66666666669, -132.000000000023, 
    -129.333333333356, -126.66666666669, -133.000000000023, 
    -130.333333333356, -127.66666666669, -131.333333333356, -128.66666666669, 
    -126.000000000023, -132.333333333356, -129.66666666669, 
    -127.000000000023, -133.333333333356, -130.66666666669, 
    -128.000000000023, -125.333333333357, -131.66666666669, 
    -129.000000000023, -126.333333333357, -132.666666666689, 
    -130.000000000023, -127.333333333357, -131.000000000023, 
    -128.333333333357, -125.66666666669, -132.000000000023, 
    -129.333333333356, -126.66666666669, -133.000000000023, 
    -130.333333333356, -127.66666666669, -131.333333333356, -128.66666666669, 
    -126.000000000023, -132.333333333356, -129.66666666669, 
    -127.000000000023, -130.66666666669, -128.000000000023, 
    -125.333333333357, -131.66666666669, -129.000000000023, 
    -126.333333333357, -132.666666666689, -130.000000000023, 
    -127.333333333357, -131.000000000023, -128.333333333357, 
    -125.66666666669, -132.000000000023, -129.333333333356, -126.66666666669, 
    -130.333333333356, -127.66666666669, -125.000000000024, 
    -131.333333333356, -128.66666666669, -126.000000000023, 
    -132.333333333356, -129.66666666669, -127.000000000023, -130.66666666669, 
    -128.000000000023, -125.333333333357, -131.66666666669, 
    -129.000000000023, -126.333333333357, -130.000000000023, 
    -127.333333333357, -131.000000000023, -128.333333333357, 
    -125.66666666669, -132.000000000023, -129.333333333356, -126.66666666669, 
    -130.333333333356, -127.66666666669, -125.000000000024, 
    -131.333333333356, -128.66666666669, -126.000000000023, -129.66666666669, 
    -127.000000000023, -130.66666666669, -128.000000000023, 
    -125.333333333357, -131.66666666669, -129.000000000023, 
    -126.333333333357, -130.000000000023, -127.333333333357, 
    -131.000000000023, -128.333333333357, -125.66666666669, 
    -129.333333333356, -126.66666666669, -130.333333333356, -127.66666666669, 
    -125.000000000024, -131.333333333356, -128.66666666669, 
    -126.000000000023, -129.66666666669, -127.000000000023, -130.66666666669, 
    -128.000000000023, -125.333333333357, -129.000000000023, 
    -126.333333333357, -130.000000000023, -127.333333333357, 
    -131.000000000023, -128.333333333357, -125.66666666669, 
    -129.333333333356, -126.66666666669, -130.333333333356, -127.66666666669, 
    -125.000000000024, -128.66666666669, -126.000000000023, -129.66666666669, 
    -127.000000000023, -130.66666666669, -128.000000000023, 
    -125.333333333357, -129.000000000023, -126.333333333357, 
    -130.000000000023, -127.333333333357, -128.333333333357, 
    -125.66666666669, -129.333333333356, -126.66666666669, -130.333333333356, 
    -127.66666666669, -125.000000000024, -128.66666666669, -126.000000000023, 
    -129.66666666669, -127.000000000023, -128.000000000023, 
    -125.333333333357, -129.000000000023, -126.333333333357, 
    -130.000000000023, -127.333333333357, -124.66666666669, 
    -128.333333333357, -125.66666666669, -129.333333333356, -126.66666666669, 
    -127.66666666669, -125.000000000024, -128.66666666669, -126.000000000023, 
    -129.66666666669, -127.000000000023, -128.000000000023, 
    -125.333333333357, -129.000000000023, -126.333333333357, 
    -127.333333333357, -124.66666666669, -128.333333333357, -125.66666666669, 
    -129.333333333356, -126.66666666669, -127.66666666669, -125.000000000024, 
    -128.66666666669, -126.000000000023, -127.000000000023, 
    -128.000000000023, -125.333333333357, -129.000000000023, 
    -126.333333333357, -127.333333333357, -124.66666666669, 
    -128.333333333357, -125.66666666669, -126.66666666669, -127.66666666669, 
    -125.000000000024, -128.66666666669, -126.000000000023, 
    -127.000000000023, -128.000000000023, -125.333333333357, 
    -126.333333333357, -127.333333333357, -124.66666666669, 
    -128.333333333357, -125.66666666669, -126.66666666669, -127.66666666669, 
    -125.000000000024, -126.000000000023, -127.000000000023, 
    -128.000000000023, -125.333333333357, -126.333333333357, 
    -127.333333333357, -124.66666666669, -125.66666666669, -126.66666666669, 
    -127.66666666669, -125.000000000024, -126.000000000023, 
    -127.000000000023, -125.333333333357, -126.333333333357, 
    -127.333333333357, -124.66666666669, -125.66666666669, -126.66666666669, 
    -125.000000000024, -126.000000000023, -127.000000000023, 
    -124.333333333357, -125.333333333357, -126.333333333357, 
    -124.66666666669, -125.66666666669, -126.66666666669, -125.000000000024, 
    -126.000000000023, -124.333333333357, -125.333333333357, 
    -126.333333333357, -124.66666666669, -125.66666666669, -125.000000000024, 
    -126.000000000023, -124.333333333357, -125.333333333357, 
    -124.66666666669, -125.66666666669, -125.000000000024, -125.333333333357, 
    -124.66666666669, -125.000000000024, -124.333333333357, -124.66666666669 ;

 obs_lat = 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3666661580404, 38.6666666666667, 38.966667175293, 
    39.3666661580404, 39.6666666666667, 39.966667175293, 40.3666661580404, 
    40.6666666666667, 40.966667175293, 41.3666661580404, 41.6666666666667, 
    41.966667175293, 42.3666661580404, 42.6666666666667, 42.966667175293, 
    43.3666661580404, 43.6666666666667, 43.966667175293, 44.3666661580404, 
    44.6666666666667, 44.966667175293, 45.3666661580404, 45.6666666666667, 
    45.966667175293, 46.3666661580404, 46.6666666666667, 46.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.966667175293, 41.3666661580404, 41.6666666666667, 41.966667175293, 
    42.3666661580404, 42.6666666666667, 42.966667175293, 43.3666661580404, 
    43.6666666666667, 43.966667175293, 44.3666661580404, 44.6666666666667, 
    44.966667175293, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    39.966667175293, 40.3666661580404, 40.6666666666667, 40.966667175293, 
    41.3666661580404, 41.6666666666667, 41.966667175293, 42.3666661580404, 
    42.6666666666667, 42.966667175293, 43.3666661580404, 43.6666666666667, 
    43.966667175293, 44.3666661580404, 44.6666666666667, 44.966667175293, 
    45.3666661580404, 45.6666666666667, 45.966667175293, 46.3666661580404, 
    46.6666666666667, 46.966667175293, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 38.3666661580404, 38.6666666666667, 
    38.966667175293, 39.3666661580404, 39.6666666666667, 39.966667175293, 
    40.3666661580404, 40.6666666666667, 40.966667175293, 41.3666661580404, 
    41.6666666666667, 41.966667175293, 42.3666661580404, 42.6666666666667, 
    42.966667175293, 43.3666661580404, 43.6666666666667, 43.966667175293, 
    44.3666661580404, 44.6666666666667, 44.966667175293, 45.3666661580404, 
    45.6666666666667, 45.966667175293, 46.3666661580404, 46.6666666666667, 
    46.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3666661580404, 38.6666666666667, 38.966667175293, 
    39.3666661580404, 39.6666666666667, 39.966667175293, 40.3666661580404, 
    40.6666666666667, 40.966667175293, 41.3666661580404, 41.6666666666667, 
    41.966667175293, 42.3666661580404, 42.6666666666667, 42.966667175293, 
    43.3666661580404, 43.6666666666667, 43.966667175293, 44.3666661580404, 
    44.6666666666667, 44.966667175293, 45.3666661580404, 45.6666666666667, 
    45.966667175293, 46.3666661580404, 46.6666666666667, 46.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.966667175293, 41.3666661580404, 41.6666666666667, 41.966667175293, 
    42.3666661580404, 42.6666666666667, 42.966667175293, 43.3666661580404, 
    43.6666666666667, 43.966667175293, 44.3666661580404, 44.6666666666667, 
    44.966667175293, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    39.966667175293, 40.3666661580404, 40.6666666666667, 40.966667175293, 
    41.3666661580404, 41.6666666666667, 41.966667175293, 42.3666661580404, 
    42.6666666666667, 42.966667175293, 43.3666661580404, 43.6666666666667, 
    43.966667175293, 44.3666661580404, 44.6666666666667, 44.966667175293, 
    45.3666661580404, 45.6666666666667, 45.966667175293, 46.3666661580404, 
    46.6666666666667, 46.966667175293, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 38.3666661580404, 38.6666666666667, 
    38.966667175293, 39.3666661580404, 39.6666666666667, 39.966667175293, 
    40.3666661580404, 40.6666666666667, 40.966667175293, 41.3666661580404, 
    41.6666666666667, 41.966667175293, 42.3666661580404, 42.6666666666667, 
    42.966667175293, 43.3666661580404, 43.6666666666667, 43.966667175293, 
    44.3666661580404, 44.6666666666667, 44.966667175293, 45.3666661580404, 
    45.6666666666667, 45.966667175293, 46.3666661580404, 46.6666666666667, 
    46.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3666661580404, 38.6666666666667, 38.966667175293, 
    39.3666661580404, 39.6666666666667, 39.966667175293, 40.3666661580404, 
    40.6666666666667, 40.966667175293, 41.3666661580404, 41.6666666666667, 
    41.966667175293, 42.3666661580404, 42.6666666666667, 42.966667175293, 
    43.3666661580404, 43.6666666666667, 43.966667175293, 44.3666661580404, 
    44.6666666666667, 44.966667175293, 45.3666661580404, 45.6666666666667, 
    45.966667175293, 46.3666661580404, 46.6666666666667, 46.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.966667175293, 41.3666661580404, 41.6666666666667, 41.966667175293, 
    42.3666661580404, 42.6666666666667, 42.966667175293, 43.3666661580404, 
    43.6666666666667, 43.966667175293, 44.3666661580404, 44.6666666666667, 
    44.966667175293, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    39.966667175293, 40.3666661580404, 40.6666666666667, 40.966667175293, 
    41.3666661580404, 41.6666666666667, 41.966667175293, 42.3666661580404, 
    42.6666666666667, 42.966667175293, 43.3666661580404, 43.6666666666667, 
    43.966667175293, 44.3666661580404, 44.6666666666667, 44.966667175293, 
    45.3666661580404, 45.6666666666667, 45.966667175293, 46.3666661580404, 
    46.6666666666667, 46.966667175293, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 38.3666661580404, 38.6666666666667, 
    38.966667175293, 39.3666661580404, 39.6666666666667, 39.966667175293, 
    40.3666661580404, 40.6666666666667, 40.966667175293, 41.3666661580404, 
    41.6666666666667, 41.966667175293, 42.3666661580404, 42.6666666666667, 
    42.966667175293, 43.3666661580404, 43.6666666666667, 43.966667175293, 
    44.3666661580404, 44.6666666666667, 44.966667175293, 45.3666661580404, 
    45.6666666666667, 45.966667175293, 46.3666661580404, 46.6666666666667, 
    46.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3666661580404, 38.6666666666667, 38.966667175293, 
    39.3666661580404, 39.6666666666667, 39.966667175293, 40.3666661580404, 
    40.6666666666667, 40.966667175293, 41.3666661580404, 41.6666666666667, 
    41.966667175293, 42.3666661580404, 42.6666666666667, 42.966667175293, 
    43.3666661580404, 43.6666666666667, 43.966667175293, 44.3666661580404, 
    44.6666666666667, 44.966667175293, 45.3666661580404, 45.6666666666667, 
    45.966667175293, 46.3666661580404, 46.6666666666667, 46.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.966667175293, 41.3666661580404, 41.6757574370413, 41.966667175293, 
    42.3523802984328, 42.5666681925456, 42.9952385312035, 43.3666659037272, 
    43.6291672388713, 43.966667175293, 44.3666661580404, 44.6809521629697, 
    44.966667175293, 45.3566660563151, 45.6666666666667, 45.9666672908899, 
    46.3757571596088, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    39.966667175293, 40.3666661580404, 40.6666666666667, 40.966667175293, 
    41.3575752720688, 41.6666666666667, 41.966667175293, 42.3666659037272, 
    42.6380956740606, 42.9666670481364, 43.3999989827474, 43.6999994913737, 
    43.9541670481364, 44.7666651407878, 44.9666675385975, 45.3666659037272, 
    45.6666666666667, 45.966667175293, 46.3666664759318, 46.6666666666667, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.966667175293, 41.3666661580404, 41.6666666666667, 41.9333337148031, 
    42.3809518359956, 42.5916678110759, 43.0333340962728, 43.3166662851969, 
    43.6999994913737, 43.9166666666667, 44.2666651407878, 44.6866663614909, 
    45.0000012715658, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3791662851969, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    39.966667175293, 40.3888884650336, 40.6666666666667, 41.006667582194, 
    41.3575752720688, 41.6444447835286, 41.9952385312035, 42.3952378772554, 
    42.5666681925456, 43.3166662851969, 43.6416670481364, 44.6999994913737, 
    44.9666675991482, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    40.4266665140788, 40.6666666666667, 40.9757580612645, 41.3380948021298, 
    41.6380956740606, 43.3166662851969, 43.6666666666667, 44.7041660944621, 
    44.9757580612645, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.657575896292, 46.9541670481364, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 44.9866671244303, 
    45.3666661580404, 45.6666666666667, 46.3666661580404, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3575752720688, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3766661326091, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.657575896292, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.9541670481364, 36.3791662851969, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6541668574015, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3266657511393, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6166674296061, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6166674296061, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.9541670481364, 33.3166662851969, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.9541670481364, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3523802984329, 32.6466669718424, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 37.5846659342448, 
    37.5846659342448, 37.5846659342448, 37.5846659342448, 37.5846659342448, 
    37.5846659342448, 37.5846659342448, 37.5846659342448, 37.5846659342448, 
    37.5846659342448, 37.5846659342448, 37.5846659342448, 37.5846659342448, 
    37.5846659342448, 37.5846659342448, 37.5846659342448, 37.5846659342448, 
    37.5846659342448, 37.5846659342448, 37.5846659342448, 37.5846659342448, 
    37.5846659342448, 37.5846659342448, 37.5846659342448, 37.5846659342448, 
    37.5846659342448, 37.5846659342448, 37.5846659342448, 37.5846659342448, 
    37.5846659342448, 37.5846659342448, 37.5846659342448, 37.5846659342448, 
    37.5846659342448, 37.5846659342448, 37.5846659342448, 37.5846659342448, 
    37.5846659342448, 38.4526659647624, 38.4526659647624, 38.4526659647624, 
    38.4526659647624, 38.4526659647624, 38.4526659647624, 38.4526659647624, 
    38.4526659647624, 38.4526659647624, 38.4526659647624, 38.4526659647624, 
    38.4526659647624, 38.4526659647624, 38.4526659647624, 38.4526659647624, 
    38.4526659647624, 38.4526659647624, 38.4526659647624, 38.4526659647624, 
    38.4526659647624, 38.4526659647624, 38.4526659647624, 38.4526659647624, 
    38.4526659647624, 38.4526659647624, 38.4526659647624, 38.4526659647624, 
    38.4526659647624, 38.4526659647624, 38.4526659647624, 38.4526659647624, 
    38.4526659647624, 38.4526659647624, 38.4526659647624, 38.4526659647624, 
    38.4526659647624, 38.4526659647624, 38.4526659647624, 38.4526659647624, 
    38.4526659647624, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3666661580404, 38.6666666666667, 38.966667175293, 
    39.3666661580404, 39.6666666666667, 39.966667175293, 40.3666661580404, 
    40.6666666666667, 40.966667175293, 41.3666661580404, 41.6666666666667, 
    41.966667175293, 42.3666661580404, 42.6666666666667, 42.966667175293, 
    43.3666661580404, 43.6666666666667, 43.966667175293, 44.3666661580404, 
    44.6666666666667, 44.966667175293, 45.3666661580404, 45.6666666666667, 
    45.966667175293, 46.3666661580404, 46.6666666666667, 46.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.966667175293, 41.3666661580404, 41.6666666666667, 41.966667175293, 
    42.3666661580404, 42.6666666666667, 42.966667175293, 43.3666661580404, 
    43.6666666666667, 43.966667175293, 44.3666661580404, 44.6666666666667, 
    44.966667175293, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    39.966667175293, 40.3666661580404, 40.6666666666667, 40.966667175293, 
    41.3666661580404, 41.6666666666667, 41.966667175293, 42.3666661580404, 
    42.6666666666667, 42.966667175293, 43.3666661580404, 43.6666666666667, 
    43.966667175293, 44.3666661580404, 44.6666666666667, 44.966667175293, 
    45.3666661580404, 45.6666666666667, 45.966667175293, 46.3666661580404, 
    46.6666666666667, 46.966667175293, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 38.3666661580404, 38.6666666666667, 
    38.966667175293, 39.3666661580404, 39.6666666666667, 39.966667175293, 
    40.3666661580404, 40.6666666666667, 40.966667175293, 41.3666661580404, 
    41.6666666666667, 41.966667175293, 42.3666661580404, 42.6666666666667, 
    42.966667175293, 43.3666661580404, 43.6666666666667, 43.966667175293, 
    44.3666661580404, 44.6666666666667, 44.966667175293, 45.3666661580404, 
    45.6666666666667, 45.966667175293, 46.3666661580404, 46.6666666666667, 
    46.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3666661580404, 38.6666666666667, 38.966667175293, 
    39.3666661580404, 39.6666666666667, 39.966667175293, 40.3666661580404, 
    40.6666666666667, 40.966667175293, 41.3666661580404, 41.6666666666667, 
    41.966667175293, 42.3666661580404, 42.6666666666667, 42.966667175293, 
    43.3666661580404, 43.6666666666667, 43.966667175293, 44.3666661580404, 
    44.6666666666667, 44.966667175293, 45.3666661580404, 45.6666666666667, 
    45.966667175293, 46.3666661580404, 46.6666666666667, 46.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.966667175293, 41.3666661580404, 41.6666666666667, 41.966667175293, 
    42.3666661580404, 42.6666666666667, 42.966667175293, 43.3666661580404, 
    43.6666666666667, 43.966667175293, 44.3666661580404, 44.6666666666667, 
    44.966667175293, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    39.966667175293, 40.3666661580404, 40.6666666666667, 40.966667175293, 
    41.3666661580404, 41.6666666666667, 41.966667175293, 42.3666661580404, 
    42.6666666666667, 42.966667175293, 43.3666661580404, 43.6666666666667, 
    43.966667175293, 44.3666661580404, 44.6666666666667, 44.966667175293, 
    45.3666661580404, 45.6666666666667, 45.966667175293, 46.3666661580404, 
    46.6666666666667, 46.966667175293, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 38.3666661580404, 38.6666666666667, 
    38.966667175293, 39.3666661580404, 39.6666666666667, 39.966667175293, 
    40.3666661580404, 40.6666666666667, 40.966667175293, 41.3666661580404, 
    41.6666666666667, 41.966667175293, 42.3666661580404, 42.6666666666667, 
    42.966667175293, 43.3666661580404, 43.6666666666667, 43.966667175293, 
    44.3666661580404, 44.6666666666667, 44.966667175293, 45.3666661580404, 
    45.6666666666667, 45.966667175293, 46.3666661580404, 46.6666666666667, 
    46.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3666661580404, 38.6666666666667, 38.966667175293, 
    39.3666661580404, 39.6666666666667, 39.966667175293, 40.3666661580404, 
    40.6666666666667, 40.966667175293, 41.3666661580404, 41.6666666666667, 
    41.966667175293, 42.3666661580404, 42.6666666666667, 42.966667175293, 
    43.3666661580404, 43.6666666666667, 43.966667175293, 44.3666661580404, 
    44.6666666666667, 44.966667175293, 45.3666661580404, 45.6666666666667, 
    45.966667175293, 46.3666661580404, 46.6666666666667, 46.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.966667175293, 41.3666661580404, 41.6666666666667, 41.966667175293, 
    42.3666661580404, 42.6666666666667, 42.966667175293, 43.3666661580404, 
    43.6666666666667, 43.966667175293, 44.3666661580404, 44.6666666666667, 
    44.966667175293, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    39.966667175293, 40.3666661580404, 40.6666666666667, 40.966667175293, 
    41.3666661580404, 41.6666666666667, 41.966667175293, 42.3666661580404, 
    42.6666666666667, 42.966667175293, 43.3666661580404, 43.6666666666667, 
    43.966667175293, 44.3666661580404, 44.6666666666667, 44.966667175293, 
    45.3666661580404, 45.6666666666667, 45.966667175293, 46.3666661580404, 
    46.6666666666667, 46.966667175293, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 38.3666661580404, 38.6666666666667, 
    38.966667175293, 39.3666661580404, 39.6666666666667, 39.966667175293, 
    40.3666661580404, 40.6666666666667, 40.966667175293, 41.3666661580404, 
    41.6666666666667, 41.966667175293, 42.3666661580404, 42.6666666666667, 
    42.966667175293, 43.3666661580404, 43.6666666666667, 43.966667175293, 
    44.3666661580404, 44.6666666666667, 44.966667175293, 45.3666661580404, 
    45.6666666666667, 45.966667175293, 46.3666661580404, 46.6666666666667, 
    46.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3666661580404, 38.6666666666667, 38.966667175293, 
    39.3666661580404, 39.6666666666667, 39.966667175293, 40.3666661580404, 
    40.6666666666667, 40.966667175293, 41.3666661580404, 41.6666666666667, 
    41.966667175293, 42.3666661580404, 42.6666666666667, 42.966667175293, 
    43.3666661580404, 43.6666666666667, 43.966667175293, 44.3666661580404, 
    44.6666666666667, 44.966667175293, 45.3666661580404, 45.6666666666667, 
    45.966667175293, 46.3666661580404, 46.6666666666667, 46.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.966667175293, 41.3666661580404, 41.6757574370413, 41.966667175293, 
    42.3523802984328, 42.5666681925456, 42.9666668574015, 43.3666659037272, 
    43.6291672388713, 43.966667175293, 44.3666661580404, 44.6809521629697, 
    44.966667175293, 45.3566660563151, 45.6666666666667, 45.9666672908899, 
    46.3866663614909, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    39.966667175293, 40.3666661580404, 40.6666666666667, 40.966667175293, 
    41.3575752720688, 41.6666666666667, 41.966667175293, 42.3666659037272, 
    42.6380956740606, 42.9666670481364, 43.3999989827474, 43.6999994913737, 
    43.9541670481364, 44.7666651407878, 44.9666675385975, 45.3666659037272, 
    45.6666666666667, 45.966667175293, 46.4000002543131, 46.6666666666667, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.9666674296061, 41.3666661580404, 41.6666666666667, 41.9333337148031, 
    42.3809518359956, 42.5916678110759, 43.0333340962728, 43.3166662851969, 
    43.6999994913737, 43.9166666666667, 44.2666651407878, 44.6866663614909, 
    45.0000012715658, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3791662851969, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    39.966667175293, 40.3888884650336, 40.6666666666667, 41.006667582194, 
    41.3575752720688, 41.6444447835286, 41.9952385312035, 42.3952378772554, 
    42.5666681925456, 43.3166662851969, 43.6416670481364, 44.6999994913737, 
    44.9666675991482, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    40.4266665140788, 40.6791664759318, 40.9757580612645, 41.3380948021298, 
    41.6380956740606, 43.3166662851969, 43.6666666666667, 44.7041660944621, 
    44.9757580612645, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.657575896292, 46.9541670481364, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 44.9866671244303, 
    45.3666661580404, 45.6666666666667, 46.3666661580404, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3575752720688, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3766661326091, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.657575896292, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.9541670481364, 36.3791662851969, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6541668574015, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3266657511393, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6166674296061, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6166674296061, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.9541670481364, 33.3166662851969, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.9541670481364, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3523802984329, 32.6466669718424, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 34.122667948405, 
    34.122667948405, 34.122667948405, 34.122667948405, 34.122667948405, 
    34.122667948405, 34.122667948405, 34.122667948405, 34.122667948405, 
    34.122667948405, 34.122667948405, 34.122667948405, 34.122667948405, 
    34.122667948405, 34.122667948405, 34.122667948405, 34.122667948405, 
    34.122667948405, 34.122667948405, 34.122667948405, 34.122667948405, 
    34.122667948405, 34.122667948405, 34.122667948405, 34.122667948405, 
    34.122667948405, 34.122667948405, 34.122667948405, 34.122667948405, 
    34.122667948405, 34.122667948405, 34.122667948405, 34.122667948405, 
    34.122667948405, 34.122667948405, 34.122667948405, 34.122667948405, 
    34.122667948405, 34.122667948405, 34.122667948405, 34.122667948405, 
    34.122667948405, 34.122667948405, 34.122667948405, 34.122667948405, 
    34.122667948405, 42.2416674296061, 42.2416674296061, 42.2416674296061, 
    42.2416674296061, 42.2416674296061, 42.2416674296061, 42.2416674296061, 
    42.2416674296061, 42.2416674296061, 42.2416674296061, 42.2416674296061, 
    42.2416674296061, 42.2416674296061, 42.2416674296061, 42.2416674296061, 
    42.2416674296061, 42.2416674296061, 42.2416674296061, 42.2416674296061, 
    42.2416674296061, 42.2416674296061, 42.2416674296061, 42.2416674296061, 
    42.2416674296061, 42.2416674296061, 42.2416674296061, 42.2416674296061, 
    42.2416674296061, 42.2416674296061, 42.2416674296061, 42.2416674296061, 
    42.2416674296061, 42.2416674296061, 42.2416674296061, 42.2416674296061, 
    42.2416674296061, 42.2416674296061, 42.2416674296061, 42.2416674296061, 
    42.2416674296061, 42.2416674296061, 42.2416674296061, 42.2416674296061, 
    42.2416674296061, 42.2416674296061, 42.2416674296061, 44.8956667582194, 
    44.8956667582194, 44.8956667582194, 44.8956667582194, 44.8956667582194, 
    44.8956667582194, 44.8956667582194, 44.8956667582194, 44.8956667582194, 
    44.8956667582194, 44.8956667582194, 44.8956667582194, 44.8956667582194, 
    44.8956667582194, 44.8956667582194, 44.8956667582194, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    39.966667175293, 40.3666661580404, 40.6666666666667, 40.966667175293, 
    41.3666661580404, 41.6666666666667, 41.966667175293, 42.3666661580404, 
    42.6666666666667, 42.966667175293, 43.3666661580404, 43.6666666666667, 
    43.966667175293, 44.3666661580404, 44.6666666666667, 44.966667175293, 
    45.3666661580404, 45.6666666666667, 45.966667175293, 46.3666661580404, 
    46.6666666666667, 46.966667175293, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 38.3666661580404, 38.6666666666667, 
    38.966667175293, 39.3666661580404, 39.6666666666667, 39.966667175293, 
    40.3666661580404, 40.6666666666667, 40.966667175293, 41.3666661580404, 
    41.6666666666667, 41.966667175293, 42.3666661580404, 42.6666666666667, 
    42.966667175293, 43.3666661580404, 43.6666666666667, 43.966667175293, 
    44.3666661580404, 44.6666666666667, 44.966667175293, 45.3666661580404, 
    45.6666666666667, 45.966667175293, 46.3666661580404, 46.6666666666667, 
    46.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3666661580404, 38.6666666666667, 38.966667175293, 
    39.3666661580404, 39.6666666666667, 39.966667175293, 40.3666661580404, 
    40.6666666666667, 40.966667175293, 41.3666661580404, 41.6666666666667, 
    41.966667175293, 42.3666661580404, 42.6666666666667, 42.966667175293, 
    43.3666661580404, 43.6666666666667, 43.966667175293, 44.3666661580404, 
    44.6666666666667, 44.966667175293, 45.3666661580404, 45.6666666666667, 
    45.966667175293, 46.3666661580404, 46.6666666666667, 46.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.966667175293, 41.3666661580404, 41.6666666666667, 41.966667175293, 
    42.3666661580404, 42.6666666666667, 42.966667175293, 43.3666661580404, 
    43.6666666666667, 43.966667175293, 44.3666661580404, 44.6666666666667, 
    44.966667175293, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    39.966667175293, 40.3666661580404, 40.6666666666667, 40.966667175293, 
    41.3666661580404, 41.6666666666667, 41.966667175293, 42.3666661580404, 
    42.6666666666667, 42.966667175293, 43.3666661580404, 43.6666666666667, 
    43.966667175293, 44.3666661580404, 44.6666666666667, 44.966667175293, 
    45.3666661580404, 45.6666666666667, 45.966667175293, 46.3666661580404, 
    46.6666666666667, 46.966667175293, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 38.3666661580404, 38.6666666666667, 
    38.966667175293, 39.3666661580404, 39.6666666666667, 39.966667175293, 
    40.3666661580404, 40.6666666666667, 40.966667175293, 41.3666661580404, 
    41.6666666666667, 41.966667175293, 42.3666661580404, 42.6666666666667, 
    42.966667175293, 43.3666661580404, 43.6666666666667, 43.966667175293, 
    44.3666661580404, 44.6666666666667, 44.966667175293, 45.3666661580404, 
    45.6666666666667, 45.966667175293, 46.3666661580404, 46.6666666666667, 
    46.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3666661580404, 38.6666666666667, 38.966667175293, 
    39.3666661580404, 39.6666666666667, 39.966667175293, 40.3666661580404, 
    40.6666666666667, 40.966667175293, 41.3666661580404, 41.6666666666667, 
    41.966667175293, 42.3666661580404, 42.6666666666667, 42.966667175293, 
    43.3666661580404, 43.6666666666667, 43.966667175293, 44.3666661580404, 
    44.6666666666667, 44.966667175293, 45.3666661580404, 45.6666666666667, 
    45.966667175293, 46.3666661580404, 46.6666666666667, 46.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.966667175293, 41.3666661580404, 41.6666666666667, 41.966667175293, 
    42.3666661580404, 42.6666666666667, 42.966667175293, 43.3666661580404, 
    43.6666666666667, 43.966667175293, 44.3666661580404, 44.6666666666667, 
    44.966667175293, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    39.966667175293, 40.3666661580404, 40.6666666666667, 40.966667175293, 
    41.3666661580404, 41.6666666666667, 41.966667175293, 42.3666661580404, 
    42.6666666666667, 42.966667175293, 43.3666661580404, 43.6666666666667, 
    43.966667175293, 44.3666661580404, 44.6666666666667, 44.966667175293, 
    45.3666661580404, 45.6666666666667, 45.966667175293, 46.3666661580404, 
    46.6666666666667, 46.966667175293, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 38.3666661580404, 38.6666666666667, 
    38.966667175293, 39.3666661580404, 39.6666666666667, 39.966667175293, 
    40.3666661580404, 40.6666666666667, 40.966667175293, 41.3666661580404, 
    41.6666666666667, 41.966667175293, 42.3666661580404, 42.6666666666667, 
    42.966667175293, 43.3666661580404, 43.6666666666667, 43.966667175293, 
    44.3666661580404, 44.6666666666667, 44.966667175293, 45.3666661580404, 
    45.6666666666667, 45.966667175293, 46.3666661580404, 46.6666666666667, 
    46.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3666661580404, 38.6666666666667, 38.966667175293, 
    39.3666661580404, 39.6666666666667, 39.966667175293, 40.3666661580404, 
    40.6666666666667, 40.966667175293, 41.3666661580404, 41.6666666666667, 
    41.966667175293, 42.3666661580404, 42.6666666666667, 42.966667175293, 
    43.3666661580404, 43.6666666666667, 43.966667175293, 44.3666661580404, 
    44.6666666666667, 44.966667175293, 45.3666661580404, 45.6666666666667, 
    45.966667175293, 46.3666661580404, 46.6666666666667, 46.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.966667175293, 41.3666661580404, 41.6666666666667, 41.966667175293, 
    42.3666661580404, 42.6666666666667, 42.966667175293, 43.3666661580404, 
    43.6666666666667, 43.966667175293, 44.3666661580404, 44.6666666666667, 
    44.966667175293, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    39.966667175293, 40.3666661580404, 40.6666666666667, 40.966667175293, 
    41.3666661580404, 41.6666666666667, 41.966667175293, 42.3666661580404, 
    42.6666666666667, 42.966667175293, 43.3666661580404, 43.6666666666667, 
    43.966667175293, 44.3666661580404, 44.6666666666667, 44.966667175293, 
    45.3666661580404, 45.6666666666667, 45.966667175293, 46.3666661580404, 
    46.6666666666667, 46.966667175293, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 38.3666661580404, 38.6666666666667, 
    38.966667175293, 39.3666661580404, 39.6666666666667, 39.966667175293, 
    40.3666661580404, 40.6666666666667, 40.966667175293, 41.3666661580404, 
    41.6888885498047, 41.966667175293, 42.2916657129923, 42.9666668574015, 
    43.2666651407878, 43.6095246814546, 43.966667175293, 44.3666661580404, 
    44.6809521629697, 44.9666674296061, 45.3666660424435, 45.6666666666667, 
    45.9666672908899, 46.3866663614909, 46.6666666666667, 46.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.966667175293, 41.3575752720688, 41.6777776082357, 41.966667175293, 
    42.3666659037272, 42.6500002543132, 42.9666670481364, 43.2666651407878, 
    43.6166674296061, 43.9541670481364, 44.7666651407878, 44.9666678110758, 
    45.3666659037272, 45.6666666666667, 45.966667175293, 46.4000002543131, 
    46.6666666666667, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3666661580404, 38.6666666666667, 38.966667175293, 
    39.3666661580404, 39.6666666666667, 39.966667175293, 40.3666661580404, 
    40.6666666666667, 40.9416672388713, 41.3666655222575, 41.6999994913737, 
    41.9000002543132, 42.3809518359956, 42.5916678110759, 43.0333340962728, 
    43.3666674296061, 43.6866663614909, 43.9166666666667, 44.2666651407878, 
    44.7666651407878, 45.0000012715658, 45.3666661580404, 45.6666666666667, 
    45.966667175293, 46.3666661580404, 46.6666666666667, 46.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.9575761737245, 40.3888884650336, 40.6566668192546, 
    40.8666674296061, 41.3466654459635, 41.5666681925456, 42.3916670481364, 
    42.5666681925456, 43.3166662851969, 43.7166659037272, 44.7166659037272, 
    44.9666675991482, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    40.4266665140788, 40.6791664759318, 40.966667175293, 41.6666666666667, 
    43.7166659037272, 44.7041660944621, 44.9757580612645, 45.3666661580404, 
    45.6666666666667, 45.966667175293, 46.3666661580404, 46.657575896292, 
    46.9541670481364, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3666661580404, 38.6666666666667, 38.966667175293, 
    39.3666661580404, 44.9866671244303, 45.3666661580404, 45.6666666666667, 
    46.3666661580404, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3575752720688, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3766661326091, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.657575896292, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.9541670481364, 
    36.3791662851969, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6541668574015, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3266657511393, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6166674296061, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6166674296061, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.9541670481364, 33.3166662851969, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.9541670481364, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3523802984329, 32.6466669718424, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 41.2626673380534, 41.2626673380534, 41.2626673380534, 
    41.2626673380534, 41.2626673380534, 41.2626673380534, 41.2626673380534, 
    41.2626673380534, 41.2626673380534, 41.2626673380534, 41.2626673380534, 
    41.2626673380534, 41.2626673380534, 40.8836657206217, 40.8836657206217, 
    40.8836657206217, 40.8836657206217, 40.8836657206217, 40.8836657206217, 
    40.8836657206217, 40.8836657206217, 40.8836657206217, 40.8836657206217, 
    40.8836657206217, 40.8836657206217, 40.8836657206217, 40.8836657206217, 
    32.6146685282389, 32.6146685282389, 32.6146685282389, 32.6146685282389, 
    32.6146685282389, 32.6146685282389, 32.6146685282389, 32.6146685282389, 
    32.6146685282389, 32.6146685282389, 32.6146685282389, 32.6146685282389, 
    32.6146685282389, 32.6146685282389, 32.5836664835612, 32.5836664835612, 
    32.5836664835612, 32.5836664835612, 32.5836664835612, 32.5836664835612, 
    32.5836664835612, 32.5836664835612, 32.5836664835612, 32.5836664835612, 
    32.5836664835612, 32.5836664835612, 32.5836664835612, 32.5836664835612, 
    32.5836664835612, 32.5836664835612, 32.5836664835612, 32.5836664835612, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.966667175293, 41.3666661580404, 41.6666666666667, 41.966667175293, 
    42.3666661580404, 42.6666666666667, 42.966667175293, 43.3666661580404, 
    43.6666666666667, 43.966667175293, 44.3666661580404, 44.6666666666667, 
    44.966667175293, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    39.966667175293, 40.3666661580404, 40.6666666666667, 40.966667175293, 
    41.3666661580404, 41.6666666666667, 41.966667175293, 42.3666661580404, 
    42.6666666666667, 42.966667175293, 43.3666661580404, 43.6666666666667, 
    43.966667175293, 44.3666661580404, 44.6666666666667, 44.966667175293, 
    45.3666661580404, 45.6666666666667, 45.966667175293, 46.3666661580404, 
    46.6666666666667, 46.966667175293, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 38.3666661580404, 38.6666666666667, 
    38.966667175293, 39.3666661580404, 39.6666666666667, 39.966667175293, 
    40.3666661580404, 40.6666666666667, 40.966667175293, 41.3666661580404, 
    41.6666666666667, 41.966667175293, 42.3666661580404, 42.6666666666667, 
    42.966667175293, 43.3666661580404, 43.6666666666667, 43.966667175293, 
    44.3666661580404, 44.6666666666667, 44.966667175293, 45.3666661580404, 
    45.6666666666667, 45.966667175293, 46.3666661580404, 46.6666666666667, 
    46.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3666661580404, 38.6666666666667, 38.966667175293, 
    39.3666661580404, 39.6666666666667, 39.966667175293, 40.3666661580404, 
    40.6666666666667, 40.966667175293, 41.3666661580404, 41.6666666666667, 
    41.966667175293, 42.3666661580404, 42.6666666666667, 42.966667175293, 
    43.3666661580404, 43.6666666666667, 43.966667175293, 44.3666661580404, 
    44.6666666666667, 44.966667175293, 45.3666661580404, 45.6666666666667, 
    45.966667175293, 46.3666661580404, 46.6666666666667, 46.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.966667175293, 41.3666661580404, 41.6666666666667, 41.966667175293, 
    42.3666661580404, 42.6666666666667, 42.966667175293, 43.3666661580404, 
    43.6666666666667, 43.966667175293, 44.3666661580404, 44.6666666666667, 
    44.966667175293, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    39.966667175293, 40.3666661580404, 40.6666666666667, 40.966667175293, 
    41.3666661580404, 41.6666666666667, 41.966667175293, 42.3666661580404, 
    42.6666666666667, 42.966667175293, 43.3666661580404, 43.6666666666667, 
    43.966667175293, 44.3666661580404, 44.6666666666667, 44.966667175293, 
    45.3666661580404, 45.6666666666667, 45.966667175293, 46.3666661580404, 
    46.6666666666667, 46.966667175293, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 38.3666661580404, 38.6666666666667, 
    38.966667175293, 39.3666661580404, 39.6666666666667, 39.966667175293, 
    40.3666661580404, 40.6666666666667, 40.966667175293, 41.3666661580404, 
    41.6666666666667, 41.966667175293, 42.3666661580404, 42.6666666666667, 
    42.966667175293, 43.3666661580404, 43.6666666666667, 43.966667175293, 
    44.3666661580404, 44.6666666666667, 44.966667175293, 45.3666661580404, 
    45.6666666666667, 45.966667175293, 46.3666661580404, 46.6666666666667, 
    46.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3666661580404, 38.6666666666667, 38.966667175293, 
    39.3666661580404, 39.6666666666667, 39.966667175293, 40.3666661580404, 
    40.6666666666667, 40.966667175293, 41.3666661580404, 41.6666666666667, 
    41.966667175293, 42.3666661580404, 42.6666666666667, 42.966667175293, 
    43.3666661580404, 43.6666666666667, 43.966667175293, 44.3666661580404, 
    44.6666666666667, 44.966667175293, 45.3666661580404, 45.6666666666667, 
    45.966667175293, 46.3666661580404, 46.6666666666667, 46.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.966667175293, 41.3666661580404, 41.6666666666667, 41.966667175293, 
    42.3666661580404, 42.6666666666667, 42.966667175293, 43.3666661580404, 
    43.6666666666667, 43.966667175293, 44.3666661580404, 44.6666666666667, 
    44.966667175293, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666661580404, 39.6666666666667, 
    39.966667175293, 40.3666661580404, 40.6666666666667, 40.966667175293, 
    41.3666661580404, 41.6666666666667, 41.966667175293, 42.3666661580404, 
    42.6666666666667, 42.966667175293, 43.3666661580404, 43.6666666666667, 
    43.966667175293, 44.3666661580404, 44.6666666666667, 44.966667175293, 
    45.3666661580404, 45.6666666666667, 45.966667175293, 46.3666661580404, 
    46.6666666666667, 46.966667175293, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 38.3666661580404, 38.6666666666667, 
    38.966667175293, 39.3666661580404, 39.6666666666667, 39.966667175293, 
    40.3666661580404, 40.6666666666667, 40.966667175293, 41.3666661580404, 
    41.6666666666667, 41.966667175293, 42.3666661580404, 42.6666666666667, 
    42.966667175293, 43.3666661580404, 43.6666666666667, 43.966667175293, 
    44.3666661580404, 44.6666666666667, 44.966667175293, 45.3666661580404, 
    45.6666666666667, 45.966667175293, 46.3666661580404, 46.6666666666667, 
    46.966667175293, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3666661580404, 38.6666666666667, 38.966667175293, 
    39.3666661580404, 39.6666666666667, 39.966667175293, 40.3666661580404, 
    40.6666666666667, 40.966667175293, 41.3666661580404, 41.6666666666667, 
    41.966667175293, 42.3666661580404, 42.6666666666667, 42.966667175293, 
    43.3666661580404, 43.6666666666667, 43.966667175293, 44.3666661580404, 
    44.6666666666667, 44.966667175293, 45.3666661580404, 45.6666666666667, 
    45.966667175293, 46.3666661580404, 46.6666666666667, 46.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.966667175293, 39.3666661580404, 
    39.6666666666667, 39.966667175293, 40.3666661580404, 40.6666666666667, 
    40.966667175293, 41.3666661580404, 41.6666666666667, 41.966667175293, 
    42.3666661580404, 42.6666666666667, 42.966667175293, 43.3666661580404, 
    43.6666666666667, 43.966667175293, 44.3666661580404, 44.6666666666667, 
    44.966667175293, 45.3666661580404, 45.6666666666667, 45.966667175293, 
    46.3666661580404, 46.6666666666667, 46.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 38.3666661580404, 
    38.6666666666667, 38.966667175293, 39.3666660424435, 39.6666666666667, 
    39.9575761737245, 40.3666661580404, 40.6666666666667, 40.966667175293, 
    41.3575752720688, 41.6809521629697, 41.9541670481364, 42.3666674296061, 
    43.966667175293, 44.3666662851969, 44.6791664759318, 44.955556233724, 
    45.3666660424435, 45.6666666666667, 45.966667175293, 46.3666661580404, 
    46.6666666666667, 46.966667175293, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 38.3666661580404, 38.6666666666667, 
    38.966667175293, 39.3666660424435, 39.6666666666667, 39.966667175293, 
    40.3666660424435, 40.6266672770182, 41.0095245724633, 41.3291660944621, 
    41.6999994913737, 41.9333335028754, 42.3166662851969, 44.3916670481364, 
    44.7166659037272, 44.916667620341, 45.3766661326091, 45.6666666666667, 
    45.966667175293, 46.3666661580403, 46.6666666666667, 46.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    34.3666661580404, 34.6666666666667, 34.966667175293, 35.3666661580404, 
    35.6666666666667, 35.966667175293, 36.3666661580404, 36.6666666666667, 
    36.966667175293, 37.3666661580404, 37.6666666666667, 37.966667175293, 
    38.3666661580404, 38.6666666666667, 38.9541670481364, 39.3541661898295, 
    39.6666666666667, 39.9523814973377, 40.3266657511393, 41.2666651407878, 
    41.7666651407878, 44.7166659037272, 45.0000006357829, 45.3666661580404, 
    45.6666666666667, 45.966667175293, 46.3666661580404, 46.6666666666667, 
    46.9541670481364, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 37.6666666666667, 
    37.966667175293, 38.3666661580404, 38.6666666666667, 38.966667175293, 
    39.3575752720688, 39.657575896292, 40.4041663805644, 40.6566668192546, 
    40.8666674296061, 42.5666681925456, 44.7166659037272, 44.9666674296061, 
    45.3666661580404, 45.6666666666667, 45.966667175293, 46.3666661580404, 
    46.6666666666667, 46.966667175293, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 38.3666661580404, 38.6666666666667, 
    38.966667175293, 39.3666661580404, 39.6380956740606, 40.4266665140788, 
    40.6666666666667, 40.8666674296061, 44.7041660944621, 44.9757580612645, 
    45.3666661580404, 45.6666666666667, 45.966667175293, 46.3666661580404, 
    46.657575896292, 46.9541670481364, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 38.3666661580404, 38.6666666666667, 
    38.966667175293, 39.3666661580404, 44.9866671244303, 45.3666661580404, 
    45.6666666666667, 46.3666661580404, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6666666666667, 35.966667175293, 
    36.3666661580404, 36.6666666666667, 36.966667175293, 37.3666661580404, 
    37.6666666666667, 37.966667175293, 38.3575752720688, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 37.6666666666667, 37.966667175293, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.6666666666667, 36.966667175293, 
    37.3666661580404, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.966667175293, 33.3666661580404, 33.6666666666667, 
    33.966667175293, 34.3666661580404, 34.6666666666667, 34.966667175293, 
    35.3666661580404, 35.6666666666667, 35.966667175293, 36.3666661580404, 
    36.6666666666667, 36.966667175293, 37.3666661580404, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.966667175293, 36.3666661580404, 36.657575896292, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3666661580404, 35.6666666666667, 
    35.9541670481364, 36.3791662851969, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    34.966667175293, 35.3666661580404, 35.6541668574015, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 35.3266657511393, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6666666666667, 33.966667175293, 34.3666661580404, 
    34.6666666666667, 34.966667175293, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6666666666667, 33.966667175293, 34.3666661580404, 34.6666666666667, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 33.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.966667175293, 33.3666661580404, 33.6666666666667, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    33.3666661580404, 33.6166674296061, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 31.6666660308838, 31.966667175293, 
    32.3666661580404, 32.6666666666667, 32.966667175293, 33.3666661580404, 
    33.6166674296061, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3666661580404, 
    32.6666666666667, 32.9541670481364, 33.3166662851969, 30.3666667938232, 
    30.6666666666667, 30.9666665395101, 31.3666667938232, 31.6666660308838, 
    31.966667175293, 32.3666661580404, 32.6666666666667, 32.966667175293, 
    30.3666667938232, 30.6666666666667, 30.9666665395101, 31.3666667938232, 
    31.6666660308838, 31.966667175293, 32.3666661580404, 32.6666666666667, 
    32.9541670481364, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 31.966667175293, 32.3523802984329, 
    32.6466669718424, 30.3666667938232, 30.6666666666667, 30.9666665395101, 
    31.3666667938232, 31.6666660308838, 30.3666667938232, 30.6666666666667, 
    30.9666665395101, 31.3666667938232, 32.3496653238932, 32.3496653238932, 
    32.3496653238932, 32.3496653238932, 32.3496653238932, 32.3496653238932, 
    32.3496653238932, 32.3496653238932, 32.3496653238932, 32.3496653238932, 
    32.3496653238932, 32.3496653238932, 32.3496653238932, 32.3496653238932, 
    32.3496653238932, 32.3496653238932, 32.3496653238932, 32.3496653238932, 
    32.013666788737, 32.013666788737, 32.013666788737, 32.013666788737, 
    32.013666788737, 32.013666788737, 32.013666788737, 32.013666788737, 
    32.013666788737, 32.013666788737, 32.013666788737, 32.013666788737, 
    32.013666788737, 32.013666788737, 32.013666788737, 32.013666788737, 
    32.013666788737, 32.013666788737, 32.013666788737, 32.013666788737, 
    32.013666788737, 32.013666788737, 32.013666788737, 32.013666788737, 
    32.013666788737, 32.013666788737, 32.013666788737, 32.013666788737, 
    32.013666788737, 32.013666788737, 30.6170631237561, 30.6170631237561, 
    30.9025056550392, 30.6170631237561, 30.9025056550392, 30.6170631237561, 
    30.9025056550392, 30.6170631237561, 30.9025056550392, 31.7536566677173, 
    30.6170631237561, 30.9025056550392, 31.7536566677173, 30.6170631237561, 
    32.0356337743697, 30.9025056550392, 31.7536566677173, 30.6170631237561, 
    32.0356337743697, 30.9025056550392, 31.7536566677173, 32.3167339917995, 
    30.6170631237561, 32.0356337743697, 30.9025056550392, 31.7536566677173, 
    32.3167339917995, 30.6170631237561, 32.0356337743697, 32.5969533019733, 
    30.9025056550392, 31.7536566677173, 32.3167339917995, 30.6170631237561, 
    32.0356337743697, 32.5969533019733, 30.9025056550392, 31.7536566677173, 
    32.3167339917995, 30.6170631237561, 32.8762877838633, 32.0356337743697, 
    32.5969533019733, 30.9025056550392, 31.7536566677173, 32.3167339917995, 
    30.6170631237561, 32.8762877838633, 32.0356337743697, 32.5969533019733, 
    30.9025056550392, 33.432287061478, 31.7536566677173, 32.3167339917995, 
    30.6170631237561, 32.8762877838633, 32.0356337743697, 32.5969533019733, 
    30.9025056550392, 33.432287061478, 31.7536566677173, 32.3167339917995, 
    30.6170631237561, 32.8762877838633, 33.7089444967663, 32.0356337743697, 
    32.5969533019733, 30.9025056550392, 33.432287061478, 31.7536566677173, 
    32.3167339917995, 30.6170631237561, 32.8762877838633, 33.7089444967663, 
    32.0356337743697, 32.5969533019733, 30.9025056550392, 33.432287061478, 
    31.7536566677173, 33.9847023820702, 32.3167339917995, 30.6170631237561, 
    32.8762877838633, 33.7089444967663, 32.0356337743697, 32.5969533019733, 
    30.9025056550392, 33.432287061478, 31.7536566677173, 33.9847023820702, 
    32.3167339917995, 30.6170631237561, 32.8762877838633, 33.7089444967663, 
    32.0356337743697, 34.2595572754987, 32.5969533019733, 30.9025056550392, 
    33.432287061478, 31.7536566677173, 33.9847023820702, 32.3167339917995, 
    30.6170631237561, 32.8762877838633, 33.7089444967663, 32.0356337743697, 
    34.2595572754987, 32.5969533019733, 30.9025056550392, 33.432287061478, 
    31.7536566677173, 33.9847023820702, 32.3167339917995, 30.6170631237561, 
    34.5335058296867, 32.8762877838633, 33.7089444967663, 32.0356337743697, 
    34.2595572754987, 32.5969533019733, 30.9025056550392, 33.432287061478, 
    31.7536566677173, 33.9847023820702, 32.3167339917995, 30.6170631237561, 
    34.5335058296867, 32.8762877838633, 33.7089444967663, 32.0356337743697, 
    34.2595572754987, 32.5969533019733, 30.9025056550392, 35.0786710006513, 
    33.432287061478, 31.7536566677173, 33.9847023820702, 32.3167339917995, 
    30.6170631237561, 34.5335058296867, 32.8762877838633, 33.7089444967663, 
    32.0356337743697, 34.2595572754987, 32.5969533019733, 30.9025056550392, 
    35.0786710006513, 33.432287061478, 31.7536566677173, 33.9847023820702, 
    32.3167339917995, 30.6170631237561, 34.5335058296867, 32.8762877838633, 
    35.3498813909852, 33.7089444967663, 32.0356337743697, 34.2595572754987, 
    32.5969533019733, 30.9025056550392, 35.0786710006513, 33.432287061478, 
    31.7536566677173, 33.9847023820702, 32.3167339917995, 30.6170631237561, 
    34.5335058296867, 32.8762877838633, 35.3498813909852, 33.7089444967663, 
    32.0356337743697, 34.2595572754987, 32.5969533019733, 30.9025056550392, 
    35.0786710006513, 33.432287061478, 31.7536566677173, 35.620172988168, 
    33.9847023820702, 32.3167339917995, 30.6170631237561, 34.5335058296867, 
    32.8762877838633, 35.3498813909853, 33.7089444967663, 32.0356337743697, 
    34.2595572754987, 32.5969533019733, 30.9025056550392, 35.0786710006513, 
    33.432287061478, 31.7536566677173, 35.620172988168, 33.9847023820702, 
    32.3167339917995, 30.6170631237561, 34.5335058296867, 32.8762877838633, 
    35.3498813909852, 33.7089444967663, 32.0356337743697, 35.8895429100474, 
    34.2595572754987, 32.5969533019733, 30.9025056550392, 35.0786710006513, 
    33.432287061478, 31.7536566677173, 35.620172988168, 33.9847023820702, 
    32.3167339917995, 30.6170631237561, 34.5335058296867, 32.8762877838633, 
    35.3498813909852, 33.7089444967663, 32.0356337743697, 35.8895429100474, 
    34.2595572754987, 32.5969533019733, 30.9025056550392, 35.0786710006513, 
    33.432287061478, 31.7536566677173, 35.620172988168, 33.9847023820702, 
    32.3167339917995, 36.4255066559906, 30.6170631237561, 34.5335058296867, 
    32.8762877838633, 35.3498813909852, 33.7089444967663, 32.0356337743697, 
    35.8895429100474, 34.2595572754987, 32.5969533019733, 30.9025056550392, 
    35.0786710006513, 33.432287061478, 31.7536566677173, 35.620172988168, 
    33.9847023820702, 32.3167339917995, 36.4255066559906, 30.6170631237561, 
    34.5335058296867, 32.8762877838633, 35.3498813909852, 33.7089444967663, 
    32.0356337743697, 35.8895429100474, 34.2595572754987, 32.5969533019733, 
    36.6920951707497, 30.9025056550392, 35.0786710006513, 33.432287061478, 
    31.7536566677173, 35.620172988168, 33.9847023820702, 32.3167339917995, 
    36.4255066559906, 30.6170631237561, 34.5335058296867, 32.8762877838633, 
    35.3498813909852, 33.7089444967663, 32.0356337743697, 35.8895429100474, 
    34.2595572754987, 32.5969533019733, 36.6920951707497, 30.9025056550392, 
    35.0786710006513, 33.432287061478, 31.7536566677173, 35.620172988168, 
    33.9847023820702, 32.3167339917995, 36.4255066559906, 30.6170631237561, 
    34.5335058296867, 32.8762877838633, 36.9577513904295, 35.3498813909852, 
    33.7089444967663, 32.0356337743697, 35.8895429100474, 34.2595572754987, 
    32.5969533019733, 36.6920951707497, 30.9025056550392, 35.0786710006513, 
    33.432287061478, 31.7536566677173, 35.620172988168, 33.9847023820702, 
    32.3167339917995, 36.4255066559906, 30.6170631237561, 34.5335058296867, 
    32.8762877838633, 36.9577513904295, 35.3498813909852, 33.7089444967663, 
    32.0356337743697, 35.8895429100474, 34.2595572754987, 32.5969533019733, 
    36.6920951707497, 30.9025056550392, 35.0786710006513, 33.432287061478, 
    37.2224728843778, 31.7536566677173, 35.620172988168, 33.9847023820702, 
    32.3167339917995, 36.4255066559906, 30.6170631237561, 34.5335058296867, 
    32.8762877838633, 36.9577513904295, 35.3498813909853, 33.7089444967663, 
    32.0356337743697, 35.8895429100474, 34.2595572754987, 32.5969533019733, 
    36.6920951707497, 30.9025056550392, 35.0786710006513, 33.432287061478, 
    37.2224728843778, 31.7536566677173, 35.620172988168, 33.9847023820702, 
    32.3167339917995, 36.4255066559906, 30.6170631237561, 34.5335058296867, 
    32.8762877838633, 36.9577513904295, 35.3498813909852, 33.7089444967663, 
    37.7491024143739, 32.0356337743697, 35.8895429100474, 34.2595572754987, 
    32.5969533019733, 36.6920951707497, 30.9025056550392, 35.0786710006513, 
    33.432287061478, 37.2224728843778, 31.7536566677173, 35.620172988168, 
    33.9847023820702, 32.3167339917995, 36.4255066559906, 30.6170631237561, 
    34.5335058296867, 32.8762877838633, 36.9577513904295, 35.3498813909852, 
    33.7089444967663, 37.749102414374, 32.0356337743697, 35.8895429100474, 
    34.2595572754987, 32.5969533019733, 36.6920951707497, 30.9025056550392, 
    35.0786710006513, 33.432287061478, 37.2224728843778, 31.7536566677173, 
    35.620172988168, 33.9847023820702, 38.0110060291271, 32.3167339917995, 
    36.4255066559906, 30.6170631237561, 34.5335058296867, 32.8762877838633, 
    36.9577513904295, 35.3498813909852, 33.7089444967663, 37.7491024143739, 
    32.0356337743697, 35.8895429100474, 34.2595572754987, 32.5969533019733, 
    36.6920951707497, 30.9025056550392, 35.0786710006513, 33.432287061478, 
    37.2224728843778, 31.7536566677173, 35.620172988168, 33.9847023820702, 
    38.0110060291271, 32.3167339917995, 36.4255066559906, 30.6170631237561, 
    34.5335058296867, 32.8762877838633, 36.9577513904295, 35.3498813909852, 
    33.7089444967663, 37.7491024143739, 32.0356337743697, 35.8895429100474, 
    34.2595572754987, 38.2719660742721, 32.5969533019733, 36.6920951707497, 
    30.9025056550392, 35.0786710006513, 33.432287061478, 37.2224728843778, 
    31.7536566677173, 35.620172988168, 33.9847023820702, 38.0110060291271, 
    32.3167339917995, 36.4255066559906, 30.6170631237561, 34.5335058296867, 
    32.8762877838633, 36.9577513904295, 35.3498813909852, 33.7089444967663, 
    37.7491024143739, 32.0356337743697, 35.8895429100474, 34.2595572754987, 
    38.2719660742721, 32.5969533019733, 36.6920951707497, 30.9025056550392, 
    35.0786710006513, 33.432287061478, 37.2224728843778, 31.7536566677173, 
    35.620172988168, 33.9847023820702, 38.0110060291271, 32.3167339917995, 
    36.4255066559906, 30.6170631237561, 34.5335058296867, 38.6615140591414, 
    32.8762877838633, 36.9577513904295, 35.3498813909852, 33.7089444967663, 
    37.7491024143739, 32.0356337743697, 35.8895429100474, 34.2595572754987, 
    38.2719660742721, 32.5969533019733, 36.6920951707497, 30.9025056550392, 
    35.0786710006513, 33.432287061478, 37.2224728843778, 31.7536566677173, 
    35.620172988168, 33.9847023820702, 38.0110060291271, 32.3167339917995, 
    36.4255066559906, 30.6170631237561, 34.5335058296867, 38.6615140591413, 
    32.8762877838633, 36.9577513904295, 35.3498813909852, 33.7089444967663, 
    37.7491024143739, 32.0356337743697, 35.8895429100474, 34.2595572754987, 
    38.2719660742721, 32.5969533019733, 36.6920951707497, 30.9025056550392, 
    35.0786710006513, 39.049165272633, 33.432287061478, 37.2224728843778, 
    31.7536566677173, 35.620172988168, 33.9847023820702, 38.0110060291271, 
    32.3167339917995, 36.4255066559906, 30.6170631237561, 34.5335058296867, 
    38.6615140591414, 32.8762877838633, 36.9577513904295, 35.3498813909852, 
    33.7089444967663, 37.7491024143739, 32.0356337743697, 35.8895429100474, 
    34.2595572754987, 38.2719660742721, 32.5969533019733, 36.6920951707497, 
    30.9025056550392, 35.0786710006513, 39.049165272633, 33.432287061478, 
    37.2224728843778, 31.7536566677173, 35.620172988168, 33.9847023820702, 
    38.0110060291271, 32.3167339917995, 36.4255066559906, 30.6170631237561, 
    34.5335058296867, 38.6615140591414, 32.8762877838633, 36.9577513904295, 
    35.3498813909853, 39.3063319434942, 33.7089444967663, 37.7491024143739, 
    32.0356337743697, 35.8895429100474, 34.2595572754987, 38.2719660742721, 
    32.5969533019733, 36.6920951707497, 30.9025056550392, 35.0786710006513, 
    39.049165272633, 33.432287061478, 37.2224728843778, 31.7536566677173, 
    35.620172988168, 33.9847023820702, 38.0110060291271, 32.3167339917995, 
    36.4255066559906, 30.6170631237561, 34.5335058296867, 38.6615140591414, 
    32.8762877838633, 36.9577513904295, 35.3498813909852, 39.3063319434942, 
    33.7089444967663, 37.7491024143739, 32.0356337743697, 35.8895429100474, 
    34.2595572754987, 38.2719660742721, 32.5969533019733, 36.6920951707497, 
    30.9025056550392, 35.0786710006513, 39.049165272633, 33.432287061478, 
    37.2224728843778, 31.7536566677173, 35.620172988168, 39.5625459179821, 
    33.9847023820702, 38.0110060291271, 32.3167339917995, 36.4255066559906, 
    30.6170631237561, 34.5335058296867, 38.6615140591414, 32.8762877838633, 
    36.9577513904295, 35.3498813909852, 39.3063319434942, 33.7089444967663, 
    37.7491024143739, 32.0356337743697, 35.8895429100474, 34.2595572754987, 
    38.2719660742721, 32.5969533019733, 36.6920951707497, 30.9025056550392, 
    35.0786710006513, 39.049165272633, 33.432287061478, 37.2224728843778, 
    31.7536566677173, 35.620172988168, 39.5625459179821, 33.9847023820702, 
    38.0110060291271, 32.3167339917995, 36.4255066559906, 30.6170631237561, 
    34.5335058296867, 38.6615140591414, 32.8762877838633, 36.9577513904295, 
    35.3498813909853, 39.3063319434942, 33.7089444967663, 37.7491024143739, 
    32.0356337743697, 35.8895429100474, 40.0721095592252, 34.2595572754987, 
    38.2719660742721, 32.5969533019733, 36.6920951707497, 30.9025056550392, 
    35.0786710006513, 39.049165272633, 33.432287061478, 37.2224728843778, 
    31.7536566677173, 35.620172988168, 39.5625459179821, 33.9847023820702, 
    38.0110060291271, 32.3167339917995, 36.4255066559906, 30.6170631237561, 
    34.5335058296867, 38.6615140591414, 32.8762877838633, 36.9577513904295, 
    35.3498813909852, 39.3063319434942, 33.7089444967663, 37.749102414374, 
    32.0356337743697, 35.8895429100474, 40.0721095592252, 34.2595572754987, 
    38.2719660742721, 32.5969533019733, 36.6920951707497, 30.9025056550392, 
    35.0786710006513, 39.049165272633, 33.432287061478, 37.2224728843778, 
    31.7536566677173, 35.620172988168, 39.5625459179821, 33.9847023820702, 
    38.0110060291271, 32.3167339917995, 36.4255066559906, 40.3254563203728, 
    30.6170631237561, 34.5335058296867, 38.6615140591414, 32.8762877838633, 
    36.9577513904295, 35.3498813909852, 39.3063319434942, 33.7089444967663, 
    37.7491024143739, 32.0356337743697, 35.8895429100474, 40.0721095592252, 
    34.2595572754987, 38.2719660742721, 32.5969533019733, 36.6920951707497, 
    30.9025056550392, 35.0786710006513, 39.049165272633, 33.432287061478, 
    37.2224728843778, 31.7536566677173, 35.620172988168, 39.5625459179821, 
    33.9847023820702, 38.0110060291271, 32.3167339917995, 36.4255066559906, 
    40.3254563203728, 30.6170631237561, 34.5335058296867, 38.6615140591413, 
    32.8762877838633, 36.9577513904295, 35.3498813909852, 39.3063319434942, 
    33.7089444967663, 37.7491024143739, 32.0356337743697, 35.8895429100474, 
    40.0721095592252, 34.2595572754987, 38.2719660742721, 32.5969533019733, 
    36.6920951707497, 40.5778445724771, 30.9025056550392, 35.0786710006513, 
    39.049165272633, 33.432287061478, 37.2224728843778, 31.7536566677173, 
    35.620172988168, 39.5625459179821, 33.9847023820702, 38.0110060291271, 
    32.3167339917995, 36.4255066559906, 40.3254563203728, 30.6170631237561, 
    34.5335058296867, 38.6615140591414, 32.8762877838633, 36.9577513904294, 
    35.3498813909852, 39.3063319434942, 33.7089444967663, 37.7491024143739, 
    32.0356337743697, 35.8895429100474, 40.0721095592252, 34.2595572754987, 
    38.2719660742721, 32.5969533019733, 36.6920951707497, 40.5778445724771, 
    30.9025056550392, 35.0786710006513, 39.049165272633, 33.432287061478, 
    37.2224728843778, 31.7536566677173, 35.620172988168, 39.5625459179821, 
    33.9847023820702, 38.0110060291271, 32.3167339917995, 36.4255066559906, 
    40.3254563203728, 30.6170631237561, 34.5335058296867, 38.6615140591414, 
    32.8762877838633, 36.9577513904295, 41.0797406188206, 35.3498813909852, 
    39.3063319434942, 33.7089444967663, 37.7491024143739, 32.0356337743697, 
    35.8895429100474, 40.0721095592252, 34.2595572754987, 38.2719660742721, 
    32.5969533019733, 36.6920951707497, 40.5778445724771, 30.9025056550392, 
    35.0786710006513, 39.049165272633, 33.432287061478, 37.2224728843778, 
    31.7536566677173, 35.620172988168, 39.5625459179821, 33.9847023820702, 
    38.0110060291271, 32.3167339917995, 36.4255066559906, 40.3254563203728, 
    34.5335058296867, 38.6615140591414, 32.8762877838633, 36.9577513904295, 
    41.0797406188206, 35.3498813909852, 39.3063319434942, 33.7089444967663, 
    37.7491024143739, 32.0356337743697, 35.8895429100474, 40.0721095592252, 
    34.2595572754987, 38.2719660742721, 32.5969533019733, 36.6920951707497, 
    40.5778445724771, 30.9025056550392, 35.0786710006513, 39.049165272633, 
    33.432287061478, 37.2224728843778, 41.3292461440167, 31.7536566677173, 
    35.620172988168, 39.5625459179821, 33.9847023820702, 38.0110060291271, 
    32.3167339917995, 36.4255066559906, 40.3254563203728, 34.5335058296867, 
    38.6615140591414, 32.8762877838633, 36.9577513904295, 41.0797406188206, 
    35.3498813909852, 39.3063319434942, 33.7089444967663, 37.7491024143739, 
    32.0356337743697, 35.8895429100474, 40.0721095592252, 34.2595572754987, 
    38.2719660742721, 32.5969533019733, 36.6920951707497, 40.5778445724771, 
    35.0786710006513, 39.049165272633, 33.432287061478, 37.2224728843778, 
    41.3292461440167, 31.7536566677173, 35.620172988168, 39.5625459179821, 
    33.9847023820702, 38.0110060291271, 32.3167339917995, 36.4255066559906, 
    40.3254563203728, 34.5335058296867, 38.6615140591413, 32.8762877838633, 
    36.9577513904295, 41.0797406188206, 35.3498813909852, 39.3063319434942, 
    33.7089444967663, 37.7491024143739, 41.5777886205734, 32.0356337743697, 
    35.8895429100474, 40.0721095592252, 34.2595572754987, 38.2719660742721, 
    32.5969533019733, 36.6920951707497, 40.5778445724771, 35.0786710006513, 
    39.049165272633, 33.432287061478, 37.2224728843778, 41.3292461440167, 
    31.7536566677173, 35.620172988168, 39.5625459179821, 33.9847023820702, 
    38.0110060291271, 32.3167339917995, 36.4255066559906, 40.3254563203728, 
    34.5335058296867, 38.6615140591414, 32.8762877838633, 36.9577513904295, 
    41.0797406188206, 35.3498813909852, 39.3063319434942, 33.7089444967663, 
    37.7491024143739, 41.5777886205734, 32.0356337743697, 35.8895429100474, 
    40.0721095592252, 34.2595572754987, 38.2719660742721, 32.5969533019733, 
    36.6920951707497, 40.5778445724771, 35.0786710006513, 39.049165272633, 
    33.432287061478, 37.2224728843778, 41.3292461440167, 35.620172988168, 
    39.5625459179821, 33.9847023820702, 38.0110060291271, 42.0719807371405, 
    32.3167339917995, 36.4255066559906, 40.3254563203728, 34.5335058296867, 
    38.6615140591414, 32.8762877838633, 36.9577513904295, 41.0797406188206, 
    35.3498813909852, 39.3063319434942, 33.7089444967663, 37.7491024143739, 
    41.5777886205734, 35.8895429100474, 40.0721095592252, 34.2595572754987, 
    38.2719660742721, 36.6920951707497, 40.5778445724771, 35.0786710006513, 
    39.049165272633, 33.432287061478, 37.2224728843778, 41.3292461440167, 
    35.620172988168, 39.5625459179821, 33.9847023820702, 38.0110060291271, 
    42.0719807371405, 32.3167339917995, 36.4255066559906, 40.3254563203728, 
    34.5335058296867, 38.6615140591413, 32.8762877838633, 36.9577513904295, 
    41.0797406188206, 35.3498813909852, 39.3063319434942, 37.749102414374, 
    41.5777886205734, 35.8895429100474, 40.0721095592252, 38.2719660742721, 
    42.3176287205335, 36.6920951707497, 40.5778445724771, 35.0786710006513, 
    39.049165272633, 33.432287061478, 37.2224728843778, 41.3292461440167, 
    35.620172988168, 39.5625459179821, 33.9847023820702, 38.0110060291271, 
    42.0719807371405, 36.4255066559906, 40.3254563203728, 34.5335058296867, 
    38.6615140591414, 36.9577513904295, 41.0797406188206, 35.3498813909852, 
    39.3063319434942, 37.7491024143739, 41.5777886205734, 35.8895429100474, 
    40.0721095592252, 38.2719660742721, 42.3176287205335, 36.6920951707497, 
    40.5778445724771, 35.0786710006513, 39.049165272633, 33.432287061478, 
    37.2224728843778, 41.3292461440167, 35.620172988168, 39.5625459179821, 
    38.0110060291271, 42.0719807371405, 36.4255066559906, 40.3254563203728, 
    38.6615140591414, 42.5623103404995, 36.9577513904295, 41.0797406188206, 
    35.3498813909852, 39.3063319434942, 37.7491024143739, 41.5777886205734, 
    35.8895429100474, 40.0721095592252, 38.2719660742721, 42.3176287205335, 
    36.6920951707497, 40.5778445724771, 39.049165272633, 37.2224728843778, 
    41.3292461440167, 35.620172988168, 39.5625459179821, 38.0110060291271, 
    42.0719807371405, 36.4255066559906, 40.3254563203728, 38.6615140591414, 
    42.5623103404995, 36.9577513904295, 41.0797406188206, 39.3063319434942, 
    37.7491024143739, 41.5777886205734, 35.8895429100474, 40.0721095592252, 
    38.2719660742721, 42.3176287205335, 36.6920951707497, 40.5778445724771, 
    39.049165272633, 43.0487719903617, 37.2224728843778, 41.3292461440167, 
    39.5625459179821, 38.0110060291271, 42.0719807371405, 36.4255066559906, 
    40.3254563203728, 38.6615140591414, 42.5623103404995, 36.9577513904295, 
    41.0797406188206, 39.3063319434942, 37.749102414374, 41.5777886205734, 
    40.0721095592252, 38.2719660742721, 42.3176287205335, 36.6920951707497, 
    40.5778445724771, 39.049165272633, 43.0487719903617, 37.2224728843778, 
    41.3292461440167, 39.5625459179821, 38.0110060291271, 42.0719807371405, 
    36.4255066559906, 40.3254563203728, 38.6615140591414, 42.5623103404995, 
    36.9577513904295, 41.0797406188206, 39.3063319434942, 43.2905509512355, 
    37.7491024143739, 41.5777886205734, 40.0721095592252, 38.2719660742721, 
    42.3176287205335, 36.6920951707497, 40.5778445724771, 39.049165272633, 
    43.0487719903617, 37.2224728843778, 41.3292461440167, 39.5625459179821, 
    38.0110060291271, 42.0719807371405, 40.3254563203728, 38.6615140591414, 
    42.5623103404995, 36.9577513904295, 41.0797406188206, 39.3063319434942, 
    43.2905509512355, 37.7491024143739, 41.5777886205734, 40.0721095592252, 
    38.2719660742721, 42.3176287205335, 40.5778445724771, 39.049165272633, 
    43.0487719903617, 37.2224728843778, 41.3292461440167, 39.5625459179821, 
    43.7712030066013, 38.0110060291271, 42.0719807371405, 40.3254563203728, 
    38.6615140591414, 42.5623103404995, 41.0797406188206, 39.3063319434942, 
    43.2905509512355, 37.749102414374, 41.5777886205734, 40.0721095592252, 
    38.2719660742721, 42.3176287205335, 40.5778445724771, 39.049165272633, 
    43.0487719903617, 37.2224728843778, 41.3292461440167, 39.5625459179821, 
    43.7712030066013, 38.0110060291271, 42.0719807371405, 40.3254563203728, 
    38.6615140591414, 42.5623103404995, 41.0797406188206, 39.3063319434942, 
    43.2905509512355, 41.5777886205734, 40.0721095592252, 44.0100754561533, 
    38.2719660742721, 42.3176287205335, 40.5778445724771, 39.049165272633, 
    43.0487719903617, 41.3292461440167, 39.5625459179821, 43.7712030066013, 
    42.0719807371405, 40.3254563203728, 38.6615140591414, 42.5623103404995, 
    41.0797406188206, 39.3063319434942, 43.2905509512355, 41.5777886205734, 
    40.0721095592252, 44.0100754561533, 38.2719660742721, 42.3176287205335, 
    40.5778445724771, 39.049165272633, 43.0487719903617, 41.3292461440167, 
    39.5625459179821, 43.7712030066013, 42.0719807371405, 40.3254563203728, 
    44.2479785386593, 38.6615140591414, 42.5623103404995, 41.0797406188206, 
    39.3063319434942, 43.2905509512355, 41.5777886205734, 40.0721095592252, 
    44.0100754561533, 42.3176287205335, 40.5778445724771, 39.049165272633, 
    43.0487719903617, 41.3292461440167, 39.5625459179821, 43.7712030066013, 
    42.0719807371405, 40.3254563203728, 44.2479785386593, 42.5623103404995, 
    41.0797406188206, 39.3063319434942, 43.2905509512355, 41.5777886205734, 
    40.0721095592252, 44.0100754561533, 42.3176287205335, 40.5778445724771, 
    44.7208760649052, 39.049165272633, 43.0487719903617, 41.3292461440167, 
    39.5625459179821, 43.7712030066013, 42.0719807371405, 40.3254563203728, 
    44.2479785386593, 42.5623103404995, 41.0797406188206, 39.3063319434942, 
    43.2905509512354, 41.5777886205734, 40.0721095592252, 44.0100754561533, 
    42.3176287205335, 40.5778445724771, 44.7208760649052, 43.0487719903617, 
    41.3292461440167, 39.5625459179821, 43.7712030066013, 42.0719807371405, 
    40.3254563203728, 44.2479785386593, 42.5623103404995, 41.0797406188206, 
    44.9558704066931, 39.3063319434942, 43.2905509512355, 41.5777886205734, 
    40.0721095592252, 44.0100754561533, 42.3176287205335, 40.5778445724771, 
    44.7208760649052, 43.0487719903617, 41.3292461440167, 39.5625459179821, 
    43.7712030066013, 42.0719807371405, 40.3254563203728, 44.2479785386593, 
    42.5623103404995, 41.0797406188206, 44.9558704066931, 43.2905509512355, 
    41.5777886205734, 40.0721095592252, 44.0100754561533, 42.3176287205335, 
    40.5778445724771, 44.7208760649052, 43.0487719903617, 41.3292461440167, 
    45.4229504848083, 43.7712030066013, 42.0719807371405, 40.3254563203728, 
    44.2479785386593, 42.5623103404995, 41.0797406188206, 44.9558704066931, 
    43.2905509512355, 41.5777886205734, 44.0100754561533, 42.3176287205335, 
    40.5778445724771, 44.7208760649052, 43.0487719903617, 41.3292461440167, 
    45.4229504848083, 43.7712030066013, 42.0719807371405, 40.3254563203728, 
    44.2479785386593, 42.5623103404995, 41.0797406188206, 44.9558704066931, 
    43.2905509512355, 41.5777886205734, 45.6550365094507, 44.0100754561533, 
    42.3176287205335, 40.5778445724771, 44.7208760649052, 43.0487719903617, 
    41.3292461440167, 45.4229504848083, 43.7712030066013, 42.0719807371405, 
    40.3254563203728, 44.2479785386593, 42.5623103404995, 41.0797406188206, 
    44.9558704066931, 43.2905509512355, 41.5777886205734, 45.6550365094507, 
    44.0100754561533, 42.3176287205335, 40.5778445724771, 44.7208760649052, 
    43.0487719903617, 41.3292461440167, 45.4229504848083, 43.7712030066013, 
    42.0719807371405, 46.0012276067282, 44.2479785386593, 42.5623103404995, 
    41.0797406188206, 44.9558704066931, 43.2905509512354, 41.5777886205734, 
    45.6550365094507, 44.0100754561533, 42.3176287205335, 40.5778445724771, 
    44.7208760649052, 43.0487719903617, 41.3292461440167, 45.4229504848083, 
    43.7712030066013, 42.0719807371405, 46.0012276067282, 44.2479785386593, 
    42.5623103404995, 44.9558704066931, 43.2905509512354, 41.5777886205734, 
    45.6550365094507, 44.0100754561533, 42.3176287205335, 46.3454815789384, 
    44.7208760649052, 43.0487719903617, 41.3292461440167, 45.4229504848084, 
    43.7712030066013, 42.0719807371405, 46.0012276067282, 44.2479785386593, 
    42.5623103404995, 44.9558704066931, 43.2905509512355, 41.5777886205734, 
    45.6550365094507, 44.0100754561533, 42.3176287205335, 46.3454815789384, 
    44.7208760649052, 43.0487719903617, 45.4229504848083, 43.7712030066013, 
    42.0719807371405, 46.0012276067282, 44.2479785386593, 42.5623103404995, 
    46.6873156862054, 44.9558704066931, 43.2905509512355, 41.5777886205734, 
    45.6550365094507, 44.0100754561533, 42.3176287205335, 46.3454815789384, 
    44.7208760649052, 43.0487719903617, 45.4229504848084, 43.7712030066013, 
    42.0719807371405, 46.0012276067282, 44.2479785386593, 42.5623103404995, 
    46.6873156862054, 44.9558704066931, 43.2905509512355, 45.6550365094507, 
    44.0100754561533, 42.3176287205335, 46.3454815789384, 44.7208760649052, 
    43.0487719903617, 45.4229504848083, 43.7712030066013, 42.0719807371405, 
    46.0012276067282, 44.2479785386593, 42.5623103404995, 46.6873156862054, 
    44.9558704066931, 43.2905509512355, 45.6550365094507, 44.0100754561533, 
    42.3176287205335, 46.3454815789384, 44.7208760649052, 43.0487719903617, 
    45.4229504848084, 43.7712030066013, 42.0719807371405, 46.0012276067282, 
    44.2479785386593, 42.5623103404995, 46.6873156862054, 44.9558704066931, 
    43.2905509512354, 45.6550365094507, 44.0100754561533, 42.3176287205335, 
    46.3454815789384, 44.7208760649052, 43.0487719903617, 45.4229504848083, 
    43.7712030066013, 46.0012276067282, 44.2479785386593, 42.5623103404995, 
    46.6873156862054, 44.9558704066931, 43.2905509512355, 45.6550365094507, 
    44.0100754561533, 42.3176287205335, 46.3454815789384, 44.7208760649052, 
    43.0487719903616, 45.4229504848083, 43.7712030066013, 46.0012276067282, 
    44.2479785386593, 42.5623103404995, 46.6873156862054, 44.9558704066931, 
    43.2905509512355, 45.6550365094507, 44.0100754561533, 46.3454815789384, 
    44.7208760649052, 43.0487719903617, 45.4229504848084, 43.7712030066013, 
    46.0012276067282, 44.2479785386593, 42.5623103404995, 46.6873156862054, 
    44.9558704066931, 43.2905509512355, 45.6550365094507, 44.0100754561533, 
    46.3454815789384, 44.7208760649052, 43.0487719903617, 45.4229504848083, 
    43.7712030066013, 46.0012276067282, 44.2479785386593, 46.6873156862054, 
    44.9558704066931, 43.2905509512355, 45.6550365094507, 44.0100754561533, 
    46.3454815789384, 44.7208760649052, 43.0487719903617, 45.4229504848083, 
    43.7712030066013, 46.0012276067282, 44.2479785386593, 46.6873156862054, 
    44.9558704066931, 43.2905509512355, 45.6550365094507, 44.0100754561533, 
    46.3454815789384, 44.7208760649052, 45.4229504848084, 43.7712030066013, 
    46.0012276067282, 44.2479785386593, 46.6873156862054, 44.9558704066931, 
    43.2905509512355, 45.6550365094507, 44.0100754561533, 46.3454815789384, 
    44.7208760649052, 45.4229504848083, 43.7712030066013, 46.0012276067282, 
    44.2479785386593, 46.6873156862054, 44.9558704066931, 43.2905509512355, 
    45.6550365094507, 44.0100754561533, 46.3454815789384, 44.7208760649052, 
    45.4229504848083, 43.7712030066013, 46.0012276067282, 44.2479785386593, 
    46.6873156862054, 44.9558704066931, 45.6550365094507, 44.0100754561533, 
    46.3454815789384, 44.7208760649052, 45.4229504848084, 43.7712030066013, 
    46.0012276067282, 44.2479785386593, 46.6873156862054, 44.9558704066931, 
    45.6550365094507, 44.0100754561533, 46.3454815789384, 44.7208760649052, 
    45.4229504848084, 46.0012276067282, 44.2479785386593, 46.6873156862054, 
    44.9558704066931, 45.6550365094507, 44.0100754561533, 46.3454815789384, 
    44.7208760649052, 45.4229504848083, 46.0012276067282, 44.2479785386593, 
    46.6873156862054, 44.9558704066931, 45.6550365094507, 46.3454815789384, 
    44.7208760649052, 45.4229504848083, 46.0012276067282, 44.2479785386593, 
    46.6873156862054, 44.9558704066931, 45.6550365094507, 46.3454815789384, 
    44.7208760649052, 45.4229504848084, 46.0012276067282, 46.6873156862054, 
    44.9558704066931, 45.6550365094507, 46.3454815789384, 44.7208760649052, 
    45.4229504848083, 46.0012276067282, 46.6873156862054, 44.9558704066931, 
    45.6550365094507, 46.3454815789384, 45.4229504848083, 46.0012276067282, 
    46.6873156862054, 44.9558704066931, 45.6550365094507, 46.3454815789384, 
    45.4229504848083, 46.0012276067282, 46.6873156862054, 44.9558704066931, 
    45.6550365094507, 46.3454815789384, 45.4229504848083, 46.0012276067282, 
    46.6873156862054, 45.6550365094507, 46.3454815789384, 45.4229504848084, 
    46.0012276067282, 46.6873156862054, 45.6550365094507, 46.3454815789384, 
    46.0012276067282, 46.6873156862054, 45.6550365094507, 46.3454815789384, 
    46.0012276067282, 46.6873156862054, 46.3454815789384, 46.6873156862054, 
    46.3454815789384, 46.6873156862054, 46.3454815789384, 46.6873156862054 ;

 obs_type = 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 7, 7, 7, 7, 7, 
    7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 
    7, 7, 7, 7, 7, 7, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 
    7, 7, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 7, 7, 7, 7, 
    7, 7, 7, 6, 6, 6, 6, 6, 6, 6, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    7, 7, 7, 7, 7, 7, 7, 7, 7, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1 ;

 obs_error = 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.169206023673944, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.236255327678716, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.17556760861175, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.223196763845215, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.235533601422048, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.228712343216355, 
    0.235744558228311, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.171836779133628, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.162895037797164, 0.16, 0.16, 0.16, 0.16, 0.16, 0.308477104980401, 
    0.166997650688514, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.420906402871828, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.171623836939502, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.231263474606969, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.255906707668323, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.180739066770684, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.27305871365506, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.210282059700098, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.168947220181749, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.326175480240323, 0.182336397522704, 0.841617820109869, 
    0.366017024386714, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.623906398614281, 0.431207267386656, 0.16, 0.16, 0.16, 
    0.177744377255522, 0.18731242704398, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.344668699428943, 0.16, 0.16, 0.16, 0.1875, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.203616172396576, 
    0.182449070394366, 0.404810133831867, 0.16, 0.740713460286497, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.265203209058028, 0.302222301430447, 
    0.16, 0.16, 0.427500114441024, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.620789541319744, 0.311053361730535, 0.16, 0.225260973199566, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.426319582634096, 0.379140454928221, 
    0.223218806743733, 0.16, 1.12154779706686, 0.16, 1.14083316802983, 0.16, 
    0.16, 0.170368834762154, 0.16, 0.175736671657219, 0.567207416934328, 
    0.51060831967175, 0.203242975359103, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.181969531788809, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.173249823331889, 0.16, 0.196412271437081, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.258867296792914, 0.16, 0.01, 0.01, 0.01, 0.01, 
    0.324375324438734, 0.0121287765138732, 0.038382151443966, 
    0.0240197479604376, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    1.62889755259069, 0.0419550288354458, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0504894010198768, 0.0221785731046111, 0.00233577516773949, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.00138104300034077, 0.0001, 0.01, 0.01, 0.01, 0.01, 1.65763796959436, 
    0.189741286346634, 0.048849569938443, 0.01, 0.0358767342185502, 
    0.058099554037949, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.0001, 0.0001, 0.0001, 0.0001, 0.0017334126799445, 
    0.0272445019581937, 0.0356001375475898, 0.00522243865998462, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.170362611578033, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.231153241230707, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.236314026755609, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.168976922597216, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.236366940216031, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.17166405154689, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.165160361550926, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.425309012322209, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.180274257448211, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.252474126695068, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.259657617495375, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.341411981870082, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.425859563795815, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.189787504936653, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.190438281970163, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.306693419502507, 0.163760513292607, 0.736021128966869, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.623906398614281, 
    0.431207267386656, 0.16, 0.16, 0.16, 0.16, 0.173249955654228, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.317612613250406, 0.16, 
    0.16, 0.16, 0.1875, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.209003817931969, 0.182449070394366, 0.404810133831867, 0.16, 
    0.740713460286497, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.265203209058028, 0.302222301430447, 0.16, 0.16, 0.427500114441024, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.620789541319744, 
    0.311053361730535, 0.16, 0.225260973199566, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.426319582634096, 0.417856958934457, 0.223218806743733, 0.16, 
    1.12154779706686, 0.16, 1.14083316802983, 0.16, 0.16, 0.170368834762154, 
    0.16, 0.175736671657219, 0.556349767466951, 0.51060831967175, 
    0.203242975359103, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.188555043171618, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.173249823331889, 
    0.16, 0.196412271437081, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.17800923363263, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.17775111871942, 0.16, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.01, 
    0.01, 0.01, 0.01, 0.0156910209739181, 0.0438008630647649, 
    0.547292163201109, 0.01, 0.01, 0.0314631155523557, 0.0151807135847169, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.000624001098913141, 
    0.0338037966459524, 0.0263323568316991, 0.00419089860952226, 
    0.000151686307799537, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.01, 0.01, 
    0.0297230925192713, 0.01, 0.01, 0.01, 0.01, 0.24514808984577, 
    0.019256473790154, 0.01, 0.01, 0.01, 0.0154299090933584, 
    0.0226917920130563, 0.0147561568154877, 0.01, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.167758493312198, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.218476031769064, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.253970290586694, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.188556690375325, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.387052559211043, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.22082990681889, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.168922335643806, 0.16, 0.16, 0.16, 0.16, 0.268183449650678, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.262984531641855, 0.16, 0.16, 0.16, 
    0.16, 0.166218503489694, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.197824004295878, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.21219825571601, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.171913918265311, 
    0.175010843616946, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.178992779608507, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.164015345904828, 0.16, 0.16, 0.16, 0.16, 
    0.175879345169278, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.635867754907122, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.172933733402274, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.180385724258734, 
    0.266562116742534, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    1.85281286716463, 0.307151112715443, 0.16, 0.16, 0.16, 0.16, 
    0.173249955654228, 0.16, 0.16, 0.16, 0.16, 0.16, 0.236560948623365, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.433475232442288, 0.16, 0.16, 0.16, 0.1875, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.209003817931969, 0.215377181021369, 
    0.392152663601792, 0.16, 0.740713460286497, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.180353030772818, 
    0.16, 0.16, 0.194176510876754, 0.16, 0.365316369772144, 0.16, 
    0.468000037193633, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.620789541319744, 0.311053361730535, 0.16, 0.225260973199566, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.491905725717697, 0.417856958934457, 
    0.165017488267823, 0.28125, 1.36124937057502, 0.16, 0.16, 
    0.170368834762154, 0.16, 0.175736671657219, 0.556349767466951, 
    0.51060831967175, 0.203242975359103, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.193488433406502, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.173249823331889, 0.16, 0.196412271437081, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.175906727605004, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.164341237621102, 0.16, 0.16, 0.16, 0.240545853331848, 
    0.16, 0.16, 0.16, 0.25061127991992, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.229806806459753, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.0688564273720011, 0.0211968311302344, 0.0321866176903616, 
    0.0439302069940496, 0.0189343745927172, 0.0284255121212581, 
    0.0495865738129722, 0.0279395934441173, 0.0217164937494265, 
    0.113565808354486, 0.0328322511322492, 0.0464301975957755, 
    0.0277489334581181, 0.01, 0.01, 0.01, 0.01, 0.01, 0.0941105779414708, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.01, 0.01, 0.01, 0.01, 0.01, 0.01, 
    0.0548090222587234, 0.0316542262025905, 0.0148340101627582, 0.0001, 
    0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0040500137329218, 
    0.00884493024204858, 0.00414046389778378, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.161494834401866, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.181779190759471, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.204750810126136, 0.16, 0.214176758009671, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.172032629036425, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.234138924188629, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.164342905655177, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.170321954357658, 0.173788603214462, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.411187648673831, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.186857271570489, 0.16, 0.16, 0.16, 
    0.16, 0.280361056149205, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.216000270656145, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.179386209794233, 0.176948346328152, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.170538680574771, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.175471568958549, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.208095779020798, 0.18113227749968, 0.16, 0.16, 
    0.161913314600745, 0.330000085830718, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.255720028948417, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.178928526469723, 0.16, 0.20812522888203, 
    0.16, 0.16, 0.16, 0.619104246457482, 0.403072977860802, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.162498701384215, 0.16, 
    0.181687655925816, 0.16, 0.16, 0.243416638692361, 0.16, 0.16, 
    0.209003817931969, 0.215377181021369, 0.216501779556388, 0.16, 
    0.631827416931044, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.170457777174559, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.203557247767941, 0.16, 
    0.224656370163046, 0.278738629818106, 0.302562340736495, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.620789541319744, 0.311053361730535, 0.16, 
    0.203623897367992, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.247499814033563, 
    0.186749908447382, 0.16, 0.16, 0.16, 0.170368834762154, 0.16, 
    0.175736671657219, 0.556349767466951, 0.51060831967175, 
    0.203242975359103, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.237740099601852, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.173249823331889, 
    0.16, 0.196412271437081, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.170997930777528, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.190835307095182, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.446182357798484, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.170163644763279, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.220951519713526, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.172033131606693, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.16, 0.181123597304602, 0.16, 0.16, 
    0.16, 0.16, 0.16, 0.01, 0.01, 0.01, 0.01, 0.01, 2.22978286072005, 0.01, 
    0.110309041844024, 0.0295305330382689, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0001, 0.00360850169090554, 0.0001, 0.0438204756792402, 
    0.00819178906385787, 0.0341147000726778, 0.01, 0.01, 0.01, 0.01, 
    1.20238138122841, 0.01, 0.0131558080029208, 0.0694856064951637, 0.01, 
    0.01, 0.01, 0.01, 0.01, 0.01, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.00145784015330719, 0.0226847665107925, 0.0139444694214035, 
    0.0030419309696299, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 0.0001, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.000732873089436909, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.00178545430973173, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.00222919926121832, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0017237827368197, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.000618576550867875, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.00146547146141529, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.00319360671211034, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.00344839172363281, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.00312514992430806, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.00306183930981205, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.00215113790524192, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.000772919896536042, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.000453614406473938, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.000614632743236143, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.000491725297656379, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 0.0004, 
    0.0004, 0.0004, 0.0004, 0.0004 ;

 obs_value = 17.8686498006185, 17.8131071726481, 17.8617830276489, 
    17.6225627263387, 17.1223834355672, 16.9473829269409, 16.7027254104614, 
    16.6388298670451, 16.740306854248, 16.4919951756795, 16.374140103658, 
    16.3761348724365, 16.0612738927205, 15.6583701769511, 15.605455716451, 
    14.8883198102315, 14.4206415812174, 14.3832081158956, 13.8395233154297, 
    13.6499096552531, 13.1701434453328, 13.2680602073669, 13.2600247065226, 
    13.4456125895182, 13.3635026613871, 13.4539214769999, 13.7342659632365, 
    13.0989408493042, 12.7016830444336, 12.7761775652568, 11.9570039113363, 
    11.7327136993408, 11.5222371419271, 11.249197324117, 10.9549608230591, 
    10.781909942627, 10.7043263117472, 10.7628067334493, 10.7439735730489, 
    11.2142833073934, 11.1918082237244, 10.9110434850057, 11.1261164347331, 
    10.8196873664856, 10.6027889251709, 10.2856755256653, 10.4315498669942, 
    9.87392600377401, 9.83848222096761, 9.58017428716024, 9.37397400538127, 
    17.902720981174, 17.7539225684272, 17.6760533650716, 17.5449314117432, 
    17.1177950965034, 16.8860143025716, 16.5799312591553, 16.5810521443685, 
    16.5950130886502, 16.4062904781765, 16.321013768514, 16.3073289659288, 
    16.1882004208035, 15.6307292514377, 15.5051152971056, 15.1281949149238, 
    14.4904933505588, 14.5163915952047, 14.2146603266398, 13.8862502574921, 
    13.6025365193685, 13.6202226479848, 13.5435059865316, 13.5756066640218, 
    13.5631836255391, 13.6322495142619, 13.5650587876638, 12.8016896247864, 
    12.4629538853963, 12.210329691569, 12.2411887645721, 11.8469492594401, 
    11.5793776512146, 11.5222968260447, 11.1392214298248, 10.9604073365529, 
    10.7619397640228, 10.9713776906331, 11.0695140361786, 11.1925318241119, 
    10.9902223745982, 11.0476109981537, 11.0335791905721, 10.7934989134471, 
    10.435835202535, 10.4300451278687, 10.1385598977407, 10.0796749591827, 
    9.62425168355306, 9.66027688980103, 9.58813381195068, 17.6685240003798, 
    17.5441362592909, 17.4093339708116, 17.3339163462321, 17.0588575998942, 
    16.579709370931, 16.4384117126465, 16.5931549072266, 16.5161732567681, 
    16.3779218461778, 16.3396731482612, 16.2868169148763, 16.3915076785617, 
    15.9734265009562, 15.6506340238783, 15.1115172704061, 14.8780102199978, 
    14.8882077534993, 14.7659137248993, 14.3006910483042, 14.0097931226095, 
    13.9310528437297, 13.9156708717346, 13.8826749324799, 13.5762342611949, 
    13.4387756983439, 13.2277731100718, 12.4343460400899, 12.3752910296122, 
    12.377716700236, 12.164178053538, 11.8559877872467, 11.7691961129506, 
    11.718638420105, 11.1890168190002, 11.1178963184357, 11.0474449793498, 
    11.1153093179067, 11.2982345422109, 11.3646145661672, 11.2251887321472, 
    11.0229583581289, 10.6965347131093, 10.7022506395976, 10.3992682298025, 
    10.0641298294067, 9.94975781440735, 9.72301204999288, 9.77265508969625, 
    9.88398782412211, 9.82052246729533, 17.8643211788601, 17.5660885704888, 
    17.3851555718316, 17.1644221411811, 16.8518784840902, 16.4433966742622, 
    16.2801149156358, 16.3657266828749, 16.4109128316243, 16.3826620313856, 
    16.2061865064833, 16.2727419535319, 16.276765399509, 16.0027279324002, 
    15.582453833686, 15.4504129621718, 15.1324907938639, 15.018320719401, 
    14.1425299114651, 13.5889497333103, 13.6990977393256, 14.0432945887248, 
    13.7892492082384, 13.6638476053874, 13.5874565972222, 13.256067276001, 
    12.8657422595554, 12.2033785714044, 12.1095161437988, 11.7979148228963, 
    11.6323902342055, 11.3136403825548, 11.4431229697333, 11.8368631998698, 
    11.263252682156, 11.4188646740384, 11.0170679092407, 11.4953223334418, 
    11.5026312934028, 10.899735238817, 11.153423945109, 10.9864328172472, 
    10.9134111404419, 10.4472222858005, 10.1945996814304, 9.97936598459879, 
    9.60224363538954, 9.62567117479112, 9.86019388834635, 9.98873117234972, 
    9.98170778486464, 18.0199442969428, 17.7590065002441, 17.2391632927789, 
    16.8445248074002, 16.6465733846029, 16.4957205454508, 16.0748896068997, 
    16.2683410644531, 16.3235003153483, 16.2869290245904, 16.1319358613756, 
    16.2453132205539, 16.1663838492499, 15.8937543233236, 15.710226588779, 
    15.5261217753092, 15.2293580373128, 14.3206237157186, 13.3676670392354, 
    13.1091509660085, 13.2072250048319, 13.5499849319458, 13.6086343129476, 
    13.6254851818085, 13.3893189430237, 12.8595005671183, 12.4759302934011, 
    12.338770866394, 11.7873073418935, 11.3035844167074, 11.2414281368256, 
    11.0850691000621, 11.0477206707001, 11.1969409783681, 11.3570636113485, 
    11.1844186782837, 10.8272945086161, 10.9952200253805, 11.0786762237549, 
    10.8792855739594, 10.9872721036275, 10.7128615379333, 10.6246434052785, 
    9.94160429636637, 9.72100361188253, 9.53459604581197, 9.4722912311554, 
    9.65840101242065, 9.6197235584259, 9.88399235407511, 9.98665579160055, 
    17.7009154425727, 17.5789824591743, 17.1332092285156, 16.9326489766439, 
    16.8175843556722, 16.5973731146918, 16.1374693976508, 16.3025512695312, 
    16.2559343973796, 16.1199090745714, 16.0837603674995, 16.0409804450141, 
    15.9943709903293, 15.673135333591, 15.5815919240316, 15.2156396441989, 
    14.5940988328722, 13.59010887146, 13.0655469894409, 12.9491009712219, 
    13.1538377602895, 13.4721104303996, 13.5177763303121, 13.6241952578227, 
    13.3411426544189, 12.5562081336975, 12.2922523021698, 11.9097426732381, 
    11.3092327912649, 11.2333728472392, 11.1744136810303, 11.2402401765188, 
    10.8076803684235, 11.0387280782064, 11.033539613088, 10.934552192688, 
    10.7047639687856, 10.7170461813609, 10.8562707901001, 10.8051074345907, 
    10.6753590901693, 10.5273989836375, 10.0264480908712, 9.84856613477071, 
    9.86593238512675, 9.51769963900248, 9.53892199198405, 9.62269139289856, 
    9.78984610239665, 9.69866625467936, 9.90589157740275, 17.6028116014269, 
    17.6113736894396, 17.3912599351671, 16.8856870863173, 16.8895681169298, 
    16.6807166205512, 16.1919623480903, 16.2148068745931, 16.0463875664605, 
    15.8665758768717, 15.8888018925985, 15.9329424964057, 15.6039623684353, 
    15.4220310846965, 15.4123918745253, 15.0238551033868, 13.74520556132, 
    13.0483843485514, 12.989968723721, 13.1687825520833, 13.3401367399428, 
    13.4320959515042, 13.5714970694648, 13.5118360519409, 13.2521700329251, 
    12.6334020826552, 11.8846242692735, 11.2785120010376, 11.1115425957574, 
    11.2083404329088, 11.1808550092909, 11.3472635481093, 11.0289876725939, 
    10.909107208252, 10.7710780037774, 10.6348027123345, 10.6212383906047, 
    10.7047668033176, 10.9113020367093, 10.8953300052219, 10.6949564615885, 
    10.3004207611084, 9.89880996280246, 10.0633770624797, 10.1181305779351, 
    9.88602574666341, 9.72119808197021, 9.7685522503323, 9.79260084364149, 
    9.20212512546115, 9.40839693281386, 17.7412052154541, 17.6021075778537, 
    17.3496534559462, 16.9679419199626, 16.8956127166748, 16.633267932468, 
    16.2120193905301, 16.1111454433865, 15.7553897433811, 15.7244053946601, 
    15.904599931505, 15.7626298268636, 15.6105767356025, 15.5001724031236, 
    15.0587934917874, 14.551583925883, 13.2095504336887, 12.9099601904551, 
    13.1324632962545, 13.3077109654744, 13.4097334543864, 13.3170934518178, 
    13.3796151479085, 13.2215209007263, 13.102506796519, 12.2115104198456, 
    11.4274423917135, 11.1176384290059, 11.1875011920929, 11.1681145826975, 
    11.2096800804138, 11.2104723453522, 11.1818552017212, 10.8214148680369, 
    10.6481671333313, 10.5365335146586, 10.7371890544891, 10.7612276871999, 
    10.7428054014842, 11.0097764333089, 10.8647513389587, 10.7389195760091, 
    10.3815069993337, 10.0843800703684, 10.2859400908152, 10.0456237792969, 
    9.72928563753764, 9.60072875022888, 9.27522460619609, 9.26683020591736, 
    9.84079869588216, 17.8264122009277, 17.6364163292779, 17.6271606021457, 
    17.259800169203, 16.9632778167725, 16.4979864756266, 16.230035993788, 
    16.0902796851264, 15.8471589618259, 15.8726453781128, 15.7299062940809, 
    14.9159389071994, 15.095788107978, 15.2666282653809, 15.0101013183594, 
    14.0720207426283, 13.042195532057, 12.7828991413116, 13.1682035923004, 
    13.4103170235952, 13.3750964005788, 13.30495540301, 13.3638764222463, 
    13.3633289337158, 12.8981987635295, 11.7944509188334, 11.2285717328389, 
    11.065572977066, 11.2689394950867, 11.3391540845235, 11.2757557233175, 
    11.1330415407817, 11.1177975336711, 10.8609031836192, 10.6383199691772, 
    10.8754473527273, 10.638486067454, 10.6567704677582, 10.6553152402242, 
    10.8320926030477, 10.9443678855896, 10.7345778942108, 10.4634408950806, 
    10.2523949146271, 10.250873486201, 10.0680010318756, 9.79902680714925, 
    9.32157532374064, 8.79749234517415, 9.53988711039225, 10.0852352778117, 
    17.8208457099067, 17.6720951928033, 17.5554358164469, 17.2240113152398, 
    16.7869582706028, 16.3353231218126, 16.3282324473063, 16.1936158074273, 
    16.0250906414456, 15.7660064697266, 15.0044167836507, 14.6308188968235, 
    14.6093427870009, 15.1613915761312, 15.0414596133762, 13.7811891767714, 
    13.0439778433906, 12.5793139139811, 13.0025089051988, 13.3656131956312, 
    13.309105237325, 13.2741913265652, 13.1729532877604, 13.0002508163452, 
    12.6922752592299, 11.6331615447998, 11.0862038930257, 11.0864955054389, 
    11.3518313301934, 11.4748825497097, 11.237471792433, 11.1656413608127, 
    11.1809567345513, 10.7635019090441, 10.631396929423, 10.5984117719862, 
    10.5454712973701, 10.4675868352254, 10.658835305108, 10.8727882173326, 
    11.0236953099569, 10.6267618603177, 10.433439678616, 10.5103601879544, 
    10.0601825714111, 10.017853418986, 10.0602272881402, 9.47212759653727, 
    9.24998537699381, 10.0335140228271, 10.028789308336, 17.806751675076, 
    17.5662708282471, 17.4335505167643, 17.3674023946126, 17.2081707848443, 
    16.6736867692735, 16.5820914374457, 16.3212912877401, 15.848478741116, 
    15.3983489142524, 14.7520723342896, 14.6551904678345, 14.3877025180393, 
    14.4336366653442, 14.5765027999878, 13.442386203342, 13.1544272104899, 
    12.6320009231567, 12.5607833862305, 12.9405498504639, 13.1890299320221, 
    13.1316666603088, 13.0223200321198, 12.882461309433, 12.6328237056732, 
    11.6320850849152, 11.1299397150675, 11.1505583922068, 11.3746054967244, 
    11.6599852244059, 11.3427301247915, 11.5044706662496, 11.2542022864024, 
    11.006786108017, 10.6719636122386, 10.6243744691213, 10.5895075798035, 
    10.4794416427612, 10.8959666093191, 10.7225592931112, 10.5128107070923, 
    10.4009798367818, 10.4326225916545, 10.3359718322754, 10.1406003634135, 
    10.0445350805918, 9.8684667746226, 9.6552050113678, 9.75360989570618, 
    10.2284070650736, 9.95206395785014, 17.4773616790771, 17.439728418986, 
    17.3446824815538, 17.4639818403456, 17.4404021369086, 17.1504692501492, 
    16.7966232299805, 16.2445588641697, 15.6625797483656, 15.131136364407, 
    14.5887150234646, 14.556719356113, 14.2977734671699, 14.0645848380195, 
    13.9321426815457, 13.2347113291423, 13.129828453064, 12.6229612827301, 
    12.5664873917898, 12.5571709473928, 13.017871538798, 12.937243382136, 
    12.8408591747284, 12.8055454889933, 12.4790213108063, 11.7397116820017, 
    11.2407761414846, 11.4613250096639, 11.9286359151204, 12.0463620821635, 
    11.2490148544312, 11.3920844395955, 11.3825311660767, 11.0961714585622, 
    10.8651951948802, 10.6444195906321, 10.7374013264974, 10.5873325665792, 
    10.8382159868876, 10.7148042519887, 10.5115649700165, 10.4034101963043, 
    10.412383556366, 10.3893005847931, 10.2036020755768, 10.0885475476583, 
    9.91014615694682, 9.42600893974304, 10.1750884056091, 10.3201859792074, 
    10.0052728652954, 17.1840029822456, 17.3383384280735, 17.2045665317112, 
    17.2749262915717, 17.3671120537652, 17.2288265228271, 16.6493184831407, 
    16.1576750013563, 15.6531579759386, 14.8095438215468, 14.5511629316542, 
    14.5960733625624, 14.2198066711426, 14.2272093031141, 14.0841466055976, 
    13.3366684383816, 13.1227495405409, 12.7298672993978, 12.9693313174778, 
    12.7153290642632, 12.726454310947, 12.8297713597616, 12.6739433076647, 
    12.6370987362332, 12.3672902848985, 12.1135889689128, 11.854240099589, 
    12.120166460673, 12.30351946089, 12.1950885984633, 11.1856772104899, 
    10.9993022282918, 11.1989393234253, 11.0322364171346, 11.0713130103217, 
    10.6779696146647, 11.0253166622586, 10.9325436486138, 11.0269550747342, 
    11.0111149681939, 10.6976925532023, 10.4212410185072, 10.4820054372152, 
    10.2026970121596, 9.98784690433078, 10.2526546054416, 10.2286703321669, 
    9.81193044450548, 10.3288114335802, 10.1794766320123, 9.80511336856418, 
    16.9263485802544, 17.2302186754015, 17.1730774773492, 17.3546373579237, 
    17.4236189524333, 17.1738957299127, 16.4787108103434, 16.2181760999892, 
    15.8224564658271, 14.8799469206068, 14.6637399461534, 14.6929047902425, 
    14.1821202172173, 14.2238669925266, 14.2059072918362, 13.545115047031, 
    13.1697787178887, 12.8228424390157, 13.2275823752085, 12.9264861742655, 
    12.5462508201599, 12.5235587755839, 12.5382173061371, 12.700515349706, 
    12.7435689767202, 12.7285847663879, 12.533770720164, 11.7227299213409, 
    11.72798426946, 11.5600167115529, 11.0773317813873, 10.9342215061188, 
    10.7637391885122, 10.9474337100983, 10.7288604216142, 10.6729708512624, 
    9.99999986376081, 10.1999998092651, 10.2910713468279, 10.533749961853, 
    10.428658246994, 10.3317415714264, 10.9522763888041, 10.4354976926531, 
    9.99507403373718, 9.85002794265747, 9.3729043006897, 9.74030009183017, 
    9.82614785974676, 9.86240369623358, 9.54256304105123, 16.7831810845269, 
    16.7887465159098, 16.8574470943875, 17.0785927242703, 17.2093717787001, 
    16.8833484649658, 16.4858462015788, 16.1154221428765, 15.9110057618883, 
    15.1512944963243, 14.5927799012926, 14.5875798331367, 14.2906640370687, 
    14.2880047692193, 14.302638053894, 13.6480691697862, 13.4153170055813, 
    12.960916519165, 13.2307871977488, 13.1495540142059, 12.5491460164388, 
    12.3106647332509, 12.3542804718018, 12.4939960638682, 12.8044987519582, 
    12.8055377006531, 12.1909607251485, 11.3653008937836, 11.3768981297811, 
    11.2964475154877, 11.2066859404246, 10.9633156458537, 10.8241041501363, 
    11.0431148355657, 10.6669385433197, 10.5407814184825, 10.1969999313354, 
    10.2910714830671, 10.178750038147, 10.375, 10.2679562568665, 
    10.2842186689377, 9.23125004768372, 9.44553579602923, 9.59716653823853, 
    9.36710691452026, 9.75086291631063, 9.14531254768372, 9.71999988555908, 
    16.8455515967475, 16.670398288303, 16.5924254523383, 16.7193902333577, 
    16.9921724531386, 17.0061558617486, 16.7068116929796, 16.2812455495199, 
    16.0771551132202, 15.2430523766412, 14.8340001636081, 14.5557398266262, 
    14.1941146850586, 14.3197728263007, 14.3050056033664, 13.815357208252, 
    13.453172577752, 13.2799819310506, 13.3244272867839, 13.2742685741848, 
    12.7056620915731, 12.4720680448744, 12.2622829013401, 12.4706433614095, 
    12.721126238505, 12.8023256725735, 11.7744862238566, 11.2716440624661, 
    11.5676364898682, 11.6010559929742, 11.4533996582031, 10.6454860899183, 
    10.9812501271566, 11.2478250927395, 10.8089843988419, 10.6052098274231, 
    10.3124081747872, 10.0362501144409, 11.0500001907349, 10.2791666984558, 
    10.3552083969116, 9.75, 10.1999998092651, 9.75749988555908, 
    9.70666631062826, 9.76518938276503, 9.79342608981662, 10.1500220828586, 
    9.88437521457672, 9.82392480638292, 9.77708339691162, 16.8266201019287, 
    16.6703048282199, 16.5996913909912, 16.5696125030518, 16.730989880032, 
    16.6187121073405, 16.3444904751248, 16.2734188503689, 16.3026496039497, 
    15.3992634879218, 14.9586522844103, 14.4224809010824, 14.101053237915, 
    14.3224902682834, 14.4494726392958, 14.1119792726305, 13.6111681196425, 
    13.430597225825, 13.433385848999, 13.249836842219, 12.7235169410706, 
    12.5479542414347, 12.3736299673716, 12.2824199994405, 12.4724773565928, 
    12.6209418773651, 11.5942851702372, 11.2586677869161, 11.7538615862528, 
    11.7440587679545, 11.3050923877292, 11.4008680184682, 11.0583333969116, 
    11.1414774114435, 10.8548458947076, 9.69999994550433, 9.99892861502511, 
    10.1999998092651, 10.3078126907349, 9.95000004768372, 9.61514854431152, 
    9.60738393995497, 9.91185609499613, 9.77400024731954, 9.18947919209798, 
    9.72964421908061, 9.82457224527995, 9.37186543146769, 16.8794000413683, 
    16.6359712812636, 16.5487177107069, 16.426879035102, 16.366141849094, 
    16.1442111333211, 16.1457302305434, 16.2361077202691, 16.4487692515055, 
    15.7744834687975, 15.3182440863715, 14.1497858895196, 13.9635717603895, 
    14.0594823625353, 13.9738202624851, 13.8740448421902, 13.7653101815118, 
    13.6771697998047, 13.4317735036214, 13.313229004542, 12.7764935493469, 
    12.4558240572611, 12.472663640976, 12.5351433753967, 12.6020941734314, 
    12.4170015652974, 11.7714300950368, 11.5159757932027, 11.6049584547679, 
    10.8580003738403, 11.5541666878594, 11.1625001213767, 10.8682735988072, 
    9.87142876216343, 9.09999990463257, 10.483333269755, 9.8746874332428, 
    9.73693171414462, 9.60545444488525, 9.44629796346029, 8.29400690396627, 
    8.48249777158101, 8.63380159031261, 8.3155323266983, 16.9477994706896, 
    16.7322296566433, 16.7102896372477, 16.4096588558621, 16.2166614532471, 
    16.132671462165, 15.9399919509888, 16.3124287923177, 16.0978140301175, 
    15.7933065626356, 15.2180204391479, 14.1952080196804, 13.8165542814467, 
    13.7741102642483, 13.6997520658705, 13.654659377204, 13.744639078776, 
    13.6563516192966, 13.0154858695136, 12.8971887164646, 12.8131279415554, 
    12.4989048639933, 12.3425937228733, 12.2767884996202, 11.9908799065484, 
    11.9892830318875, 11.7684735192193, 11.604575475057, 8.24499979019165, 
    8.83703136444092, 8.65571673711141, 8.13243993123372, 16.9899828169081, 
    16.9137054019504, 16.7561863793267, 16.5123842027452, 16.3484032948812, 
    16.2034346262614, 16.205540339152, 16.0671242607964, 15.7848572201199, 
    15.2138847774929, 14.6135743459066, 14.1822698381212, 14.0229782528347, 
    13.8245691723294, 13.6361236572266, 13.361542807685, 13.5420999526978, 
    13.6583212216695, 13.0707894166311, 12.8432679971059, 12.6996172269185, 
    12.8230729897817, 12.5431199073792, 12.2545596758525, 11.8099154559049, 
    16.7619681888156, 16.6501060061985, 16.6135035620795, 16.5191546546088, 
    16.3023495144314, 16.1949738396539, 15.6564608679877, 15.0288678275214, 
    14.5090747409397, 14.2524926927355, 14.2437662548489, 14.2262574301826, 
    14.2550700505575, 14.0618057250977, 13.6228618621826, 13.2174592547947, 
    13.3244410620795, 13.5286852518717, 13.0062580903371, 12.7373469670614, 
    12.8005523681641, 12.5572541554769, 12.4020782311757, 12.0418565273285, 
    16.7299904293484, 16.6391531626383, 16.5906564924452, 16.4295488993327, 
    16.1397125456068, 15.9153903325399, 14.9179495705499, 14.4562714894613, 
    14.2276825375027, 14.0060107972887, 14.2044010162354, 14.1288526323107, 
    14.2445563210381, 14.0602705213759, 13.5728641086155, 13.2653001149495, 
    13.2593864864773, 13.3914142184787, 12.9605952368842, 13.0803106096056, 
    12.95032787323, 12.4206313027276, 16.6830965677897, 16.605015012953, 
    16.5303145514594, 16.261223687066, 15.8899359173245, 15.5614006254408, 
    14.3891898261176, 14.2678381601969, 14.1427737341987, 14.0319456524319, 
    14.2769354714288, 14.1349148220486, 14.1219362682766, 14.0160848829481, 
    13.4087260564168, 13.2726073794895, 13.2335738076104, 13.4217456181844, 
    13.3300819396973, 12.8728590806325, 12.6099591255188, 11.7611373901367, 
    16.5453073713515, 16.6594751146105, 16.504063712226, 16.1471852196587, 
    15.7476727167765, 14.9186386532254, 14.2192540698581, 14.2322626113892, 
    14.1901455985175, 14.1077641381158, 14.2853445476956, 14.2372908062405, 
    13.9810821745131, 13.652629216512, 13.3071416219076, 13.1505865520901, 
    13.3366417355008, 13.3675328890483, 13.2597035566966, 12.7523018230091, 
    16.4850802951389, 16.7009355756972, 16.597372478909, 16.4319118923611, 
    15.7308297687107, 15.0302744971381, 14.3462080425686, 14.3078046374851, 
    14.2378835678101, 14.2541847229004, 14.3674765692817, 14.1940219667223, 
    13.9387115902371, 13.4876976013184, 13.3458997938368, 13.3540137608846, 
    13.3433936436971, 13.0555456876755, 12.7493443489075, 16.3583819071452, 
    16.6582137213813, 16.6750068664551, 16.6297707027859, 16.2797036700779, 
    15.6099002626207, 14.688078350491, 14.5009901258681, 14.3117105695936, 
    14.2169443766276, 14.2467801835802, 14.1134147644043, 14.1093176735772, 
    13.8649740219116, 13.7368135452271, 13.5462412304348, 13.1887452602386, 
    16.1676298777262, 16.1829718483819, 16.4308105044895, 16.5501015981038, 
    16.573269950019, 16.4100894927979, 15.6922904120551, 15.0853894551595, 
    14.4374317593045, 14.2810617023044, 13.9479375415378, 13.7754980723063, 
    13.6865578757392, 13.6298183865017, 13.5630769729614, 13.287286567688, 
    16.1440082126194, 15.9405457178752, 16.1725900438097, 16.4159437815348, 
    16.5625470479329, 16.5255928039551, 16.170125219557, 15.4327919218275, 
    14.7020237180922, 14.5902191797892, 14.023085170322, 13.4801154666477, 
    13.3690653906928, 13.3497232860989, 13.1888695822822, 16.2841705746121, 
    15.991359922621, 15.7365686628554, 16.2172402275933, 16.4982920752631, 
    16.4266986846924, 16.2690940433078, 15.7190099292331, 15.2130666308933, 
    14.4114251666599, 13.792090733846, 13.491589334276, 13.1007482210795, 
    13.0359231630961, 16.3576833936903, 16.2014168633355, 15.7058262295193, 
    15.92268731859, 16.3095866309272, 16.1635761260986, 15.9240901735094, 
    15.4498772091336, 14.9578783247206, 14.1020731396145, 13.4668126106262, 
    13.5386196772257, 16.3922928704156, 16.1941201951769, 15.7281476126777, 
    15.588354534573, 15.6562995910645, 15.4005977842543, 14.9456764856974, 
    14.5571029451158, 14.4692549175686, 13.790209558275, 13.5639472007751, 
    13.6707068549262, 16.3683717515733, 16.1618849436442, 15.706549220615, 
    15.5398908191257, 15.2471912172106, 15.008531888326, 14.8845717112223, 
    14.2954171498617, 14.186283853319, 13.6932436625163, 13.7802093823751, 
    13.5170142915514, 16.2615411546495, 16.0834242502848, 15.6941484875149, 
    15.6018696890937, 15.6059975094265, 15.591246287028, 14.6508352491591, 
    14.1529490152995, 13.8686939875285, 13.7975871827867, 13.9659023284912, 
    16.2397570080227, 15.9259145524767, 15.6842571894328, 15.7019195556641, 
    15.767831908332, 15.6611891852485, 14.3862484825982, 14.4069890975952, 
    14.1475509007772, 14.048377778795, 14.0315143267314, 16.093297428555, 
    15.6071000629001, 15.6697368621826, 15.8300728268094, 15.7446065478855, 
    15.4587413999769, 14.7541980743408, 14.6405990388658, 14.4917744530572, 
    14.4027310477363, 14.2200627326965, 15.7957474390666, 15.479488796658, 
    15.4125658671061, 15.6371079550849, 15.1254260804918, 15.0618999269274, 
    15.0161162482368, 14.9064904318915, 14.8707484006882, 14.5494068463643, 
    15.6825097401937, 15.4692361619737, 15.3576439751519, 15.2585238350762, 
    15.0796634886, 15.1348473230998, 14.9781494140625, 15.0079839494493, 
    15.0627092785305, 15.9849858813816, 15.7069696850247, 15.4619029362996, 
    15.2038567860921, 15.2228181627062, 15.2203339470757, 15.061680369907, 
    15.1132759518094, 14.9453402757645, 16.3220885594686, 16.1109341515435, 
    15.9966684977214, 15.5056640836928, 15.4451687071058, 14.9691705703735, 
    14.8884754180908, 14.8138809204102, 16.5040844811334, 16.2422099643283, 
    15.9943749109904, 15.3377110163371, 14.9511218600803, 16.1232522328695, 
    15.9359462526109, 15.467033068339, 14.8854451179504, 13.5994353294373, 
    13.5979795455933, 13.5995578765869, 13.5986251831055, 9.31532955169678, 
    8.70725421905518, 8.33609848022461, 7.74068880081177, 6.13158750534058, 
    5.19000482559204, 4.59018754959106, 4.12346506118774, 3.58884763717651, 
    3.06718969345093, 2.74898195266724, 2.37187910079956, 2.04651880264282, 
    12.3035481770833, 6.71296739578247, 32.5345001220703, 32.5349998474121, 
    32.5349998474121, 32.5354995727539, 32.9124008178711, 33.6688003540039, 
    33.9573997497559, 34.0235992431641, 34.0849990844727, 34.1889991760254, 
    34.298999786377, 34.3860015869141, 34.4630012512207, 34.4879989624023, 
    34.5289993286133, 34.5589981079102, 34.5810012817383, 32.5649998982747, 
    34.0623334248861, 12.7304906845093, 12.7311878204346, 12.7328443527222, 
    12.72651720047, 11.7412452697754, 8.79164543151856, 7.69488296508789, 
    7.55984725952148, 7.06394948959351, 6.39525003433228, 5.37227010726929, 
    4.68950748443604, 4.17570924758911, 3.81572961807251, 3.30136156082153, 
    2.90579581260681, 2.54541397094727, 2.28822183609009, 2.04689741134644, 
    1.84791898727417, 32.5050010681152, 32.5050010681152, 32.5040016174316, 
    32.5034999847412, 32.5343335469564, 32.823600769043, 33.4916000366211, 
    33.8880004882812, 33.9651992797852, 33.9822006225586, 34.0699996948242, 
    34.1269989013672, 34.2529983520508, 34.3610000610352, 34.4519996643066, 
    34.4970016479492, 34.5349998474121, 34.560001373291, 34.5830001831055, 
    34.6030006408691, 17.6937446594238, 17.730001449585, 17.9029378890991, 
    17.4762090047201, 17.0930430094401, 16.9600601196289, 16.7098439534505, 
    16.5314207077026, 16.6710096995036, 16.526294708252, 16.3527167638143, 
    16.3751169840495, 16.0161083539327, 15.5816133817037, 15.2764863967896, 
    14.8742070198059, 14.4290722211202, 14.3898981412252, 13.8408015569051, 
    13.6516863505046, 13.1773961385091, 13.2379206021627, 13.1906150182088, 
    13.4185662269592, 13.3045722643534, 13.426969687144, 13.8271678288778, 
    12.6630237897237, 12.6465126673381, 12.4903418223063, 11.7005270322164, 
    11.6904576619466, 11.4702774683634, 11.1652231216431, 10.91193262736, 
    10.747181892395, 10.5829645792643, 10.586002667745, 10.5524668693542, 
    10.8295833269755, 10.9150748252869, 10.7833188374837, 10.9186166127523, 
    10.6432709693909, 10.5113304456075, 10.2855242093404, 10.1239002545675, 
    9.7872314453125, 9.7298747698466, 9.59417994817098, 9.1812268892924, 
    17.8198748694526, 17.6392057206896, 17.5643804338243, 17.5420337253147, 
    17.0952847798665, 16.8775628407796, 16.6725476582845, 16.5505373213026, 
    16.5457897186279, 16.4281154208713, 16.343317243788, 16.3123306698269, 
    16.1716673109267, 15.6803780661689, 15.5035287009345, 15.1462027231852, 
    14.5049866570367, 14.5207765897115, 14.2151068051656, 13.8870411713918, 
    13.5750086307526, 13.5723111629486, 13.5509833494822, 13.4924126466115, 
    13.5302048524221, 13.5381878217061, 13.4089523156484, 12.5501164595286, 
    12.3746281464895, 12.2436544895172, 11.954217672348, 11.7154717445374, 
    11.490690946579, 11.5040876865387, 11.0936754544576, 10.8819674650828, 
    10.6620230674744, 10.7876935005188, 10.8478193283081, 10.9172400633494, 
    10.8042500019073, 10.8612916469574, 10.8216832478841, 10.6228350798289, 
    10.3714328606923, 10.3506693840027, 10.0106611251831, 9.81047145525614, 
    9.44192910194397, 9.50626516342163, 9.41678277651469, 17.5836211310493, 
    17.4016123877631, 17.3076881832547, 17.2938783433702, 17.0205296410455, 
    16.5892908308241, 16.444886525472, 16.4671819474962, 16.4605950249566, 
    16.3788876003689, 16.358287387424, 16.2349806891547, 16.3441537221273, 
    15.967924118042, 15.6431670718723, 15.106320699056, 14.8781006071303, 
    14.8887236913045, 14.7658449014028, 14.3005955219269, 13.992699543635, 
    13.8920055230459, 13.9328811168671, 13.8702554702759, 13.563724120458, 
    13.3598176638285, 13.1823342641195, 12.3871296246847, 12.4543976783752, 
    12.3695323467255, 12.1202133496602, 11.8451909224192, 11.7435890038808, 
    11.7068467140198, 11.1854019959768, 11.100014368693, 11.0835076967875, 
    11.0870052178701, 11.290478626887, 11.2015292644501, 10.602162361145, 
    10.6968416372935, 10.5739465554555, 10.5508950551351, 10.2892010211945, 
    10.0159233411153, 9.88308580716451, 9.47754645347595, 9.54642979303996, 
    9.60847687721252, 9.59736084938049, 17.8578737046983, 17.4757580227322, 
    17.3423444959852, 17.136117723253, 16.8266557057699, 16.4237306382921, 
    16.2261781692505, 16.3233759138319, 16.3644104003906, 16.4055105845133, 
    16.2233325110541, 16.1807969411214, 16.2578639984131, 15.9792802598741, 
    15.5553878148397, 15.4405717849731, 15.1334377924601, 15.018320719401, 
    14.1424502266778, 13.5896589491102, 13.6089785893758, 14.0257547166612, 
    13.7773008346558, 13.6662279764811, 13.5769941541884, 13.2475368711683, 
    12.8621546427409, 12.1886682510376, 12.1545068952772, 11.7826271057129, 
    11.4144153594971, 11.2593588299221, 11.4101370705499, 11.8091465632121, 
    11.2342240015666, 11.3353686862522, 11.0408602820502, 11.5133555730184, 
    11.5053944057888, 10.8783693313599, 10.9018621444702, 10.7666864395142, 
    10.5701333151923, 10.2417536841498, 10.0768080817329, 9.78638490041097, 
    9.40688652462429, 9.40613248613146, 9.59667587280273, 9.64232455359565, 
    9.70053556230333, 18.0488764444987, 17.6874226464166, 17.2139708201091, 
    16.7603969573975, 16.5977562798394, 16.5083401997884, 15.9480610953437, 
    16.1968622207642, 16.2883911132812, 16.2963922288683, 16.1492309570312, 
    16.238774617513, 16.1791896820068, 15.8920379214817, 15.6881240208944, 
    15.512035369873, 15.2317394680447, 14.3131673336029, 13.3686785697937, 
    13.0937016010284, 13.1980386575063, 13.5436470508575, 13.6028870741526, 
    13.6169222195943, 13.3935787677765, 12.8424541950226, 12.4858194986979, 
    12.1658274332682, 11.6716759204865, 11.2865296999613, 11.1014885107676, 
    10.9867877960205, 10.9677430788676, 11.1730676492055, 11.2838368415833, 
    11.2536792755127, 10.9494264125824, 11.0426816940308, 11.1063735485077, 
    10.8888674577077, 10.8158638477325, 10.4961854616801, 10.2884578704834, 
    9.84350482622782, 9.5776302019755, 9.37283190091451, 9.34943087895711, 
    9.41421914100647, 9.58926304181417, 9.63160339991252, 9.64310669898987, 
    17.7513412899441, 17.5036349826389, 17.0402200486925, 16.8896609412299, 
    16.7908520168728, 16.6004967159695, 16.1334100299411, 16.2982090844048, 
    16.2104697757297, 16.124932607015, 16.0962270100911, 16.0330641004774, 
    16.0026455985175, 15.6726339128282, 15.5646432240804, 15.1958654191759, 
    14.5252039167616, 13.5518030325572, 13.0654783248901, 12.937236626943, 
    13.1541740894318, 13.4190465609233, 13.46657594045, 13.5723748207092, 
    13.3312193552653, 12.5441193580627, 12.232275724411, 11.79958264033, 
    11.2710422674815, 11.209298213323, 11.0212182998657, 11.0891395409902, 
    10.7412243684133, 10.9143273830414, 11.004249493281, 11.1027876536051, 
    10.9007859230042, 10.8055682182312, 10.8819371859233, 10.7995351950328, 
    10.7382980982463, 10.328110853831, 9.85271469751994, 9.7894766330719, 
    9.698619445165, 9.43217730522156, 9.41277432441711, 9.49573953946432, 
    9.66675964991252, 9.64011073112488, 9.58169007301331, 17.6035073598226, 
    17.5943400065104, 17.3976018693712, 16.8465008205838, 16.9019198947483, 
    16.6852887471517, 16.191753493415, 16.2127687666151, 15.9862818188137, 
    15.8714865578545, 15.8788563410441, 15.9447668923272, 15.5844176610311, 
    15.4065341949463, 15.3983361985948, 15.0272776285807, 13.7392331229316, 
    13.0319796668159, 12.9851797951592, 13.159310552809, 13.3343562020196, 
    13.3898849487305, 13.5241437488132, 13.4872890048557, 13.2164336310493, 
    12.5225928624471, 11.7971421347724, 11.2028819190131, 11.0694305631849, 
    11.1828544404772, 11.1338216993544, 11.1642991171943, 10.9823678334554, 
    10.6853509479099, 10.6373866399129, 10.6441168255276, 10.6786989635891, 
    10.7393777635362, 10.8137979507446, 10.881268925137, 10.6596859825982, 
    10.1933857599894, 9.86532274881999, 9.92752022213406, 9.92485374874539, 
    9.75587452782525, 9.58518674638536, 9.6163420147366, 9.5298408932156, 
    9.55176226298014, 9.59445646074083, 17.8232216305203, 17.7993960910373, 
    17.4004737006293, 16.9378689659966, 16.8744475046794, 16.6244667900933, 
    16.2127684487237, 16.1646341747708, 15.6907200283474, 15.7386397255792, 
    15.8974473741319, 15.7422457800971, 15.5820118586222, 15.4756342569987, 
    15.0400630103217, 14.5560195710924, 13.2131905025906, 12.8973366419474, 
    13.1204452514648, 13.2991565068563, 13.4008554617564, 13.3070964813232, 
    13.3286213080088, 13.1996954282125, 13.053169965744, 12.2082912127177, 
    11.3724638621012, 11.0728227297465, 11.1757430235545, 11.1569720109304, 
    11.1440397898356, 11.1022510528564, 11.1525371869405, 10.7519336541494, 
    10.537723382314, 10.5064031283061, 10.7146492799123, 10.7242278258006, 
    10.606997013092, 11.0008883476257, 10.8405505021413, 10.665420850118, 
    10.175589799881, 9.94765988985697, 10.0212404727936, 9.86375157038371, 
    9.66036359469096, 9.64508748054504, 9.30817635854085, 9.48144205411275, 
    9.91018295288086, 17.9198691050212, 17.6129336886936, 17.6962846120199, 
    17.1957715352376, 17.0172687106662, 16.5033164554172, 16.2304840087891, 
    16.1439954969618, 15.8119518491957, 15.8972210354275, 15.70753426022, 
    14.8973132239448, 15.0877508587307, 15.2614866892497, 15.0096100701226, 
    14.0767629411485, 13.0367517471313, 12.7686416308085, 13.1524867216746, 
    13.4040497144063, 13.381637096405, 13.3032680352529, 13.3224405447642, 
    13.3534615039825, 12.8783390522003, 11.804424683253, 11.1811677614848, 
    11.0586311022441, 11.3020377159119, 11.3470168908437, 11.2274162769318, 
    11.1118377049764, 11.1096940835317, 10.842182079951, 10.6069476604462, 
    10.8009316126506, 10.552343527476, 10.4983580907186, 10.6097234884898, 
    10.8122088909149, 10.9093942642212, 10.68412510554, 10.2358697255452, 
    10.0641175111135, 9.99645884831746, 9.8703285853068, 9.74492979049683, 
    9.42668867111206, 9.14692068099976, 9.47405815124512, 10.0737017790476, 
    17.8784493340386, 17.725341796875, 17.5648905436198, 17.2703062693278, 
    16.694860458374, 16.2659132215712, 16.3099185095893, 16.2484171125624, 
    16.0808562172784, 15.795166015625, 14.9516269895766, 14.6167897118462, 
    14.6110917197333, 15.1670979393853, 15.0547364552816, 13.788050227695, 
    13.0440475675795, 12.5728293524848, 12.9914990531074, 13.3674942652384, 
    13.3184143702189, 13.2921698888143, 13.175066947937, 13.0230136447483, 
    12.6941702100966, 11.6363002989027, 11.0365765889486, 11.0892339282566, 
    11.3495619032118, 11.4744086795383, 11.1871983210246, 11.1445175806681, 
    11.1997865041097, 10.767770131429, 10.6248502731323, 10.5768300162421, 
    10.5051353242662, 10.4831972122192, 10.6759746339586, 10.84071720971, 
    10.9569389555189, 10.5881834030151, 10.3544262780084, 10.3075529734294, 
    9.92250156402588, 9.79712581634521, 9.97758928934733, 9.52689711252848, 
    9.30525557200114, 9.90899011823866, 9.98599296145969, 17.8575579325358, 
    17.5838911268446, 17.5293602413601, 17.1865906185574, 17.177942276001, 
    16.6429621378581, 16.4565052456326, 16.3173242145114, 15.8799634509616, 
    15.4684620963203, 14.7323178185357, 14.6386131710476, 14.3932049009535, 
    14.4424351586236, 14.589706103007, 13.4534349441528, 13.1558331383599, 
    12.6311225891113, 12.5563387870789, 12.9378110567729, 13.1962159474691, 
    13.1397460301717, 13.0272949536641, 12.8885877927144, 12.6423428853353, 
    11.6248348553975, 11.0736499627431, 11.1259814898173, 11.4179697036743, 
    11.6311333179474, 11.3230783939362, 11.5112370649974, 11.2563999493917, 
    11.0130527814229, 10.7334837118785, 10.672067006429, 10.5905209382375, 
    10.5231002966563, 10.9278486569722, 10.6903898715973, 10.4878570238749, 
    10.3676682313283, 10.353929678599, 10.2997822761536, 10.0132249991099, 
    9.90369002024333, 9.89982096354167, 9.60605986913045, 9.69349964459737, 
    10.1795384089152, 9.95627236366272, 17.4917736053467, 17.4664827982585, 
    17.427858988444, 17.3796819051107, 17.4359192318386, 17.1134018368191, 
    16.8423716227214, 16.2502483791775, 15.6992734273275, 15.1520607206557, 
    14.5940441555447, 14.5505153867933, 14.302891837226, 14.0680945714315, 
    13.9383125305176, 13.2382972505358, 13.1347823672824, 12.6253323554993, 
    12.5671638647715, 12.5567539532979, 13.0168108145396, 12.9289659659068, 
    12.8320221106211, 12.8042879899343, 12.491091410319, 11.7960019906362, 
    11.2173762321472, 11.4647114276886, 11.9478599230448, 12.2364477316538, 
    11.2483568986257, 11.3553188641866, 11.3606896400452, 11.1350758075714, 
    10.965448141098, 10.7341481844584, 10.7847356001536, 10.6277194023132, 
    10.8504501183828, 10.6708690325419, 10.4891974131266, 10.3830798467, 
    10.3069052696228, 10.2867267926534, 9.99286468823751, 9.89801359176636, 
    9.98685932159424, 9.39051556587219, 10.1737484137217, 10.2835642496745, 
    10.0157055854797, 17.1913159688314, 17.3917713165283, 17.2457093132867, 
    17.288361231486, 17.3820669386122, 17.1072118547228, 16.7282307942708, 
    16.1454696655273, 15.5512924194336, 14.815819952223, 14.5415954589844, 
    14.5863242679172, 14.2200298309326, 14.230518023173, 14.0888669755724, 
    13.3389869266086, 13.1271486282349, 12.7360253863864, 12.9757295184665, 
    12.7225756115384, 12.7328098085192, 12.8271376291911, 12.6503926383124, 
    12.6276279025608, 12.3777878019545, 12.1371737586127, 11.7804435094198, 
    12.094886885749, 12.3164033889771, 12.221930609809, 11.1599800321791, 
    10.9656209945679, 11.174190097385, 10.9967477586534, 11.1361507839627, 
    10.732189072503, 11.0445665783352, 10.9317961798774, 11.0215794245402, 
    10.9545832739936, 10.6683674918281, 10.4168854819404, 10.4643559985691, 
    10.1686414082845, 9.97388044993083, 10.041015625, 9.90664037068685, 
    9.69203588697645, 10.3209598329332, 10.1847699483236, 9.81614759233263, 
    16.9579802619086, 17.2916526794434, 17.2281307644314, 17.4965534210205, 
    17.4044592115614, 17.1574242909749, 16.4474059210883, 16.1636621687147, 
    15.7707703908285, 14.8302983178033, 14.627046585083, 14.648770014445, 
    14.1851296954685, 14.2288015153673, 14.2114686965942, 13.5477084053887, 
    13.1695155037774, 12.8259863853455, 13.2424849669139, 12.953651825587, 
    12.5603220462799, 12.5214128494263, 12.5291795730591, 12.701931476593, 
    12.7497297128042, 12.720405737559, 12.4349336624146, 11.6567958990733, 
    11.7119430700938, 11.5628360112508, 11.086980899175, 10.9215311209361, 
    10.7400667667389, 10.9284597237905, 10.7274704846469, 10.6769940853119, 
    9.99999986376081, 10.1999998092651, 10.3875000476837, 10.533749961853, 
    10.428658246994, 10.3270554542542, 10.8476403554281, 10.3791363579886, 
    9.9888870716095, 9.83368062973022, 9.34434620539347, 9.67870911684903, 
    10.1049786567688, 9.86479715867476, 9.54644044240316, 16.8101618025038, 
    16.8340515560574, 16.8954230414497, 17.0987381405301, 17.0843221876356, 
    16.6996739705404, 16.4336982303196, 15.9715741475423, 15.8004233042399, 
    15.0859494739109, 14.532747692532, 14.5420604281955, 14.2711844974094, 
    14.2711011038886, 14.2851909001668, 13.6191870371501, 13.3917134602865, 
    12.9598387082418, 13.2413777510325, 13.1666126251221, 12.5602582295736, 
    12.3210634390513, 12.362070719401, 12.4999029636383, 12.8081270853678, 
    12.8076260884603, 12.1857833067576, 11.3487754662832, 11.3504402637482, 
    11.2916509310404, 11.2155196666718, 10.9667645295461, 10.8280895551046, 
    11.1761148626154, 10.672611951828, 10.5407814184825, 10.1969999313354, 
    10.2910714830671, 10.197500038147, 10.375, 10.2679562568665, 
    10.2842186689377, 9.23125004768372, 9.44553579602923, 9.60299987792969, 
    9.40031266212463, 9.75086291631063, 9.67499987284342, 9.70499992370605, 
    16.8869599236382, 16.7085613674588, 16.6881190405952, 16.7675493028429, 
    16.9711772070991, 16.7388899061415, 16.5291025373671, 16.2812351650662, 
    15.8937301635742, 15.1891639497545, 14.7872800827026, 14.5336057874891, 
    14.1863159603543, 14.3047397401598, 14.2858152389526, 13.7970335218641, 
    13.4382271236844, 13.2771546045939, 13.34112962087, 13.2800630993313, 
    12.7100060780843, 12.4916163550483, 12.2745282914903, 12.4712777667575, 
    12.721126238505, 12.8023256725735, 11.7744862238566, 11.2545075946384, 
    11.5732632742988, 11.6051670710246, 11.3573787477281, 10.5458994971381, 
    10.8525001525879, 11.2906250423855, 10.8532552719116, 10.6052098274231, 
    10.3124081747872, 10.0362501144409, 11.0500001907349, 10.2791666984558, 
    10.3552083969116, 9.75, 10.1999998092651, 9.75749988555908, 
    9.70666631062826, 9.76518938276503, 9.78986114925808, 10.1500220828586, 
    9.88437521457672, 9.82392480638292, 9.77708339691162, 16.8460528055827, 
    16.6969028049045, 16.6693053775364, 16.6027007632785, 16.8233432769775, 
    16.4415020412869, 16.0996532440186, 16.230062590705, 16.2292363908556, 
    15.3381661309136, 14.9258574379815, 14.3943520651923, 14.0936975479126, 
    14.3146342171563, 14.4334565268623, 14.0916333728366, 13.6051068835788, 
    13.432475010554, 13.4415332476298, 13.2520198822021, 12.749720176061, 
    12.5567207336426, 12.3796145121257, 12.2824199994405, 12.4724773565928, 
    12.6209418773651, 11.5978225866954, 11.2709999879201, 11.7634595235189, 
    11.7419753869375, 11.3050923877292, 11.4008680184682, 11.0583333969116, 
    11.1414774114435, 10.8548458947076, 9.69999994550433, 9.99892861502511, 
    10.1999998092651, 10.3078126907349, 9.95000004768372, 9.61514854431152, 
    9.58363395267063, 9.91185609499613, 9.77400024731954, 9.18947919209798, 
    9.72964421908061, 9.82457224527995, 9.37186543146769, 16.9208236270481, 
    16.6820299360487, 16.5760112338596, 16.4555568695068, 16.3555111355252, 
    16.1306425730387, 16.0809540218777, 16.3536508348253, 16.5325609842936, 
    15.6816308763292, 15.2450415293376, 14.1262573666043, 13.9475469589233, 
    14.0432411829631, 13.9594891866048, 13.8594152662489, 13.7654229270087, 
    13.6826733748118, 13.4467675685883, 13.3324186007182, 12.8468386332194, 
    12.4868791898092, 12.472663640976, 12.5351433753967, 12.6020941734314, 
    12.4170015652974, 11.8058098951975, 11.5054933230082, 11.5939283370972, 
    10.8580003738403, 11.6250001192093, 11.1625001213767, 10.8682735988072, 
    9.87142876216343, 9.09999990463257, 10.483333269755, 9.8746874332428, 
    9.73693171414462, 9.60545444488525, 9.44629796346029, 8.29400690396627, 
    8.50310778617859, 8.63380159031261, 8.3155323266983, 16.9304105970595, 
    16.7285346984863, 16.718334197998, 16.3896410200331, 16.1789390775892, 
    16.1237291759915, 15.8911561965942, 16.1852672364977, 16.0732000139025, 
    15.7409620285034, 15.2056303024292, 14.1742097006904, 13.7991377512614, 
    13.7555203967624, 13.6778740353054, 13.6212106280857, 13.7321102354262, 
    13.7196203867594, 13.1563532087538, 13.0029147466024, 12.8011322021484, 
    12.4927955203586, 12.3390264511108, 12.2767884996202, 11.9908799065484, 
    11.9892830318875, 11.7705237070719, 11.604575475057, 8.24499979019165, 
    8.83703136444092, 8.65571673711141, 8.13243993123372, 16.9150602552626, 
    16.8731257120768, 16.7148259480794, 16.4834679497613, 16.3424186706543, 
    16.1645090315077, 16.1189714007907, 16.0495785607232, 15.8201479381985, 
    15.2510902616713, 14.5936047236125, 14.1666332880656, 14.0119410620795, 
    13.8103545506795, 13.5956364737617, 13.3327444924249, 13.5320729149712, 
    13.6787450313568, 13.1607396602631, 12.8429358800252, 12.6888354619344, 
    12.8184821605682, 12.5547772248586, 12.2545596758525, 11.8099154559049, 
    16.6500432756212, 16.5723567538791, 16.5567027197944, 16.4666697184245, 
    16.2542209625244, 16.1898556815253, 15.6560639275445, 14.9813301298353, 
    14.5080601374308, 14.2438420189752, 14.205491065979, 14.1945614284939, 
    14.2472356160482, 14.0375741322835, 13.5961010191176, 13.1873145633274, 
    13.3213895161947, 13.5384578704834, 13.0494287014008, 12.7496828238169, 
    12.7807025114695, 12.5487875143687, 12.4100335439046, 12.0418565273285, 
    16.7167063819038, 16.6062689887153, 16.5582692888048, 16.390574561225, 
    16.1514792972141, 15.9296471277873, 14.8804454803467, 14.4534637663099, 
    14.2308008405897, 14.0397000842624, 14.227807574802, 14.1478486590915, 
    14.222783724467, 14.0418914159139, 13.544380929735, 13.2363941404555, 
    13.2634728749593, 13.4129254023234, 12.9704467985365, 13.0891261630588, 
    12.9389547771878, 12.4134928385417, 16.7234944237603, 16.6337297227648, 
    16.5562148623996, 16.251942952474, 15.9043377770318, 15.5893025928073, 
    14.388891643948, 14.289000193278, 14.1575982835558, 14.0553369522095, 
    14.2832481596205, 14.1568938361274, 14.1120427449544, 14.0046656926473, 
    13.3942487504747, 13.2395684983995, 13.2389114167955, 13.4611438115438, 
    13.3420360883077, 12.8663490613302, 12.5922852357229, 11.767521572113, 
    16.5187507205539, 16.6738529205322, 16.5254272884793, 16.1311232248942, 
    15.705591307746, 14.8826036453247, 14.2167616950141, 14.2471878263685, 
    14.2252396477593, 14.1434471342299, 14.3034642537435, 14.2403863271077, 
    13.9984793133206, 13.660028245714, 13.302926381429, 13.1349129147, 
    13.3327792485555, 13.3654622236888, 13.254326581955, 12.7463287006725, 
    16.4282684326172, 16.7031091054281, 16.6201962365044, 16.3743000030518, 
    15.7320693333944, 14.9624101850722, 14.3652086257935, 14.3763501909044, 
    14.2819900512695, 14.2773803075155, 14.357508553399, 14.1819967693753, 
    13.9337762196859, 13.5071983337402, 13.3438786400689, 13.3531330956353, 
    13.3523423936632, 13.0436960458755, 12.7420965433121, 16.3700389862061, 
    16.6647330390082, 16.6897926330566, 16.6506565941705, 16.230073928833, 
    15.5506753921509, 14.8662859598796, 14.6224585639106, 14.4423459370931, 
    14.3043140835232, 14.2257910834418, 14.1017989052667, 14.0819370481703, 
    13.8633456759983, 13.7263580958048, 13.5428926679823, 13.1832609176636, 
    16.1560103098551, 16.1870237986247, 16.4139876895481, 16.5496135287815, 
    16.597290886773, 16.4025463528103, 15.7143149905735, 15.2816406885783, 
    14.548161400689, 14.4151511722141, 14.0122577879164, 13.7738244798448, 
    13.6713432735867, 13.6146290037367, 13.5428795284695, 13.2911334991455, 
    16.1948632134332, 15.9619491365221, 16.1278898451063, 16.4467860327827, 
    16.5890375773112, 16.6035957336426, 16.190395143297, 15.6050075954861, 
    14.7484658559163, 14.6686903635661, 14.1396536297268, 13.4697051578098, 
    13.3605552249485, 13.3454692628649, 13.1741477118598, 16.3400446573893, 
    16.0223497814602, 15.7546922895643, 16.2794257269965, 16.5503819783529, 
    16.4987733629015, 16.3173364003499, 15.8189455668132, 15.2600491841634, 
    14.4556562635634, 13.8633808559842, 13.4991920259264, 13.096159140269, 
    13.0249026616414, 16.370738559299, 16.2104663848877, 15.7471460766262, 
    16.0429756376478, 16.3412776523166, 16.1532973183526, 15.8721218109131, 
    15.4567687776354, 15.0524798499213, 14.1434533860948, 13.4882436990738, 
    13.5612008836534, 16.4268656836616, 16.2122660742866, 15.7546354929606, 
    15.6148114734226, 15.6239806281196, 15.3284576204088, 14.9734172821045, 
    14.699456108941, 14.6190871132745, 13.9916317198012, 13.6137543916702, 
    13.6740821202596, 16.399057176378, 16.2187564637926, 15.7605288823446, 
    15.565821117825, 15.2564761903551, 15.0411933263143, 14.8318073484633, 
    14.3370991812812, 14.254535039266, 13.741199069553, 13.8378376960754, 
    13.5181556277805, 16.2690987057156, 16.0941608217027, 15.7425896326701, 
    15.6051549911499, 15.6006045871311, 15.5933791266547, 14.6668214797974, 
    14.3171984354655, 14.0433803134494, 13.9103853437636, 14.006888601515, 
    16.2057395511203, 15.8962050543891, 15.7133515675863, 15.718627081977, 
    15.767907778422, 15.7143564224243, 14.4076065487332, 14.4246826171875, 
    14.2096020380656, 14.1505030526055, 14.1717019081116, 16.0270653830634, 
    15.5376519097222, 15.7218840916952, 15.859214146932, 15.7409678565131, 
    15.4992487165663, 14.79220061832, 14.6972401936849, 14.540459950765, 
    14.4677571190728, 14.2809767723083, 15.7460888756646, 15.4975696139865, 
    15.4366044998169, 15.6886438793606, 15.1006814108955, 15.0863129297892, 
    15.0219135284424, 14.9261100557115, 14.89275431633, 14.6215642293294, 
    15.6736613379584, 15.5040584140354, 15.3619737625122, 15.3058924145169, 
    15.091618431939, 15.1621013217502, 15.0464191436768, 15.018789185418, 
    15.0707364612155, 15.9488146040175, 15.7705305947198, 15.5051981608073, 
    15.2187773386637, 15.2492617501153, 15.2279349433051, 15.1302349302504, 
    15.1409287982517, 14.9575517177582, 16.3364404042562, 16.1462031470405, 
    16.0858464770847, 15.5420289569431, 15.5157400767008, 14.9886971579658, 
    14.8799578802926, 14.7411727905273, 16.5501147376166, 16.2896082136366, 
    16.0546145968967, 15.3607108857897, 14.9214821921455, 16.1607813305325, 
    15.9212759865655, 15.5850780275133, 14.9529047012329, 13.660737991333, 
    13.6543226242065, 13.6519346237183, 13.6475734710693, 13.5557880401611, 
    12.320969581604, 10.9682931900024, 9.3370189666748, 9.09381484985352, 
    8.71106433868408, 7.90615367889404, 7.44208955764771, 6.51879835128784, 
    6.36768102645874, 5.95759439468384, 5.44174098968506, 5.31588220596313, 
    5.07773685455322, 4.81876945495605, 4.48915863037109, 4.3190770149231, 
    4.09442853927612, 3.94832134246826, 33.0390014648438, 33.0410003662109, 
    33.0419998168945, 33.0429992675781, 33.0460014343262, 33.1069984436035, 
    33.4220008850098, 33.6570014953613, 33.9179992675781, 34.0260009765625, 
    34.0579986572266, 34.1319999694824, 34.1189994812012, 34.226001739502, 
    34.2350006103516, 34.306999206543, 34.3440017700195, 34.3549995422363, 
    34.3779983520508, 34.4150009155273, 34.4290008544922, 34.4309997558594, 
    34.4529991149902, 11.9808597564697, 11.979567527771, 11.9672937393188, 
    11.8038272857666, 11.5040793418884, 11.1912132898966, 8.86040439605713, 
    7.94273729324341, 7.68683080673218, 7.27129459381104, 6.4627062479655, 
    5.905433177948, 4.96015405654907, 4.36980199813843, 3.99167037010193, 
    3.61798858642578, 3.20025634765625, 2.93255996704102, 2.66319346427917, 
    2.38115048408508, 2.12302207946777, 2.01422190666199, 1.83520793914795, 
    32.609001159668, 32.6080017089844, 32.6049995422363, 32.5929985046387, 
    32.5665016174316, 32.5890007019043, 32.863200378418, 33.4963996887207, 
    33.8833999633789, 33.9877998352051, 34.0226669311523, 34.0349998474121, 
    34.1080017089844, 34.1699981689453, 34.2569999694824, 34.3660011291504, 
    34.423999786377, 34.4700012207031, 34.5040016174316, 34.5349998474121, 
    34.5610008239746, 34.576000213623, 34.5909996032715, 8.24374903165377, 
    8.07208486703726, 7.40963862492488, 10.1993227005005, 10.1984163920085, 
    10.1972808837891, 10.1961441040039, 9.74515962600708, 8.72219058445522, 
    8.59093364079793, 8.52049914995829, 8.14381901423136, 7.83411924044291, 
    6.89342304070791, 6.35731637477875, 6.05581331253052, 17.4521064758301, 
    17.5186147689819, 17.7798026402791, 17.2524731953939, 16.8908859888713, 
    16.841423034668, 16.6067616144816, 16.4914929072062, 16.4654572804769, 
    16.3707898457845, 16.310320854187, 16.2978836695353, 15.9055972099304, 
    15.5073030789693, 15.2727502187093, 14.7865436871847, 14.3055931727091, 
    14.2342782020569, 13.8623596827189, 13.5598425865173, 13.2206937472026, 
    13.1862414677938, 13.1362455685933, 13.1925018628438, 13.2313092549642, 
    13.3542019526164, 13.3689521153768, 12.9612310727437, 12.3907348314921, 
    11.9085378646851, 11.7606477737427, 11.8396237691243, 11.6014156341553, 
    11.2889803250631, 11.0234769185384, 10.8983608881632, 10.5983700752258, 
    10.7106485366821, 10.7239500681559, 10.8712759017944, 10.4368408521016, 
    10.269420782725, 10.5252105394999, 10.2006138165792, 10.1269243558248, 
    9.92950487136841, 9.83324750264486, 9.70593372980754, 9.47948582967122, 
    9.28510999679565, 8.92641830444336, 17.6219306521946, 17.4285803900825, 
    17.6011778513591, 17.4277763366699, 16.9896969265408, 16.806791305542, 
    16.5446597205268, 16.4778535630968, 16.4132408565945, 16.3403911590576, 
    16.3200971815321, 16.301718182034, 16.0416741900974, 15.5963178210788, 
    15.4450531005859, 14.9978722466363, 14.3880194558038, 14.4419848124186, 
    14.050444761912, 13.7898867925008, 13.550878127416, 13.4420030117035, 
    13.3393286863963, 13.3702449798584, 13.4143737951914, 13.3680259386698, 
    13.3220423857371, 12.8759008248647, 12.3103707631429, 12.0574643611908, 
    11.7251416842143, 11.6445637543996, 11.4323325157166, 11.4365921815236, 
    11.1384031772614, 10.8755568663279, 10.7099364598592, 10.8574593861898, 
    11.0625181992849, 11.0488599141439, 10.765119155248, 10.4057608445485, 
    10.4253056049347, 10.3070116837819, 10.070229212443, 9.99454148610433, 
    9.66588393847148, 9.56306902567546, 9.2147487004598, 9.27773412068685, 
    9.13771017392476, 17.4306439293755, 17.100271013048, 17.2871918148465, 
    17.294442070855, 16.9547742207845, 16.5289906395806, 16.3720082177056, 
    16.4089387257894, 16.343271891276, 16.2679996490479, 16.2781829833984, 
    16.1842695871989, 15.917549027337, 15.7824754714966, 15.5193818410238, 
    15.1113849216037, 14.7047296100193, 14.6815431118011, 14.4707549413045, 
    14.1779828866323, 13.9392410119375, 13.8542853196462, 13.7608026663462, 
    13.7187414169312, 13.6086111863454, 13.287735303243, 13.1619271437327, 
    12.7353624502818, 12.1838668982188, 11.8532002766927, 11.8354760805766, 
    11.7362672487895, 11.7333873907725, 11.5870920022329, 11.2722353935242, 
    11.0725568135579, 10.9285651048025, 11.0542931556702, 11.1458199818929, 
    11.0035116672516, 10.7099262078603, 10.6812395254771, 10.4409442742666, 
    10.2368634541829, 9.98233977953593, 9.76400502522787, 9.53174328804016, 
    9.26571981112162, 9.24029572804769, 9.33757742245992, 9.35421347618103, 
    17.569976594713, 17.2467642890082, 17.290078692966, 17.1035338507758, 
    16.788572523329, 16.3662221696642, 16.2446363237169, 16.2455399831136, 
    16.1274789174398, 16.2404865688748, 16.1693587832981, 16.0955412122938, 
    16.0071778827243, 15.9049780103895, 15.5378581153022, 15.2406288782756, 
    14.9144949383206, 14.8854532241821, 14.1397955152724, 13.6351191202799, 
    13.6026152504815, 14.0081446965535, 13.8747368918525, 13.7173813713921, 
    13.5757745107015, 13.1989316940308, 12.9187299940321, 12.3610553741455, 
    11.7746045854357, 11.4823514090644, 11.4825720257229, 11.4868247773912, 
    11.4990451600817, 11.7097430759006, 11.2997133466933, 11.2384759055244, 
    10.964741812812, 11.0447864532471, 11.0755052566528, 10.8023805618286, 
    10.8496902253893, 10.8572898440891, 10.2761414845785, 9.75024318695068, 
    9.85389433966743, 9.49061563279894, 9.12722259097629, 9.2241399553087, 
    9.19973776075575, 9.32647874620226, 9.29020108116998, 17.8756773206923, 
    17.6297878689236, 17.0689252217611, 16.7287686665853, 16.5870543585883, 
    16.4807275136312, 16.1611103481717, 16.198420630561, 16.1590167151557, 
    16.0821250279744, 16.0825830035739, 16.0507758458455, 15.9843485090468, 
    15.8028156492445, 15.608029683431, 15.3899722629123, 15.121560520596, 
    14.2839774290721, 13.3028551737467, 13.0803511937459, 13.1461062431335, 
    13.4151796499888, 13.5497903029124, 13.5905869801839, 13.4388221899668, 
    12.8800951639811, 12.587162733078, 12.1518103281657, 11.5915264288584, 
    11.3111531734467, 11.095096429189, 11.0714058081309, 11.0993487040202, 
    11.3157296975454, 11.2154105504354, 11.0974852244059, 10.8645830154419, 
    10.8171068032583, 10.8643432458242, 10.7589556376139, 10.4802484512329, 
    10.6074829101562, 10.0276446342468, 9.64030305544535, 9.38900009791056, 
    9.19114589691162, 9.26121393839518, 9.3174409866333, 9.32460363705953, 
    9.28718034426371, 9.28494834899902, 17.460947672526, 17.2921045091417, 
    16.9064945644803, 16.8219634162055, 16.7925391727024, 16.5447442796495, 
    16.2759034898546, 16.1724580128988, 15.9177476035224, 15.9008036719428, 
    15.866995493571, 15.8210973739624, 15.7004843817817, 15.5838333765666, 
    15.5269913143582, 15.1475962532891, 14.5017631318834, 13.5341317653656, 
    12.9784826437632, 12.9189412593842, 13.1180390516917, 13.3457023302714, 
    13.4151781400045, 13.4620412985484, 13.2540368239085, 12.5827696323395, 
    12.2628451188405, 11.7487033208211, 11.3881251811981, 11.2123995621999, 
    11.060887893041, 11.0526096820831, 10.7692728837331, 11.0099306106567, 
    10.8564976851145, 10.7845520178477, 10.6250243186951, 10.7084084351858, 
    10.7724155584971, 10.4239570299784, 10.3792924880981, 10.0790359179179, 
    9.70093472798665, 9.5265306631724, 9.55407087008158, 9.14119784037272, 
    9.26633985837301, 9.46097207069397, 9.31397517522176, 9.11934463183085, 
    9.28313080469767, 17.3682842254639, 17.2471894158257, 16.9193670484755, 
    16.8115914662679, 16.8810886806912, 16.6719301011827, 16.2131411234538, 
    16.1612383524577, 15.795837826199, 15.6934294170803, 15.6967204411825, 
    15.6943811840481, 15.3774884541829, 15.3446379767524, 15.3773932986789, 
    14.9805707931519, 13.7670423719618, 13.0132239659627, 12.9265489578247, 
    13.1503536436293, 13.295097457038, 13.2833137512207, 13.3486553827922, 
    13.4184143278334, 13.0149866739909, 12.3825714323256, 11.7942488988241, 
    11.2635938856337, 11.0550860299004, 11.1337244245741, 11.1229219436646, 
    11.0452704959446, 10.8799964057075, 10.6041901906331, 10.4979076385498, 
    10.3600741492377, 10.5765366024441, 10.5863953696357, 10.4602131313748, 
    10.6872665617201, 10.4889279471503, 10.1740267011854, 9.657593621148, 
    9.80379030439589, 9.77239269680447, 9.59166929456923, 9.33735423617893, 
    9.36344146728516, 9.21082602606879, 9.00909847683377, 9.38681104448107, 
    17.6048810746935, 17.2099829779731, 16.8422730763753, 16.8244101206462, 
    16.8669668833415, 16.6695868174235, 16.177431318495, 16.1357449425591, 
    15.6615494622125, 15.6309589809842, 15.5704087151421, 15.4403504265679, 
    15.3234673606025, 15.2438584433662, 15.1414667765299, 14.4632595909966, 
    13.1980572806464, 12.8490618069967, 13.0770213603973, 13.2958097457886, 
    13.3580228487651, 13.3060825665792, 13.2893598079681, 13.2881183624268, 
    12.780524969101, 12.1601657072703, 11.3866142431895, 11.1056428750356, 
    11.2059735457102, 11.1468830108643, 11.0570120811462, 11.059386809667, 
    10.9563518365224, 10.6054191589355, 10.3788825670878, 10.3714208602905, 
    10.5570543607076, 10.5125839710236, 10.4468135039012, 10.8159352938334, 
    10.6987140973409, 10.4728709856669, 9.88036672274272, 9.73555493354797, 
    9.77897310256958, 9.55955600738525, 9.44276229540507, 9.36133503913879, 
    9.26112524668376, 9.25328882535299, 9.84788568814596, 17.3467415703668, 
    17.0314617156982, 17.1708937750922, 17.0271538628472, 16.8579906887478, 
    16.3788168165419, 16.1856293148465, 16.1105258729723, 15.544707192315, 
    15.6890062756009, 15.185282919142, 14.6420967313978, 15.0363584094577, 
    15.0997334586249, 15.0147565205892, 14.0352684656779, 12.9967965020074, 
    12.7035621007284, 13.1184571584066, 13.318962097168, 13.3493412335714, 
    13.2460509141286, 13.293865998586, 13.2275763352712, 12.7051961421967, 
    11.8372422854106, 11.1144257386525, 11.0139896869659, 11.2271356582642, 
    11.2823483149211, 10.9825354417165, 10.9881097475688, 11.0766909917196, 
    10.6976267496745, 10.3821472326914, 10.285730044047, 10.5012300014496, 
    10.4193830490112, 10.5050875345866, 10.7123951117198, 10.7778221766154, 
    10.5599930286407, 10.0907887617747, 9.78257417678833, 9.8262669245402, 
    9.6224148273468, 9.54590805371602, 9.23143712679545, 9.25817863146464, 
    9.5073143641154, 10.0336559613546, 17.4319311777751, 17.2045957777235, 
    17.1266655392117, 17.1037693023682, 16.4507217407227, 16.2148696051704, 
    16.2770983378092, 16.2024088965522, 15.8356399536133, 15.6362585491604, 
    14.8103292253282, 14.3505212995741, 14.4962063895331, 15.0458743837145, 
    14.9758562511868, 13.791389465332, 12.9701467090183, 12.5238242679172, 
    12.920093536377, 13.2651773028904, 13.2902026706272, 13.2864519755046, 
    13.1227703094482, 13.1418646706475, 12.5879309972127, 11.6451784769694, 
    10.965217060513, 10.996886783176, 11.1746135287815, 11.2091870837741, 
    11.0596073998345, 11.1919777128432, 11.1708173751831, 10.732323328654, 
    10.383118947347, 10.2475580639309, 10.430459022522, 10.4234550264147, 
    10.5280135472616, 10.6547223197089, 10.4994524849786, 10.4587461683485, 
    10.2879297468397, 9.99062559339735, 9.73448912302653, 9.66484949323866, 
    9.67306031121148, 9.12308523390028, 8.60857031080458, 9.73774878184001, 
    9.93783940209283, 17.7426310645209, 17.2467839982775, 17.2558591630724, 
    17.0870255364312, 16.9140588972304, 16.6114891899957, 16.3309302859836, 
    16.2349757088555, 15.8012108272976, 15.3949406941732, 14.6569734149509, 
    14.4836086697049, 14.2996658749051, 14.3127856784397, 14.631756040785, 
    13.4556488460965, 13.0547329584757, 12.6089690526327, 12.5262390772502, 
    12.9076915582021, 13.1352797349294, 13.0529099305471, 12.9721416632334, 
    12.9142814477285, 12.631405433019, 11.639627456665, 11.005117336909, 
    10.9757498900096, 11.2637555599213, 11.290357430776, 11.1141438484192, 
    11.1396334966024, 11.0966595013936, 10.9864366849264, 10.6796259085337, 
    10.5795420805613, 10.4898873964945, 10.377782980601, 10.740374883016, 
    10.5609070460002, 10.4552805423737, 10.4709061781565, 10.2105224927266, 
    10.1404983997345, 9.89640402793884, 9.55968356132507, 9.61736567815145, 
    9.15096513430277, 9.5605727036794, 10.1349766254425, 9.917990843455, 
    17.3022912343343, 17.2915376027425, 17.3734007941352, 17.1806040869819, 
    17.290882534451, 17.0435678693983, 16.8217046525743, 16.2223552068075, 
    15.646653175354, 15.1500265333388, 14.4833731121487, 14.524974822998, 
    14.2387347751194, 14.0251733991835, 13.9268012576633, 13.2087199952867, 
    13.0942366917928, 12.6067266464233, 12.5793677171071, 12.5140307744344, 
    12.9733895460765, 12.9117290178935, 12.8015755812327, 12.7889177799225, 
    12.4964071114858, 11.8304862181346, 11.1511138280233, 11.2855168978373, 
    11.565601905187, 11.8879539966583, 11.2252229849497, 11.0755345026652, 
    10.9929705460866, 11.0652424494425, 11.0222911039988, 10.652756690979, 
    10.7282264232635, 10.6755494276683, 10.7168610095978, 10.51473681132, 
    10.512821038564, 10.501638174057, 10.0050985018412, 10.1516427199046, 
    9.78515823682149, 9.57314658164978, 9.57317193349203, 9.07371536890666, 
    10.0849494139353, 10.2379088401794, 9.95501446723938, 16.9740746815999, 
    16.8942970699734, 17.1102587381999, 17.2111373477512, 17.0644520653619, 
    16.9884149763319, 16.6795817481147, 16.1292503145006, 15.5100816090902, 
    14.8457256952922, 14.3423201243083, 14.6093082427979, 14.1656976275974, 
    14.2082139121162, 13.9503124025133, 13.2660470538669, 13.0683804617988, 
    12.7118395699395, 12.9518695407444, 12.7414744695028, 12.7286059061686, 
    12.7921856774224, 12.5535247590807, 12.5680008994208, 12.3134245342678, 
    12.077379544576, 11.7108671400282, 11.757499270969, 11.9454306496514, 
    12.0341949462891, 11.376263194614, 10.9505405426025, 11.1207387712267, 
    11.044123755561, 11.0109824074639, 10.6947761111789, 10.9235778384739, 
    10.8852110968696, 11.0443112055461, 10.9042001300388, 10.6588489744398, 
    10.6422628826565, 10.4492073059082, 10.1562774446276, 10.0087998708089, 
    9.61215782165527, 9.40678066677517, 9.37638007269965, 10.2657016118368, 
    10.141212993198, 9.82807985941569, 16.5641589694553, 16.7864089541965, 
    16.769844479031, 17.4961310492622, 17.0218609703912, 17.0287634531657, 
    16.4525731404622, 16.0954038831923, 15.723658879598, 14.8906761805216, 
    14.6168660057916, 14.6325047810872, 14.1287395689223, 14.1722588009304, 
    14.1593129899767, 13.505649778578, 13.077345000373, 12.7536098162333, 
    13.0262541770935, 12.9246857961019, 12.4908056259155, 12.3561503887177, 
    12.3698318799337, 12.5346681276957, 12.5720755259196, 12.3355650901794, 
    12.2937006950378, 11.7628772258759, 11.6831323305766, 11.6334730784098, 
    11.3377277056376, 10.9273862838745, 10.8067313035329, 10.7725114822388, 
    10.7135492960612, 10.6291739940643, 10.224999666214, 10.3875000476837, 
    10.359375, 10.4455355235509, 10.3803132375081, 10.5753334363302, 
    10.2445140566145, 9.7616774559021, 9.48951825228604, 9.23490405082703, 
    9.48468780517578, 10.0812103271484, 9.84556796334007, 9.52770177523295, 
    16.4022036658393, 16.3657383388943, 16.5491631825765, 16.7517846425374, 
    16.8795532650418, 16.6773317125108, 16.4428257412381, 15.9536216523912, 
    15.7590149773492, 15.0648759206136, 14.5261031256782, 14.5532442728678, 
    14.1375183529324, 14.1608899434408, 14.2248752382067, 13.5711562898424, 
    13.2958799997965, 12.9092145760854, 13.1161286036173, 13.1967673301697, 
    12.5328164100647, 12.253123998642, 12.1907619635264, 12.2594504356384, 
    12.7503277460734, 12.7308425108592, 12.3270847002665, 11.2912915547689, 
    11.4126833279928, 11.3542092641195, 11.0436531702677, 10.8888442516327, 
    10.8517874876658, 11.0424999757247, 10.7374998728434, 10.4382292429606, 
    10.1969999313354, 10.3062500953674, 10.197500038147, 10.1999998092651, 
    10.453125, 10.2929686307907, 9.16249990463257, 9.2854167620341, 
    9.59549989700317, 9.39770857493083, 9.78677225112915, 9.67499987284342, 
    9.70499992370605, 16.4472365909153, 16.324092441135, 16.5015936957465, 
    16.6630365583632, 16.5830006069607, 16.64574347602, 16.4932539198134, 
    16.2474066416423, 15.8686803181966, 15.1726971732246, 14.7735238605075, 
    14.5325618320041, 14.1010141372681, 14.2442448933919, 14.2043594784207, 
    13.7759033838908, 13.4057109620836, 13.2190894020928, 13.2015274895562, 
    13.2613598505656, 12.6793841256036, 12.3790841632419, 12.2591648101807, 
    12.3432820638021, 12.768692334493, 13.1034721798367, 11.9586341645983, 
    11.2172819773356, 11.5160697301229, 11.5247788959079, 11.334097120497, 
    10.2851851781209, 10.6541669368744, 10.3499999046326, 10.7302083969116, 
    11.0625, 10.3839288439069, 10.0362501144409, 11.0500001907349, 10.3125, 
    10.3862501144409, 9.75, 10.1999998092651, 9.54166666666667, 
    9.70666631062826, 9.76518938276503, 9.78986114925808, 10.2694665061103, 
    9.81944465637207, 9.82392480638292, 9.77708339691162, 16.3727325863308, 
    16.425689485338, 16.2975966135661, 16.4487592909071, 16.7254473368327, 
    16.3970553080241, 16.1210779613919, 16.212546772427, 16.112735218472, 
    15.3696445888943, 14.9236612319946, 14.3538378609551, 14.0494588216146, 
    14.263196627299, 14.4109831915961, 14.0616061952379, 13.5564122729831, 
    13.4027311007182, 13.4057706197103, 13.2890654404958, 12.7095372676849, 
    12.4876538912455, 12.2729818026225, 12.2731535434723, 12.4404068787893, 
    12.9239672025045, 11.819731314977, 11.1846250693003, 11.8114964167277, 
    11.560378854925, 11.2263888253106, 11.6118750572205, 11.8500003814697, 
    10.8900003433228, 10.4500001271566, 10.0406248569489, 10.1999998092651, 
    10.3078126907349, 10.2000002861023, 9.64204216003418, 9.58363395267063, 
    9.91185609499613, 9.77400024731954, 9.18947919209798, 9.72964421908061, 
    9.82457224527995, 9.37186543146769, 16.5706799825033, 16.604513168335, 
    16.4184457990858, 16.2329580518934, 16.1707442601522, 15.7429925070869, 
    16.0372923745049, 16.3541675143772, 16.4783642027113, 15.6719504462348, 
    15.2432831658257, 14.0683244069417, 13.909828291999, 14.0342269473606, 
    13.9330061806573, 13.8282095591227, 13.7222871780396, 13.6324714024862, 
    13.4452963670095, 13.3711846669515, 12.8486223220825, 12.4256115754445, 
    12.3681372801463, 12.5341523488363, 12.6078248818715, 12.5849274794261, 
    11.9713631470998, 11.4750076135, 11.6180965900421, 10.8225004196167, 
    11.6250001192093, 11.2763890160455, 8.625, 10.875, 9.8746874332428, 
    9.73693171414462, 9.60545444488525, 9.44629796346029, 8.29400690396627, 
    8.50310778617859, 8.63380159031261, 8.3155323266983, 16.6619249979655, 
    16.3247612847222, 16.3966727786594, 16.2913282182482, 16.2184419631958, 
    16.0607453452216, 15.978674782647, 16.1271110110813, 16.0291413201226, 
    15.7388139300876, 15.2097872628106, 14.1112162272135, 13.7374059889052, 
    13.6531474855211, 13.622554037306, 13.6083008448283, 13.725484000312, 
    13.6882996029324, 13.156261338128, 13.0467420154148, 12.7939172320896, 
    12.5313848919339, 12.3456312815348, 12.2808001836141, 12.0348637898763, 
    11.9450873268975, 11.7764410442776, 11.5850460264418, 8.24499979019165, 
    8.83703136444092, 8.65571673711141, 8.13243993123372, 16.5140448676215, 
    16.3230234781901, 16.3522012498644, 16.2969786326091, 16.2689734564887, 
    16.015230178833, 15.8514700995551, 15.931361940172, 15.805475446913, 
    15.2505209181044, 14.5980223549737, 14.1234780417548, 13.9184607399835, 
    13.7328272925483, 13.5142168468899, 13.2741550869412, 13.4903222190009, 
    13.6399835745494, 13.1961416403453, 12.9007976055145, 12.6945463816325, 
    12.8498746554057, 12.5563952128092, 12.2713366349538, 11.8334614146839, 
    16.5331645541721, 16.364187028673, 16.2841521369086, 16.1686462826199, 
    15.92754067315, 15.7410028245714, 15.4230078591241, 14.9539959165785, 
    14.5129081938002, 14.2449222140842, 14.1970852745904, 14.1741861767239, 
    14.1869130664402, 14.0097263124254, 13.5460466808743, 13.2326777776082, 
    13.2805486255222, 13.5336263179779, 13.2016479174296, 12.766566435496, 
    12.8220920562744, 12.5599935849508, 12.4218448003133, 12.07634973526, 
    16.6038597954644, 16.5156673855252, 16.3608623080783, 16.0791866514418, 
    15.8101507822673, 15.499446551005, 14.5192971759372, 14.2581359015571, 
    14.2023625903659, 14.0265281465318, 14.2044197718302, 14.1248016357422, 
    14.1972006691827, 14.1889118618435, 13.6775290171305, 13.2093381881714, 
    13.2615043852064, 13.3953879674276, 13.1230317221748, 13.1849196751912, 
    13.0083642535739, 12.4394025802612, 16.6424590216743, 16.4437077840169, 
    16.5516276889377, 16.087976137797, 15.7279567718506, 15.2799331876967, 
    14.1046301523844, 14.0488941404555, 14.1358157263862, 13.9478526645237, 
    14.1516244676378, 14.0654578738742, 14.2287861506144, 14.1602827707926, 
    13.6579386393229, 13.20754898919, 13.2424987157186, 13.459893544515, 
    13.5103556315104, 12.9808926582336, 12.6556489467621, 11.7840672492981, 
    16.4998965793186, 16.6501901414659, 16.5171930525038, 16.1847087012397, 
    15.5334700478448, 14.8879103130764, 13.9995861053467, 14.1505849626329, 
    14.1780576705933, 13.9164016511705, 14.0218182669746, 13.956203672621, 
    14.0840938356188, 13.7737268871731, 13.4711937374539, 13.1570962270101, 
    13.3236507839627, 13.3783466815948, 13.2886896928151, 12.7979076558893, 
    16.3950642479791, 16.7268986172146, 16.6561029222276, 16.4220485687256, 
    15.7097977532281, 14.9390098783705, 14.1184793048435, 14.2552797529433, 
    14.231750064426, 14.0930458704631, 14.0609507030911, 13.8806876076592, 
    14.0591660605537, 13.5774208704631, 13.4326086044312, 13.5325814353095, 
    13.4106767442491, 13.0715370178223, 12.7530767917633, 16.439006169637, 
    16.7028528849284, 16.7325738271077, 16.6549725002713, 16.1856139500936, 
    15.4497060775757, 14.7032270431519, 14.5607945124308, 14.4572270711263, 
    14.1499063703749, 13.9991596009996, 13.8610765669081, 13.8843505647447, 
    13.9023983213637, 13.735852877299, 13.6126681433784, 13.2512315511703, 
    16.0899913575914, 16.0525305006239, 16.2904851701525, 16.6302602556017, 
    16.6716819339328, 16.3437392976549, 15.6239958869086, 15.2742275661892, 
    14.5786729388767, 14.3867282867432, 13.9765875074599, 13.6398431989882, 
    13.478899108039, 13.5777011447483, 13.5028555128309, 13.3067380905151, 
    16.2068144480387, 15.9232803980509, 16.0462001164754, 16.53820376926, 
    16.6030871073405, 16.5839795006646, 16.1331043243408, 15.5778775744968, 
    14.7687424553765, 14.6740702523126, 14.1620410283407, 13.3845592074924, 
    13.2746832105849, 13.3051026662191, 13.1336999469333, 16.3684741126166, 
    16.0874963336521, 15.7142188813951, 16.3143032921685, 16.5479772355821, 
    16.5178209940592, 16.2935203976101, 15.8225991990831, 15.2659853829278, 
    14.4704221089681, 13.8783077663845, 13.5206939909193, 13.0379188855489, 
    12.8501987457275, 16.394600338406, 16.2023684183757, 15.7180952495999, 
    15.9947347640991, 16.3293688032362, 16.1478969785902, 15.8493882285224, 
    15.4642003377279, 15.0793790817261, 14.161416053772, 13.4991675615311, 
    13.563195016649, 16.4593230353461, 16.1983723110623, 15.750404993693, 
    15.5719236797757, 15.5858874850803, 15.3222267362807, 14.9526377783881, 
    14.7208382288615, 14.6554622650146, 13.9821109771729, 13.6062479019165, 
    13.6595776875814, 16.4533333248562, 16.2513015535143, 15.9043964809842, 
    15.5947280459934, 15.2626521852281, 15.0579289330377, 14.8063691457113, 
    14.3365809122721, 14.2872684266832, 13.7550080617269, 13.8551460901896, 
    13.5207580990261, 16.3158927493625, 16.2043800354004, 15.8539445665148, 
    15.6470822228326, 15.5958701239692, 15.606875843472, 14.6812529034085, 
    14.3407680723402, 14.0926985210843, 13.9365146425035, 14.0482921600342, 
    16.2094508277045, 15.8767967224121, 15.7680886586507, 15.727460331387, 
    15.7971051534017, 15.7167098787096, 14.4850766923692, 14.4568254682753, 
    14.2645647260878, 14.184963438246, 14.2129074732463, 15.9832297431098, 
    15.6064812342326, 15.7826724582248, 15.8883006837633, 15.778157764011, 
    15.5188763936361, 14.8337375852797, 14.752785258823, 14.589465353224, 
    14.5044542948405, 14.3177603085836, 15.764713605245, 15.584216647678, 
    15.4937999513414, 15.737473487854, 15.1769664552477, 15.1558961868286, 
    15.0613864262899, 14.9855097664727, 14.9620975255966, 14.6877051989237, 
    15.4131152894762, 15.5294861263699, 15.2924204932319, 15.3540030585395, 
    15.1913794411553, 15.2409071392483, 15.1095952987671, 15.0799673928155, 
    15.1124964820014, 15.7624419530233, 15.7824169794718, 15.4803779390123, 
    15.1959829330444, 15.2595366372002, 15.259891404046, 15.1860720316569, 
    15.1839969423082, 14.9985092878342, 16.298166486952, 16.1154217190213, 
    16.2535994847616, 15.7027917438083, 15.4867106543647, 15.0263305240207, 
    15.0185871124268, 14.8061496734619, 16.5446578131782, 16.3696399264865, 
    16.5107989841037, 15.477232615153, 14.9267551634047, 16.1303270128038, 
    15.6558390723334, 15.7767386966281, 14.8098753293355, 11.2923981802804, 
    11.2992696762085, 11.2982950210571, 11.2970762252808, 11.2958545684814, 
    11.294629573822, 11.2391742070516, 10.14399822553, 8.83433310190837, 
    7.81750647226969, 9.48060637253981, 8.3945129101093, 7.37896112295297, 
    9.05040022043081, 7.81111368766198, 6.78067544790415, 9.78600271542867, 
    8.49324591954549, 7.2356166044871, 6.28707544008891, 11.3992643356323, 
    11.3982839584351, 11.397057056427, 11.395827293396, 11.3945941925049, 
    11.0060035387675, 11.4494684764317, 14.2498426437378, 14.1591596603394, 
    13.9784469604492, 12.437292098999, 12.0860271453857, 11.6548728942871, 
    11.4536552429199, 33.2130012512207, 33.2099990844727, 33.2060012817383, 
    33.1650009155273, 33.2050018310547, 33.2439994812012, 33.3199996948242, 
    14.5496816635132, 14.5485038757324, 14.547080039978, 14.5456113815308, 
    13.9343614578247, 12.113597869873, 11.5768885612488, 10.8239393234253, 
    10.4896655082703, 33.2140007019043, 33.2169990539551, 33.2190017700195, 
    33.2140007019043, 33.1669998168945, 33.185001373291, 33.2880001068115, 
    33.5415000915527, 33.751501083374, 17.4407428105672, 17.5064427057902, 
    17.764352162679, 17.2335424423218, 16.8680308659871, 16.827561378479, 
    16.5930344263713, 16.4485470453898, 16.3762029012044, 16.3291994730632, 
    16.2919165293376, 16.2883930206299, 15.9193553924561, 15.5074424743652, 
    15.2779763539632, 14.8105263710022, 14.2899905840556, 14.2428450584412, 
    13.9191869099935, 13.5803155899048, 13.2652708689372, 13.2064512570699, 
    13.1351172129313, 13.1786985397339, 13.2495759328206, 13.3462985356649, 
    13.3576793670654, 12.9369489351908, 12.384074529012, 11.8705547650655, 
    11.7326839764913, 11.8096005121867, 11.6234501202901, 11.2959068616231, 
    10.8587563832601, 10.7948732376099, 10.5698078473409, 10.6259299914042, 
    10.7241797447205, 10.8368198076884, 10.4992993672689, 10.4059850374858, 
    10.6148476600647, 10.4257300694784, 10.3511358896891, 10.4992863337199, 
    10.1503248214722, 9.89671421051025, 9.70059219996134, 9.35493564605713, 
    9.22393369674683, 17.5388819376628, 17.3847348954942, 17.5870585971408, 
    17.4175179799398, 16.9635384877523, 16.7779210408529, 16.5465571085612, 
    16.4346084594727, 16.3184941609701, 16.3516354031033, 16.2787736256917, 
    16.2906379699707, 16.0462183422512, 15.6532618204753, 15.4636304643419, 
    14.9801843431261, 14.3810562557644, 14.4178789456685, 14.0910464127858, 
    13.8216909567515, 13.5610047181447, 13.4476498762767, 13.3211879730225, 
    13.361141761144, 13.4090408484141, 13.3806128501892, 13.3229986826579, 
    12.8492257595062, 12.1944622993469, 11.9729450543722, 11.7037199338277, 
    11.6540182431539, 11.3939089775085, 11.3173433144887, 10.9852752685547, 
    10.7588144938151, 10.6383197307587, 10.8193749586741, 11.0014649232229, 
    10.9779201348623, 10.7009816964467, 10.5188834667206, 10.53559923172, 
    10.4537117481232, 10.4813772837321, 10.3381107648214, 9.92720603942871, 
    9.91082525253296, 9.4888121287028, 9.82123525937398, 9.43304228782654, 
    17.2280868954129, 17.0269304911296, 17.2656375037299, 17.2895035213894, 
    16.9593048095703, 16.5276118384467, 16.3826402028402, 16.3707754347059, 
    16.2427618238661, 16.2650176154243, 16.2123875088162, 16.1479350195991, 
    15.9141688876682, 15.7642867830065, 15.5199688805474, 15.134042845832, 
    14.7055932150947, 14.6951745351156, 14.4936854044596, 14.2109311421712, 
    13.9432559013367, 13.8570148150126, 13.7737342516581, 13.6777450243632, 
    13.5949985186259, 13.31573955218, 13.1705929438273, 12.7601448694865, 
    12.0645410219828, 11.772305727005, 11.8752253055573, 11.6757500171661, 
    11.6573831240336, 11.4326567649841, 11.1641902923584, 10.9662425518036, 
    10.8254458109538, 10.9798767566681, 11.1079564889272, 10.98406513532, 
    10.6595888137817, 10.6160031159719, 10.5024708112081, 10.3648361365, 
    10.2591973145803, 10.0444253285726, 9.70507113138835, 9.57716075579325, 
    9.78680316607157, 9.72938895225525, 9.77437766393026, 17.2973376380073, 
    17.1524969736735, 17.2719898223877, 17.0888646443685, 16.7700231340196, 
    16.3436459435357, 16.231930202908, 16.1967368655735, 16.0700204637316, 
    16.2520463731554, 16.1152317259047, 16.0562629699707, 16.0002245373196, 
    15.8805467817518, 15.5060858196682, 15.2457278569539, 14.9094950358073, 
    14.8931783040365, 14.1325806511773, 13.6351594924927, 13.5974298053318, 
    13.9370345009698, 13.9151313569811, 13.7510693868001, 13.5764740837945, 
    13.2057483461168, 12.9598259396023, 12.4068162706163, 11.7518193986681, 
    11.4442266888089, 11.4316877788968, 11.4834878709581, 11.523166762458, 
    11.6120381885105, 11.2007990943061, 11.1372691260444, 10.9677833980984, 
    11.0022110409207, 11.1484022140503, 10.893433464898, 10.7816914452447, 
    10.6569577323066, 10.3810400433011, 10.0717275407579, 9.89221668243408, 
    9.69908693101671, 9.28733942243788, 9.38884109920926, 9.55215930938721, 
    9.75488313039144, 9.34801959991455, 17.7018775939941, 17.4660538567437, 
    17.0549979739719, 16.7113265991211, 16.5339397854275, 16.4405858781603, 
    16.1599079767863, 16.1559916602241, 16.0877589119805, 16.0775277879503, 
    16.0705021752252, 16.0257070329454, 15.9832550684611, 15.8134645885891, 
    15.6235647201538, 15.3505655924479, 15.1098574532403, 14.2944447199504, 
    13.2946399052938, 13.0783290068309, 13.149749994278, 13.388511578242, 
    13.5594705740611, 13.6090795993805, 13.4336241881053, 12.8791151841482, 
    12.6679384708405, 12.1780090332031, 11.5887352625529, 11.3268880049388, 
    11.0781365235647, 11.0822907288869, 11.1047673225403, 11.375014146169, 
    11.216010093689, 11.0769859949748, 10.8608965873718, 10.8306731383006, 
    10.9714101155599, 10.8616866270701, 10.5439930756887, 10.5260449250539, 
    10.1821023623149, 9.71200331052144, 9.47475401560465, 9.3314962387085, 
    9.24781084060669, 9.48219537734985, 9.5135924021403, 9.69603045781454, 
    9.38164075215658, 17.2075252532959, 16.9164377848307, 16.7531000773112, 
    16.5877537197537, 16.7883904774984, 16.5199752383762, 16.2837166256375, 
    16.1371264987522, 15.8683258692423, 15.8821942011515, 15.853571150038, 
    15.8107686572605, 15.7012091742622, 15.6009178161621, 15.5611710018582, 
    15.1619083616469, 14.4493289523655, 13.5348171393077, 12.9620436827342, 
    12.9337914784749, 13.1298352877299, 13.3412856260935, 13.4175929228465, 
    13.4418710072835, 13.1746949354808, 12.5877104600271, 12.3172214031219, 
    11.8356481393178, 11.4718464215597, 11.2276880741119, 11.049028635025, 
    11.045089006424, 10.777866601944, 11.0523693561554, 10.8674148718516, 
    10.7759142716726, 10.638058423996, 10.6974539756775, 10.7858820756276, 
    10.5803984006246, 10.3985203107198, 10.176100174586, 9.82352526982625, 
    9.50128157933553, 9.58844033877055, 9.41781783103943, 9.30671898523966, 
    9.43633111317953, 9.37206546465556, 9.26343854268392, 9.26848371823629, 
    17.1495793660482, 17.160275777181, 16.6843255360921, 16.7523517608643, 
    16.8459964328342, 16.7128092447917, 16.2409269544813, 16.1007401148478, 
    15.760520723131, 15.6748655107286, 15.7049721611871, 15.6856836742825, 
    15.3641019397312, 15.3640046649509, 15.3919418123033, 14.9956979751587, 
    13.8114958869086, 13.0324186748928, 12.9487299389309, 13.1909761428833, 
    13.307394557529, 13.2388354407416, 13.3503861957126, 13.4363278283013, 
    12.8917186525133, 12.3260537253486, 11.8344400193956, 11.3805688222249, 
    11.1254505581326, 11.2302769554986, 11.1426777309842, 11.0945937898424, 
    10.8149979909261, 10.605357170105, 10.4693428675334, 10.3603999879625, 
    10.6697557237413, 10.6357243855794, 10.6634780036079, 10.5452874501546, 
    10.412646399604, 10.0837711758084, 9.7818816502889, 9.75718678368462, 
    9.78448602888319, 9.74895371331109, 9.32527054680718, 9.30478074815538, 
    9.29707770877414, 8.99779510498047, 9.13979456159804, 17.4451722039117, 
    17.2140373653836, 16.7872655656603, 16.7631732092963, 16.7930043538411, 
    16.6958406236437, 16.1672666337755, 16.1281063291762, 15.6475074556139, 
    15.6268667644925, 15.5411672592163, 15.3998907936944, 15.2880375120375, 
    15.2221475177341, 15.1643510394626, 14.420831574334, 13.2205651601156, 
    12.8584336439768, 13.0872968037923, 13.3223929405212, 13.3420946598053, 
    13.2794845104218, 13.3202245235443, 13.393151919047, 12.6596268018087, 
    12.1054422855377, 11.4106761614482, 11.1398917039235, 11.2859503428141, 
    11.1817394892375, 11.0647996266683, 11.0475951830546, 10.9447310765584, 
    10.5362267494202, 10.3696255683899, 10.404568751653, 10.4971151351929, 
    10.5301187038422, 10.5467182000478, 10.7386531829834, 10.6735095977783, 
    10.2884788513184, 9.90359576543172, 9.87823494275411, 9.85761181513468, 
    9.80824685096741, 9.50787790616353, 9.24784366289775, 9.21554613113403, 
    9.22816379865011, 9.68614284197489, 17.2389657762316, 17.332245932685, 
    17.255656560262, 16.7640213436551, 16.6935878329807, 16.249267578125, 
    16.1523412068685, 16.1110719045003, 15.5311112933689, 15.6546027925279, 
    15.165211253696, 14.6333677503798, 15.0711234410604, 15.144739151001, 
    15.1143581602308, 14.0374298095703, 13.0008378558689, 12.7053413391113, 
    13.142558892568, 13.3481151262919, 13.3473348617554, 13.2762741247813, 
    13.3252313931783, 13.280979235967, 12.5711283683777, 11.8401406606038, 
    11.1244633992513, 10.9418803056081, 11.1679409344991, 11.2313680648804, 
    10.8518197536469, 10.9485379060109, 11.0215732256571, 10.6116544405619, 
    10.3708675702413, 10.2186657587687, 10.2908293406169, 10.4383146762848, 
    10.5260616143545, 10.8519035975138, 10.7561483383179, 10.4498000144958, 
    10.1359905401866, 10.1063567002614, 10.1439924240112, 9.93781924247742, 
    9.61387777328491, 9.01830410957336, 9.17745772997538, 9.38219960530599, 
    9.75135882695516, 17.3454564412435, 17.3196603986952, 17.2995476192898, 
    16.920093536377, 16.2710818184747, 16.1630704667833, 16.2776605818007, 
    16.2184268103706, 15.7960197660658, 15.4518435796102, 14.8270867665609, 
    14.3459048800998, 14.5228421952989, 15.0626765357123, 15.0173397064209, 
    13.8168202506171, 12.9780972798665, 12.5278317133586, 12.8998722500271, 
    13.2642650604248, 13.2913848029243, 13.2883005142212, 13.1246996985541, 
    13.2212892108493, 12.6469249725342, 11.6443809933133, 10.9356098175049, 
    10.8593222300212, 10.9832741419474, 11.1199855804443, 10.8565094206068, 
    11.0441283120049, 11.1678572760688, 10.6329860687256, 10.4844217300415, 
    10.2186432944404, 10.3461641735501, 10.5795370737712, 10.6958471934001, 
    10.8045403162638, 10.5442174275716, 10.2853151957194, 10.202297422621, 
    10.216908454895, 9.97555213504367, 9.84572675493028, 9.47333611382378, 
    9.00349892510308, 8.55416059494019, 9.40628221299913, 9.61893325381809, 
    17.3993856641981, 17.3096018897163, 17.1915726131863, 17.1112217373318, 
    16.7407631344265, 16.5061451594035, 16.20858446757, 16.2470009062025, 
    15.8547709782918, 15.295890490214, 14.6251624425252, 14.4858654869927, 
    14.3394242392646, 14.3275000254313, 14.6703714794583, 13.4823314878676, 
    13.0550354851617, 12.6083656946818, 12.5174624125163, 12.9023237228394, 
    13.1393434206645, 13.0521223545074, 13.0329984823863, 12.9624485174815, 
    12.6550550460815, 11.6068156560262, 10.9220371246338, 10.9105775356293, 
    11.112429857254, 11.2496868769328, 11.0048973560333, 11.1257005532583, 
    11.0968091487885, 11.1034553845723, 10.8463124434153, 10.6015605926514, 
    10.3745791912079, 10.3327125708262, 10.724063316981, 10.5063453515371, 
    10.3605902194977, 10.216811577479, 10.2523464361827, 10.1469423770905, 
    9.83370288213094, 9.70165681838989, 9.54609886805216, 8.98902837435404, 
    9.36967412630717, 9.76374459266663, 9.75933615366618, 17.3326816558838, 
    17.1926663716634, 17.2495405409071, 17.1791195339627, 17.1378752390544, 
    16.7347558339437, 16.8453004625108, 16.2091883553399, 15.429412206014, 
    15.2000592549642, 14.4381632275052, 14.5834415223863, 14.2839691374037, 
    14.0598793029785, 13.9551079008314, 13.2249391343859, 13.1161798901028, 
    12.6196520328522, 12.6025187969208, 12.4885989824931, 13.0020501613617, 
    12.9303077061971, 12.8759775161743, 12.8731809457143, 12.5235437552134, 
    11.8249980608622, 11.0693385601044, 11.0548654397329, 11.2647552490234, 
    11.6467224756877, 11.24707086881, 11.1310584545135, 10.982291618983, 
    11.1407237052917, 11.1377499898275, 10.6342956225077, 10.645429054896, 
    10.5664873917898, 10.5935509204865, 10.3854250907898, 10.429660876592, 
    10.1516771316528, 10.0595843791962, 9.98465387026469, 9.75417447090149, 
    9.62610459327698, 9.50410087903341, 8.85821111996969, 9.95434641838074, 
    10.0515115261078, 9.7966882387797, 16.9656567043728, 16.831217235989, 
    16.9842688242594, 17.1450551350911, 17.0702472262912, 16.7899434831407, 
    16.6386144426134, 16.1530777613322, 15.299816555447, 14.9069203270806, 
    14.342488500807, 14.6631540722317, 14.2362846798367, 14.2684552934435, 
    14.0251836776733, 13.2357094022963, 13.054008907742, 12.7317117055257, 
    12.9805680380927, 12.7424490186903, 12.7436338000827, 12.8523179160224, 
    12.6534523434109, 12.6879812876383, 12.3202108807034, 11.9466883341471, 
    11.6239674886068, 11.3508372836643, 11.4637777540419, 11.66117699941, 
    11.3213027318319, 10.9387145572239, 11.0763154559665, 11.1426271862454, 
    10.9717258877224, 10.6548399395413, 10.7726944817437, 10.7227221594916, 
    10.7728110419379, 10.6327815585666, 10.5591249465942, 10.6058443917169, 
    10.0873055987888, 10.0147630903456, 9.80386585659451, 9.53582106696235, 
    9.47573068406847, 9.36817889743381, 9.93648264143202, 9.94683922661675, 
    9.72611151801215, 16.5090866088867, 16.6492144266764, 16.5952010684543, 
    17.0870407952203, 17.0446253882514, 16.9105008443197, 16.5867349836561, 
    16.0734278361003, 15.5878033108181, 14.935258547465, 14.5920299953885, 
    14.7352751625909, 14.19295946757, 14.2609718110826, 14.2289105521308, 
    13.4687583711412, 13.072898334927, 12.7608649730682, 13.0300293763479, 
    12.9030222098033, 12.5059202512105, 12.3714435100555, 12.3716680208842, 
    12.5713256994883, 12.5846848487854, 12.2934060891469, 12.2442331314087, 
    11.5323920683427, 11.5366507371267, 11.2615408463912, 10.8983155091604, 
    10.9227740547874, 10.792551279068, 10.7312454743819, 10.650000163487, 
    10.5281248092651, 10.4249992370605, 10.6836331685384, 10.1145162582397, 
    9.95956659317017, 9.50840441385905, 9.49896543676203, 9.39450287818909, 
    9.59418145815531, 9.91887863477071, 9.61937618255615, 9.44110608100891, 
    16.4035523732503, 16.3142681121826, 16.5729031032986, 16.7710522545709, 
    16.8290365007189, 16.6737128363715, 16.3198290930854, 16.1466997994317, 
    15.6035884221395, 14.8371493021647, 14.4870315127903, 14.5612229241265, 
    14.179835319519, 14.2306594848633, 14.2765067418416, 13.602996190389, 
    13.3350132836236, 12.8932615915934, 13.0981513659159, 13.1980506579081, 
    12.5831123193105, 12.2895526091258, 12.2410128911336, 12.3164131641388, 
    12.7605063120524, 12.7312200069427, 12.7159857749939, 11.3623367656361, 
    11.4062498410543, 11.1837647755941, 10.8795456452803, 10.9799999237061, 
    11.0142856325422, 10.5843750238419, 10.2750002543132, 10.5166666242811, 
    10.3874998092651, 10.03125, 9.65416669845581, 8.96875023841858, 
    9.49319038391113, 9.40146327018738, 9.73913892110189, 9.74921894073486, 
    9.62161461512248, 9.37903650601705, 16.3795827229818, 16.2851816813151, 
    16.5504048665365, 16.6814301808675, 16.5837773217095, 16.3863308164809, 
    16.2746351030138, 16.1323926713732, 15.8835319942898, 15.1011437310113, 
    14.7245102988349, 14.5585074954563, 14.126759952969, 14.3155279159546, 
    14.238107363383, 13.7243324915568, 13.3479553858439, 13.1800669564141, 
    13.1059674157037, 13.2116081449721, 12.6628757052951, 12.4210115008884, 
    12.4139116075304, 12.400127198961, 12.8697915607029, 13.4221063190036, 
    12.3515621423721, 11.2529466152191, 11.6287038591173, 11.5458333151681, 
    10.7699998855591, 10.5, 10.5, 9.63333320617676, 9.37395842870077, 
    9.76518938276503, 9.78986114925808, 10.2694665061103, 9.90138891008165, 
    9.76132678985596, 9.47968745231628, 16.3703763749864, 16.4563965267605, 
    16.3210928175184, 16.4553356170654, 16.6786566840278, 16.3975166744656, 
    16.1324668460422, 16.14061027103, 16.1756214565701, 15.3383597267999, 
    14.9030765957303, 14.3666244082981, 14.0920908186171, 14.329021135966, 
    14.43235206604, 14.0709100299411, 13.505552927653, 13.378001610438, 
    13.3943320115407, 13.2420449256897, 12.7390654881795, 12.5082244873047, 
    12.3541289965312, 12.3027341365814, 12.6718462308248, 13.0088854630788, 
    11.9913904666901, 11.1067533493042, 11.7124998786233, 11.3156249523163, 
    11.7225001335144, 11.8500003814697, 10.1999998092651, 9.62381303310394, 
    9.61759195327759, 9.91185609499613, 9.77400024731954, 9.18947919209798, 
    9.72964421908061, 9.80972862243652, 9.35545913378398, 16.5448188781738, 
    16.5985190073649, 16.4025565253364, 16.2700097825792, 16.2002195782132, 
    15.7051146825155, 16.0710322062174, 16.1290545993381, 16.5095568762885, 
    15.7875632180108, 15.2732830047607, 14.0392749574449, 13.9646011988322, 
    14.0643662346734, 13.9311156802707, 13.703929371304, 13.6686912112766, 
    13.6177020867666, 13.392098903656, 13.3191967010498, 12.8195343812307, 
    12.4510075251261, 12.4402766227722, 12.5910322666168, 12.664484500885, 
    12.7201476891836, 12.1219833691915, 11.2848091920217, 11.44553565979, 
    11.3250001907349, 11.9250001907349, 11.8500003814697, 9.8746874332428, 
    9.73693171414462, 9.60545444488525, 9.44629796346029, 8.29400690396627, 
    8.50310778617859, 8.63380159031261, 8.3155323266983, 16.6686242421468, 
    16.2902003394233, 16.3084083133274, 16.3120678795709, 16.3031611972385, 
    16.0414367251926, 16.0379333496094, 16.1350136862861, 16.0906114578247, 
    15.7648499806722, 15.3466540442573, 14.1293622122871, 13.7447201410929, 
    13.7007037268745, 13.6676157845391, 13.6110110812717, 13.7058689329359, 
    13.7111066182454, 13.178112771776, 13.1209448708428, 13.0040133794149, 
    12.666385544671, 12.4482323328654, 12.3404637442695, 12.1623722712199, 
    11.9744389851888, 11.8500232696533, 11.2524299621582, 8.24499979019165, 
    8.83703136444092, 8.65571673711141, 8.13243993123372, 16.5403406355116, 
    16.2991564008925, 16.3235251108805, 16.2656892140706, 16.2426399654812, 
    15.9517093234592, 15.8531581030952, 15.9068330128988, 15.7737753126356, 
    15.285098499722, 14.560937139723, 14.0976078245375, 13.8938873079088, 
    13.746277279324, 13.5482607947456, 13.3171566857232, 13.4715812471178, 
    13.6405780315399, 13.2797427972158, 13.0696603457133, 12.8959363301595, 
    12.9297362963359, 12.6171340942383, 12.3343273003896, 11.930721282959, 
    16.5466471778022, 16.3573864830865, 16.2689880794949, 16.1528973049588, 
    15.8969090779622, 15.7134613460965, 15.3852313359578, 14.9673113293118, 
    14.5700451533, 14.1746077007718, 14.0748168097602, 14.1612963146634, 
    14.1691550148858, 14.0053785112169, 13.5664491653442, 13.273754119873, 
    13.341518719991, 13.5921570460002, 13.3301290671031, 12.8692685763041, 
    12.974893172582, 12.5955250263214, 12.3460294405619, 11.9625511964162, 
    16.5912823147244, 16.4888617197673, 16.3214685651991, 16.0676229265001, 
    15.811291164822, 15.4803152084351, 14.4917457368639, 14.2731217278375, 
    14.2016354666816, 13.9625874625312, 14.123663160536, 14.1206193500095, 
    14.1267320844862, 13.9399176703559, 13.6106033325195, 13.2470088534885, 
    13.2922394010756, 13.4491234885322, 13.2477052476671, 13.2772703170776, 
    12.8879157172309, 12.101151254442, 16.5681726667616, 16.4052965376112, 
    16.3595566219754, 16.0470709270901, 15.7064392301771, 15.2620561387804, 
    14.0825543933445, 14.0308244493273, 14.1257830725776, 13.9278650283813, 
    14.1307524575127, 14.0774013731215, 14.1947414610121, 13.967144648234, 
    13.5602890650431, 13.082618077596, 13.1582802666558, 13.5898067951202, 
    13.608067035675, 13.0262001355489, 12.7287352879842, 11.4739905463325, 
    16.4649800194634, 16.5980508592394, 16.3801023695204, 16.0660315619575, 
    15.5540285110474, 14.9219880633884, 13.9893618689643, 14.1293178134494, 
    14.1629536946615, 13.9036535686917, 13.9691696166992, 13.9478034973145, 
    13.9750117195977, 13.7919626235962, 13.5572706858317, 13.3497524261475, 
    13.4293732113308, 13.4464832146962, 13.4504771232605, 12.8857918652621, 
    16.3486164940728, 16.6404033237033, 16.4792291853163, 16.2229801813761, 
    15.5113397174411, 14.9442427953084, 14.0887400309245, 14.2185688018799, 
    14.1997281180488, 14.0008041593764, 13.9454485575358, 13.7786398993598, 
    13.8965869479709, 13.5396828121609, 13.4341702991062, 13.6906346215142, 
    13.4519143634372, 13.1300687789917, 12.8366248607635, 16.3872392442491, 
    16.5062005784776, 16.5732460021973, 16.4525623321533, 16.0209333631727, 
    15.3451657825046, 14.5566850238376, 14.3687194188436, 14.2715724309285, 
    14.0126350190904, 13.8952207565308, 13.7502189212375, 13.7664789623684, 
    13.8529929055108, 13.7643551296658, 13.7043863932292, 13.2737722396851, 
    15.9179693857829, 15.9174177381727, 16.184186829461, 16.5807469685872, 
    16.5858296288384, 16.1775312423706, 15.3630091349284, 15.0879450903998, 
    14.529887093438, 14.2942399978638, 14.0433411068386, 13.6355029212104, 
    13.3580771552192, 13.4330078760783, 13.3101497226291, 13.2927070617676, 
    16.1044073104858, 15.8153400421143, 15.8336805767483, 16.4906862046983, 
    16.5301130082872, 16.475759294298, 15.9965153800117, 15.3403729332818, 
    14.7022546132406, 14.6283237669203, 14.183831108941, 13.3352387746175, 
    13.0657759772407, 13.0975022845798, 12.9501637352837, 16.1508238050673, 
    15.9797801971436, 15.533943494161, 16.2363501654731, 16.4382199181451, 
    16.3980880313449, 16.1896562576294, 15.6999911202325, 15.2381004757351, 
    14.4418787426419, 13.8279796176487, 13.4138003455268, 12.935110727946, 
    12.7844624519348, 16.2123974694146, 16.0621469285753, 15.6485826704237, 
    15.908673286438, 16.136890411377, 15.9293148252699, 15.6358903249105, 
    15.5702592002021, 15.0375299453735, 14.1145265367296, 13.4959172010422, 
    13.5376958847046, 16.2105462816026, 16.020029703776, 15.7237539291382, 
    15.3971811930339, 15.4040927886963, 14.8364209069146, 14.515329890781, 
    14.5084833568997, 14.4978573057387, 13.7617637846205, 13.4182469844818, 
    13.5606429841783, 16.2186965942383, 16.1408280266656, 15.8971775902642, 
    15.4921375910441, 15.0573002497355, 14.8071065478855, 14.4910953309801, 
    14.012776904636, 13.9995483822293, 13.4567006429036, 13.6281622250875, 
    13.5268115997314, 16.2446433173286, 16.0896283255683, 15.8415665096707, 
    15.4797661039564, 15.3096743689643, 15.2935651143392, 14.5714815987481, 
    14.0180371602376, 13.8443880081177, 13.6807550854153, 13.9667943318685, 
    16.1735319561428, 15.7790868547228, 15.7452500661214, 15.5913184483846, 
    15.4693118201362, 15.4816409216987, 14.4053270551893, 14.3087112638685, 
    14.1790743933784, 14.1159703996446, 14.2450405756632, 15.9771455128988, 
    15.5414890713162, 15.6925684611003, 15.7076189253065, 15.5450375874837, 
    15.428720580207, 14.8341129091051, 14.6506801181369, 14.5217547946506, 
    14.5445288552178, 14.3421430587769, 15.5865556928847, 15.6450942357381, 
    15.5338409211901, 15.6636292139689, 15.2317417992486, 15.1451901329888, 
    15.0424250496758, 15.1217485004001, 14.9169813394547, 14.5601162910461, 
    15.4519237942166, 15.7415877448188, 15.6251748402913, 15.3610517713759, 
    15.3192720413208, 15.3796740637885, 15.2405783335368, 15.1997252570258, 
    15.0989309946696, 15.8144754833645, 16.1962887446086, 16.1938959757487, 
    15.4698594411214, 15.5309147304959, 15.4333029852973, 15.2230326334635, 
    15.1915273666382, 14.949490070343, 16.700472301907, 16.595744450887, 
    16.7995482550727, 16.1722103754679, 15.5820879406399, 14.944575521681, 
    14.7628289631435, 14.679020690918, 16.8256736331516, 16.7021617889404, 
    16.6389781104194, 15.6932711071438, 14.9854067696465, 16.5309825473362, 
    16.0329845216539, 15.9251018100315, 14.8757115999858, 14.9297780990601, 
    14.8884220123291, 14.8870038986206, 14.8955249786377, 14.8840341567993, 
    13.2351795832316, 11.0896244049072, 10.2727085749308, 9.39949893951416, 
    33.185001373291, 33.185001373291, 33.1860008239746, 33.1839981079102, 
    33.185001373291, 33.1126670837402, 33.2529983520508, 33.6459999084473, 
    34.0149993896484, 14.7791595458984, 14.617115020752, 14.6057024002075, 
    14.6041698455811, 14.4727430343628, 12.4565010070801, 10.8639149665833, 
    10.0750846862793, 9.47451257705688, 9.07508945465088, 8.74132251739502, 
    8.067458152771, 7.35319900512695, 6.89866304397583, 6.34328508377075, 
    33.1900005340576, 33.1889991760254, 33.1940002441406, 33.189998626709, 
    33.1749992370605, 33.1359996795654, 33.4914989471436, 33.8134994506836, 
    34.1079998016357, 34.1990013122559, 34.2270011901855, 34.2589988708496, 
    34.2700004577637, 34.3019981384277, 34.3190002441406, 0.212599942698479, 
    0.192569131261999, 0.186839991967246, 0.1624202385672, 0.17125966474767, 
    0.152691910106491, 0.146031144711369, 0.176656513774725, 0.1348015039948, 
    0.196810728421345, 0.213358404662935, 0.156765985592722, 
    0.180619047954168, 0.226560081928098, 0.207255486524237, 
    0.196013042496556, 0.153787041517729, 0.212368519736534, 
    0.188540460109794, 0.219034055699219, 0.135877917161369, 
    0.203849114453924, 0.192228451632657, 0.159163592833512, 
    0.220391871304086, 0.132698624667742, 0.193613397121513, 
    0.185316122295004, 0.13873319565751, 0.187544003597041, 
    0.206840486321561, 0.140153379016548, 0.178375476378434, 
    0.189879470447559, 0.131266283973526, 0.192476386362354, 
    0.190877864015158, 0.158797417202507, 0.159229716653604, 
    0.186730455619295, 0.161533416395419, 0.133754848955624, 
    0.203181411961557, 0.181360249032948, 0.176701251530931, 
    0.13724620340712, 0.172981160029312, 0.181072427578701, 
    0.147862717384563, 0.195725181429943, 0.170200980298433, 
    0.0912231296053067, 0.172483917087538, 0.123530239580624, 
    0.171583434476126, 0.213740190417576, 0.164966228226658, 
    0.159621184785021, 0.158900262589309, 0.126065558610503, 
    0.150649242556255, 0.130654465431438, 0.182281570045718, 
    0.220499482447659, 0.0843297692879802, 0.163648368880922, 
    0.124864876720244, 0.163739237794475, 0.171729689857581, 
    0.132089284924213, 0.15085291645908, 0.178807922120056, 
    0.182203255578128, 0.116154925343958, 0.144601868916778, 
    0.125835649954296, 0.176666248764831, 0.194565451964035, 
    0.125656084372902, 0.0951966210946208, 0.154974357650454, 
    0.168772842309619, 0.139275560794601, 0.154757899364474, 
    0.129484572267521, 0.152559342177834, 0.176254276864559, 
    0.186633040052655, 0.125069578592439, 0.121059100148645, 
    0.137982911397246, 0.174034401284763, 0.141161124197121, 
    0.171404984700515, 0.128036341067311, 0.109148560224565, 
    0.164344103597518, 0.171835957308029, 0.178019850639175, 
    0.126770975643962, 0.15612172993088, 0.12310014233588, 0.18427215654897, 
    0.176204986264325, 0.173547243987089, 0.130903852754604, 
    0.127725787316048, 0.151375091860373, 0.179945264085907, 
    0.189834190001491, 0.130580396459516, 0.173335984456374, 
    0.125435480471608, 0.184314576186854, 0.120800315709439, 
    0.196173015628708, 0.18358172736331, 0.135984461231908, 
    0.155981523178682, 0.134354566451351, 0.192457189271989, 
    0.213286255193696, 0.137141906313331, 0.174419436369902, 
    0.134747389131557, 0.177906011191179, 0.127593617173957, 
    0.188946197511486, 0.2003258058779, 0.141387771187489, 0.174471591302939, 
    0.131149743454265, 0.198898887094371, 0.111413908850674, 
    0.229361462292454, 0.14757731753431, 0.183833497382841, 
    0.145608789845189, 0.164105325834176, 0.14647705355381, 
    0.168893903303636, 0.21279306882401, 0.144506790450027, 
    0.169930653567971, 0.139393742478665, 0.200723049149477, 
    0.108039058459723, 0.235911675494728, 0.159236916386634, 
    0.202126190399384, 0.150087874947255, 0.130759577328282, 
    0.158447413422126, 0.152873223372957, 0.0867883385720827, 
    0.217450887006753, 0.148472017344834, 0.167502181064347, 
    0.150592866691246, 0.188429626976068, 0.112689401577857, 0.2316305351423, 
    0.16716879307099, 0.214625496802526, 0.146595718672683, 
    0.0887384103705287, 0.148015362405907, 0.150352481363271, 
    0.0923169915991004, 0.227306005377937, 0.151147851548721, 
    0.181857037975724, 0.152515036510108, 0.152791794382232, 
    0.097626915106148, 0.21784515754257, 0.175607888751122, 
    0.0768635644021609, 0.213144551557534, 0.145429414805772, 
    0.0591345235840816, 0.137063634491517, 0.154285576316962, 
    0.0982554816898909, 0.236893961070653, 0.150344228945373, 
    0.198697856801141, 0.143992565215689, 0.11336875028027, 
    0.0678875739619216, 0.20024688042595, 0.191890905029911, 
    0.0826006524877724, 0.214859411139656, 0.142434625230361, 
    0.0408866853814332, 0.143608556730717, 0.152950605022543, 
    0.0798086852914453, 0.236912834747342, 0.151399295782453, 
    0.0844769135886295, 0.199059280511541, 0.13649857726566, 
    0.0904039626149169, 0.054833184914719, 0.181314832557419, 
    0.203360231123154, 0.0876878547367659, 0.224868661998387, 
    0.136521902285216, 0.0313668759942612, 0.157551731513166, 
    0.143161799241976, 0.0448863754235078, 0.227482082648751, 
    0.161822631885461, 0.0843065941059268, 0.19076073107741, 
    0.129524722250593, 0.077314663230628, 0.0600347162776729, 
    0.169021413559023, 0.199461185237027, 0.0732850952035547, 
    0.234648125274686, 0.13494849011839, 0.0857869061906988, 
    0.045490407671542, 0.158706001903253, 0.127696221619965, 
    0.0335974282708369, 0.208846818227487, 0.173393123072065, 
    0.0857374772630198, 0.194658132897222, 0.1238608864997, 
    0.0723668448102527, 0.0667710625878339, 0.162148670409668, 
    0.187840206390679, 0.0451798019371798, 0.236331112189767, 
    0.140228546192102, 0.0885896922599249, 0.0723596192357564, 
    0.149731236287278, 0.112521201061473, 0.0491173789061043, 
    0.187714857740232, 0.179261985413747, 0.0779430055298373, 
    0.21149088844508, 0.124747954069233, 0.0877922016380722, 
    0.0957436113508148, 0.0716862463378918, 0.145759478285662, 
    0.166482136479877, 0.0388148660149774, 0.222461625356393, 
    0.146043422144331, 0.0927576457934852, 0.094395577686176, 
    0.152338314205216, 0.106802271324462, 0.0660189901140265, 
    0.167860888525907, 0.182138687231461, 0.0625148668043827, 
    0.223265285803411, 0.126146296391452, 0.0937729357053701, 
    0.130197392459757, 0.0805622451543081, 0.10486465234704, 
    0.133694999464701, 0.0590632102049324, 0.195817732496092, 
    0.152449699036794, 0.0851876232528266, 0.11309593872781, 
    0.171517987257798, 0.108693977565871, 0.0885101276634629, 
    0.0722875130311398, 0.141939073110885, 0.165418796214676, 
    0.0580573293761953, 0.213639994441002, 0.122421042522264, 
    0.101915876695454, 0.144648333335375, 0.0933086358163868, 
    0.0568254044936266, 0.112786384096192, 0.0816832052019172, 
    0.163785571143094, 0.161106735327164, 0.0649399319516154, 
    0.131719700648381, 0.187228621414072, 0.103242802065824, 
    0.0991830919553701, 0.07461505596538, 0.092007252787039, 
    0.127512181128934, 0.0699976979083551, 0.187407783709607, 
    0.122632612956361, 0.0875321944868269, 0.141514740519587, 0.103262539826, 
    0.0247494439936839, 0.0873945934217513, 0.121148197250351, 
    0.0874974739686398, 0.125611711050338, 0.152932681712723, 
    0.05607569562586, 0.138169020515048, 0.182391995823147, 
    0.0882332081114841, 0.106815016099751, 0.081241909273943, 
    0.0284309582010843, 0.106241530373731, 0.0862088489111991, 
    0.15801593552704, 0.128883398291666, 0.0545201248269491, 
    0.141259482681558, 0.109791761218426, 0.0043857125965379, 
    0.101596832508043, 0.138820465726932, 0.0793458909263174, 
    0.0691428729042265, 0.121878483619169, 0.0592021209211985, 
    0.123216973194215, 0.163126032650346, 0.0820159000542423, 
    0.0873385604536237, 0.0875045596214472, -0.0163261241250303, 
    0.0865503211102296, 0.11820711185942, 0.0917400671408126, 
    0.122703309875294, 0.126858893801642, 0.0347760667238501, 
    0.146201844540412, 0.11571216639536, -0.0113855810564673, 
    0.105144170970055, 0.128169492304487, 0.0762069666469898, 
    0.00509080927530317, 0.105487135842481, 0.0531266274054616, 
    0.0813687791182764, 0.143862095678848, 0.0925961796155693, 
    0.0478868240456991, 0.0909667081392817, -0.0353075618210043, 
    0.110544291129836, 0.131853806605533, 0.0807901147161291, 
    0.0680032705573078, 0.110105537993245, 0.0258587298121571, 
    0.143089549416845, 0.12066470034339, -0.00337777752377674, 
    0.0859380609457383, 0.0797405364228571, 0.0809657107444941, 
    -0.0353269786172177, 0.0902749823574875, 0.122717152142623, 
    0.0472141807872889, 0.0256529024835687, 0.123127309200045, 
    0.0999163246174781, 0.0110716905031469, 0.0974074177763509, 
    -0.0427439984620037, 0.116192917433645, 0.101177705856158, 
    0.0709501347177028, 0.00708054447174309, 0.103176928253667, 
    0.00288715673934535, 0.121676799412608, 0.115205335007285, 
    0.0346594722523939, 0.0499760540532925, 0.0365795248771256, 
    0.0836827725924067, -0.0475048274460043, 0.116136475570454, 
    0.134353806605533, 0.0550519565523709, -0.0327576762995762, 
    0.0847338799894805, 0.0978918201274395, -0.0262031903538584, 
    0.103050625445822, -0.0328043284932975, 0.104838915039341, 
    0.0214630267708272, 0.072262670526513, -0.0280061768495358, 
    0.0982942389492844, 0.120076443514089, -0.0119601807331553, 
    0.0891109471919628, 0.102423887151548, 0.0603047542551269, 
    -0.000356833527703779, 0.0261639717736745, 0.079810982229476, 
    -0.048591471606535, 0.126089091531774, 0.0846135273893609, 
    0.062403282122079, -0.0792766629615696, 0.034422630033488, 
    0.0997354882198928, -0.0704632155751079, 0.0932669119663942, 
    0.00293418471060767, 0.08249379924541, -0.0443960438569357, 
    0.070147624548214, -0.0344510945689051, 0.11726837254311, 
    0.120688343814853, 0.00713949688739561, 0.0491508383795209, 
    0.0875812806660259, 0.0547112517308683, -0.0684239082552415, 
    0.0391179158937507, 0.0676342130923061, -0.0390079417745474, 
    0.111504138091401, -0.0235919048697978, 0.0631233548202655, 
    -0.0997268451033869, 0.00147501256170948, 0.11451068805994, 
    0.106330539959121, -0.0875633606647959, 0.0628643093255001, 
    0.0273970288749848, 0.0286421405015813, -0.0629875009979665, 
    0.0469654823300767, -0.0271670642487514, 0.122992778055211, 
    0.0579111087031687, 0.0364946066367782, 0.0037758445502225, 
    0.0682237510848011, 0.0450187663398328, -0.132511338207424, 
    0.0672459627969688, 0.0404223685093629, -0.0145458262757206, 
    0.086350184406845, -0.113008714755373, 0.0523752407370296, 
    -0.0845728595157573, -0.00510338749735029, 0.112414265012941, 
    0.0839710535073439, -0.0543412160032293, 0.0228331042071658, 
    0.0159090412786291, -0.0641597412089065, -0.0496573356733888, 
    0.00727040264603179, -0.00987128466090484, 0.102806170562104, 
    -0.0521070330618309, 0.0540855733640889, -0.0323412064852972, 
    0.0465286841958633, 0.108692204430391, 0.0355219813041529, 
    -0.148670524816478, 0.10244819846972, -0.00865348242254689, 
    -0.00110089592970274, 0.0456877651649693, -0.141683179708904, 
    0.0184618434508156, -0.0472321368674927, 0.0063137824839318, 
    0.0985993194000374, 0.0103157138925369, -0.00119124541400305, 
    -0.00793274303730017, -0.00481644656039906, -0.146086526629891, 
    -0.00824544477603002, -0.0404157048700442, 0.00859601949064756, 
    0.0788007459302826, -0.141090934104238, 0.0547995564488219, 
    -0.0372972367668081, 0.0296594215337583, 0.10584583804235, 
    0.00268581028206361, -0.100510863769283, 0.13462278521669, 
    -0.0668547009686154, -0.0162216960260585, -0.0285188130124534, 
    -0.126738176737842, -0.0257239041629776, -0.0141823467545363, 
    0.0354883767690438, 0.081240094763644, -0.0782374488925752, 
    0.0389938680418233, -0.0258177585789707, 0.087059056237032, 
    -0.014469244220697, -0.165537512206547, 0.0474237098420337, 
    -0.0902950043163488, 0.0110109249605596, 0.061607870145438, 
    -0.177107318003082, 0.0350047757410135, -0.0132716386302624, 
    0.0264266635645424, 0.0903788233376498, -0.0518185283561811, 
    -0.0276863272151381, 0.141583251148766, -0.103934787715034, 
    -0.0437480261502428, -0.105492506633772, -0.0802335124029831, 
    -0.0645029395879873, 0.00714045361232655, 0.058970481945987, 
    0.0737892355615101, -0.139731878499435, 0.0593068501499937, 
    -0.0348112820127294, 0.0956956915579755, -0.0256693678795052, 
    -0.119323313106812, 0.0975146962882129, -0.131132327728079, 
    -0.00765137101703385, 0.0178704997316872, -0.171291121335519, 
    0.0113813172368638, 0.0164349507991004, 0.0502028777633764, 
    0.0821508833399804, -0.0937522188010662, 0.0287368028069366, 
    0.104673992101793, -0.115115091342642, 0.0645446962981016, 
    -0.0594275877265563, -0.132630259788553, -0.0165098533903884, 
    -0.0781640245735273, 0.00900482431161937, 0.0566905395775436, 
    0.0853433843127985, -0.172976198189294, 0.0601184537195292, 
    -0.0372045929137839, 0.0942150354958528, -0.0459441227775153, 
    -0.0424606491298663, 0.118668441214405, -0.152231759773772, 
    -0.0479802829283275, -0.0492515093193193, -0.134188986887782, 
    -0.00688120817838031, 0.0346376339784631, 0.0772892495462132, 
    0.0892446073811557, -0.112677319477987, 0.0661350270315066, 
    0.0460981865012321, -0.115495180938511, 0.0849958564573901, 
    -0.0590165358482553, -0.0991982497597393, 0.0478616811514942, 
    -0.0679126140191884, -0.0213195391593495, 0.0324155222002493, 
    0.0800877407671267, -0.182710386959751, 0.0558973084478013, 
    -0.0243751865762781, 0.0924153181544336, -0.0623639870786972, 
    0.0256444373090725, 0.0912681059136325, -0.156974685471693, 
    0.0442432526016787, -0.0863495085603242, -0.0872835801010528, 
    -0.0746379596407106, -0.00348372993153055, 0.0314619602513589, 
    0.0763240161044408, 0.115756052067633, -0.123014332169004, 
    0.087461473912577, 0.0171020012619889, -0.115217135638393, 
    0.0943319729489141, -0.0536974186759529, -0.0299716446577413, 
    0.0873708337925302, -0.0617708531230524, -0.0642068845896527, 
    -0.0256830125137786, 0.0398348647067075, -0.16062103384361, 
    0.0547435476809949, -0.00218490243992556, 0.102168801717093, 
    -0.0746326931352005, 0.0696240140900393, 0.0361023937316997, 
    -0.156588936444514, 0.0766140099947058, -0.0941911084231147, 
    -0.0698757399941144, -0.0041565169607127, 0.0114747161845069, 
    -0.00166988432033166, 0.0470633139099867, 0.133121813092228, 
    -0.135755911670089, 0.0972992082776693, 0.025367814177696, 
    -0.107716251029403, 0.0938964991747171, -0.0492876626158066, 
    0.0351160162440884, 0.0782845548882419, -0.0739068850083846, 
    0.0451003387833193, -0.0822611611723553, -0.0931158496226017, 
    0.00290822841658495, -0.110825776895376, 0.0705999797852665, 
    0.0108462488488515, 0.126484659245367, -0.0881312490903048, 
    0.0904203706390785, 0.00432910888308123, -0.156352876138038, 
    0.0916500175663526, -0.0839965545439225, -0.0112840531050068, 
    0.0534895375357919, 0.0119623327935335, -0.0437916963033693, 
    -0.0128314106110337, 0.118064631001535, -0.135365014364471, 
    0.105820566910339, 0.0303113309508253, -0.090912319432113, 
    0.0985504419044934, -0.0537791164750444, 0.0665977201146679, 
    0.0363779674621684, -0.0985074491212009, 0.0775267907564246, 
    -0.0590928170494807, -0.121592024627609, 0.00320159649008188, 
    -0.0492773873818161, 0.0829020233134131, 0.00630694131050501, 
    0.140084245953556, -0.105636481150035, 0.100390246117452, 
    0.00586701652535115, -0.151902667968029, 0.0887951773026146, 
    -0.07382324399899, 0.048341266488229, 0.068244658777988, 
    -0.0128724688103557, 0.047363113323875, -0.0629085949563844, 
    -0.0802930287314033, 0.0902571048188344, -0.116384511085524, 
    0.126648752006957, 0.0114029193163233, -0.0691658055945079, 
    0.110545271329771, -0.0650527883969454, 0.0707320983361994, 
    0.00494113891237812, -0.124265238415449, 0.0997931755253369, 
    -0.0340760232195748, -0.114884985838445, 0.0330085760014328, 
    0.00851530407757918, 0.0702669287407992, -0.0269274165269166, 
    0.125950983540598, -0.115375588727231, 0.111872419670727, 
    0.00227571239498797, -0.143403990408176, 0.0819018788215322, 
    -0.0693323065008059, 0.0691859159154491, 0.0433463071197936, 
    -0.0577059281873746, 0.0746690208633865, -0.0408275921421037, 
    -0.116278206421958, 0.0784395688705087, -0.0923776757681495, 
    0.13294144167469, -0.0218066954048127, -0.0483968855937918, 
    0.113467987717939, -0.0818739689430042, 0.077685164474357, 
    -0.00627012947074257, -0.137328783324833, 0.104720775447146, 
    -0.031408194516804, -0.10722624759526, 0.0611843106337311, 
    0.0380413908959471, 0.0310270673224568, 0.0429429914763443, 
    -0.0716072846559777, 0.0986280764985217, -0.103180846266031, 
    0.127499656305852, -0.0184419722232853, -0.125083343112372, 
    0.0828186431925622, -0.0632060760789571, 0.0601128966760431, 
    0.0152616110538719, -0.101177645704279, 0.103475780388158, 
    -0.0194913708219633, -0.110269104644512, 0.0730296348678434, 
    -0.0680763458217148, 0.108331268793595, -0.0462893870630766, 
    -0.0468694331284791, 0.10001094695184, -0.0980512173893402, 
    0.0910621874868995, -0.0200189043042309, -0.134384340957514, 
    0.0954110951301259, -0.100655994911529, 0.0644342654674867, 
    0.0301023922508332, -0.0277155412244841, 0.0464626084752208, 
    -0.0939884889578605, 0.0802324765853525, -0.0820614057159447, 
    0.11825483843507, -0.0391164252833186, -0.0965133672034531, 
    0.0943796587955442, -0.0645462763211706, 0.0593169393767008, 
    -0.00372496394509453, -0.121607065857804, 0.117238747188321, 
    -0.00659494731126046, -0.0922768180526139, 0.0493610247411094, 
    -0.0394109388562407, 0.0649010527927174, 0.0470744612029068, 
    -0.0577982933209897, -0.0601992036012902, 0.0760004437509048, 
    -0.0931112661879064, 0.097461671436477, -0.0373399824771916, 
    -0.120666430572616, 0.0899266449015466, -0.0855298255248363, 
    0.0505319742571117, 0.0123009718235624, -0.078818331739435, 
    0.0635239054360527, -0.0826700915261183, 0.0624542259322965, 
    -0.0654251758671661, 0.0928283767129976, -0.0485401082541421, 
    -0.0728342728924371, 0.104125342713045, -0.0765212843132895, 
    0.062116264635337, -0.0215230318639828, -0.121052149857672, 
    0.107122070647712, -0.0808185485290903, 0.0241674585061501, 
    -0.0283505123595164, 0.013115699371735, 0.0471599351353772, 
    -0.0579774533606919, -0.0634902894949699, 0.0561753245644529, 
    -0.075071964797976, 0.0806043962903054, -0.0417650458887874, 
    -0.104631442957508, 0.101629414654919, -0.0753886007534449, 
    0.032221250078498, -0.000405695948841567, -0.103545847596085, 
    0.080606179072071, -0.0655681105121444, 0.0252785357274377, 
    -0.0418366731985671, 0.0677628815662848, 0.0561708333513106, 
    -0.0512248567972115, -0.0603253751146246, 0.0897112953039367, 
    -0.0759711341372464, 0.0515891738778832, -0.0352952181302211, 
    -0.110107371796993, 0.0914246077238198, -0.0793116610088547, 
    0.00509556585513413, -0.0222581016959416, -0.0306198798793254, 
    0.0578433634438653, -0.0601279632789866, -0.0489535082741651, 
    0.0379165200751214, -0.0617356006718536, 0.0595897114761648, 
    -0.0351479268576577, -0.0918230142931075, 0.115713324890779, 
    -0.0742024972307032, -0.00451520679631327, -0.0129953073378032, 
    -0.112458247269781, 0.0772561712140156, -0.054254926984503, 
    -0.0104388647360375, -0.0381190125374193, 0.0475851941609274, 
    0.0648227360730963, -0.0553467626832331, -0.0481572567174697, 
    0.0549484492434983, -0.0662620484143279, 0.0262786821789773, 
    -0.0340355222636342, -0.0986273186992354, 0.0919527307374278, 
    -0.0888884969391996, -0.0368089544357442, -0.00855709039348918, 
    -0.06051214740023, 0.0683086632029305, -0.0441578932269881, 
    0.00611219044757472, -0.0405123628958326, 0.0396490554823868, 
    0.0607050318292112, -0.0285962252054147, -0.0800466585496452, 
    0.100564414200421, -0.065254214730441, -0.0538084718701733, 
    -0.0269573087881189, -0.115000102509884, 0.0594321893330042, 
    -0.0494825705901361, -0.0428603667620533, -0.0371225399576368, 
    0.0252654015981332, 0.0738909241637195, -0.0312148580698463, 
    0.0231099644158261, -0.0614565443709571, 0.00793779497225861, 
    -0.0871360126582197, 0.0983612821830744, -0.0885137032311289, 
    -0.11241765224717, -0.00482759404121512, -0.0816066720367744, 
    0.0618237371319845, -0.0494642775704404, -0.0291099553420813, 
    -0.041579095545232, 0.0171400240115436, 0.0793543138789188, 
    -0.04312187865003, -0.062598610911551, 0.0561245967044358, 
    -0.0636566680781261, -0.0901600707468136, -0.0238467158000905, 
    -0.114260405857439, 0.0398099496535075, -0.0618802533535043, 
    -0.10155657406465, -0.00231511464995466, 0.0752103395041276, 
    -0.0346209128235062, -0.00555256005541232, -0.00588988494730074, 
    0.0617130274346799, -0.0746344066706165, 0.085219581594417, 
    -0.0730055287317548, -0.181868665732583, -0.0201383198567652, 
    -0.100194159618408, 0.0435390924091762, -0.0496797141448236, 
    -0.0712715910659562, -0.0459450192056837, -0.00512280424802208, 
    0.0904346784832138, -0.0315532525673187, 0.011906351134576, 
    -0.0710545299555481, -0.103538540338852, -0.101514979943376, 
    0.0212286645638935, -0.0734358490497304, -0.175986530420999, 
    -0.0273520785551247, 0.0618023482476705, -0.0540322166007847, 
    -0.0373300719759971, -0.0241287442990032, 0.0731079759882938, 
    -0.0537708316889471, 0.0472603387103085, -0.0771601349940996, 
    -0.206448217307488, -0.0414527756968616, -0.117953400129699, 
    0.0217546823195233, -0.0600481305507701, -0.137240157636851, 
    -0.0186133546757973, 0.0894358804898526, -0.00707893914496135, 
    -0.0216437160612717, -0.110231052729149, 0.0661062801665477, 
    -0.0750534130182729, 0.0153462353453495, -0.0804836743062159, 
    -0.22445579341813, -0.0485537285080542, 0.0391506285877051, 
    -0.062358754884781, -0.0766131918867235, -0.0399009414550534, 
    0.0768072065593857, -0.0190246638337283, 0.00104761682208946, 
    -0.20963326814997, -0.115973980603232, -0.000230380846262968, 
    -0.073180111745043, -0.196900435633527, -0.0303901257098735, 
    0.0732596012807356, -0.00216163807914405, -0.0516093993685752, 
    -0.111234273878351, 0.0669357297982892, -0.0379238163080876, 
    0.0153549194080557, -0.234828802024284, -0.0795200613045014, 
    0.0129960244731884, -0.0694401887736173, -0.110563325840431, 
    -0.0410834474492346, 0.07410568029454, 0.00501187493042585, 
    -0.0394435209303991, -0.213467509547701, 0.04738910583934, 
    -0.0818239983326247, -0.0105694445862912, -0.218286905968869, 
    -0.0453567465974659, 0.0372830154731377, -0.0398499540621203, 
    -0.0805440085371141, -0.09604428187144, 0.0592069551085165, 
    0.00540053758228723, -0.00213913836414011, -0.234195493491767, 
    -0.105657707207722, -0.0127546729834938, -0.116740936965002, 
    -0.0445933117450299, 0.0607280155873761, 0.00948237365536357, 
    -0.068769039786403, -0.194103833113895, 0.0294459724632242, 
    -0.0325641742249566, -0.0143572998302256, -0.222505603441136, 
    -0.0655928233039834, -0.0135563355479066, -0.0680276194103311, 
    -0.0925822162212905, -0.0709864009027309, 0.0499526799382996, 
    0.0180735509558164, -0.0341801347563096, -0.233404643336763, 
    0.015891760868637, -0.101563514161697, -0.0332699645426877, 
    -0.107200558488745, -0.0516683921052784, 0.0250982620551691, 
    -0.0331732885190191, -0.0864938165814718, -0.142364668398839, 
    0.0134907582939958, 0.00871474730410384, -0.0250799647801557, 
    -0.225816930904478, -0.0772651382873746, -0.0596697344206046, 
    -0.077671570509924, -0.0687157018440337, 0.0357568459302097, 
    0.00578745788387907, -0.0631311749106654, -0.205259228621708, 
    -0.00343687055435381, -0.0693419519124615, -0.0487999067465645, 
    -0.107466501927213, -0.0540950205696083, -0.031648223975641, 
    -0.085651275010767, -0.0917233354560615, 0.00563703228343506, 
    0.00811851624527355, -0.0353471269438095, -0.224257195135527, 
    -0.0394003164929176, -0.0803807952760972, -0.0886116922395639, 
    -0.0610698822192139, -0.0791190760213127, 0.00327330222658251, 
    -0.090856934303305, -0.145677198916417, -0.0124504038153792, 
    -0.0287264825318385, -0.059241509549328, -0.123394422053683, 
    -0.0478713699768278, -0.0854003252409171, -0.0640463823745674, 
    -0.0789483954252614, -0.00679320724223304, -0.0200370417891714, 
    -0.0448409222251185, -0.193067683935661, -0.0641158089093891, 
    -0.0699670943549873, -0.0994220887792265, -0.0615659281967441, 
    -0.074200483490128, -0.0503374082250916, -0.108678129929549, 
    -0.0954399187080147, -0.00955797504078358, -0.052842665670481, 
    -0.133389862065907, -0.0544997838941716, -0.0473020294069567, 
    -0.118428586770814, -0.0447597575604469, -0.0961847253795878, 
    -0.032756670379454, -0.0766110236587738, -0.133800417612521, 
    -0.0671913844067424, -0.0925361874233121, -0.0747802252763389, 
    -0.056310369482163, -0.103030997313027, -0.109910885614386, 
    -0.0843931891264333, -0.0130343571445766, -0.0431450150378105, 
    -0.118170918083353, -0.0816499686934558, -0.0478851851752998, 
    -0.126514526523367, -0.04214708337839, -0.106703068273208, 
    -0.0658644481281602, -0.117897642869002, -0.0925040375199039, 
    -0.051304687237391, -0.0793981236549709, -0.0860970764213753, 
    -0.0684040502515935, -0.0483013513879497, -0.138173857655829, 
    -0.109498015530385, -0.0993097253795879, -0.0315825065610944, 
    -0.0677099996116547, -0.099573324005355, -0.0867928861482574, 
    -0.111849389327609, -0.0510423297953734, -0.0938009761158289, 
    -0.0907540319695819, -0.141494595331183, -0.0885414153836671, 
    -0.0350418427255168, -0.0751053811779882, -0.0911616407396033, 
    -0.0967851615645494, -0.148109263576494, -0.113207210373704, 
    -0.113770176427505, -0.0534245677570663, -0.119066198900008, 
    -0.10559444879555, -0.0715587891949905, -0.0915297764870021, 
    -0.0617722930091569, -0.0896706550246361, -0.0860557443100122, 
    -0.097961899733228, -0.155420561917103, -0.097659542759149, 
    -0.0263606585854969, -0.091110337675674, -0.105281942169417, 
    -0.103283975015445, -0.129861075747254, -0.11370244647679, 
    -0.113137829143173, -0.0634090612664569, -0.160351565233906, 
    -0.124258169432751, -0.0513951878471788, -0.0797831155529881, 
    -0.081634787696809, -0.114618930587339, -0.0876119973151953, 
    -0.166885036301439, -0.105836763430247, -0.0177065712723066, 
    -0.126255197038208, -0.129047207584613, -0.088965405405928, 
    -0.0992152789691814, -0.111335326921726, -0.0820888679152613, 
    -0.112317035813918, -0.0571591348406498, -0.185506175090125, 
    -0.124950148999044, -0.0326782981407527, -0.0847698530565334, 
    -0.117726115931053, -0.109513229377368, -0.0710479220348001, 
    -0.166086174504133, -0.106190135916662, -0.00549898714503639, 
    -0.162112626718784, -0.141806082030407, -0.065300064556163, 
    -0.073670190198921, -0.12047089072895, -0.100082645186949, 
    -0.0423475625007422, -0.198182655089694, -0.108794690079121, 
    -0.0103623178581545, -0.108251351823365, -0.14620636018091, 
    -0.0809954298047246, -0.0582829854442793, -0.152188293230319, 
    -0.0616822752975348, 0.00479040506824083, -0.180969171389469, 
    -0.12866520637209, -0.0388994590294244, -0.0653275283053829, 
    -0.137966897651409, -0.0900070037914307, -0.0324848422008156, 
    -0.195767822707813, 0.0106511565037822, -0.131748246835972, 
    -0.143675779190502, -0.0500729976636619, -0.0508208176853535, 
    -0.14177933189106, -0.0691792627153728, 0.0124303046471256, 
    -0.177074357197241, -0.0997279176181835, -0.0104578378776857, 
    -0.0792804623509891, -0.135188077801881, -0.0578589857129277, 
    -0.0340678975536544, -0.178308402802579, -0.0618313536666755, 
    0.0183421295276062, -0.139244165285953, -0.115445887897359, 
    -0.0309799164640545, -0.0507656886318991, -0.140562875434613, 
    -0.0684147202100926, 0.0136031741880422, -0.164364998327278, 
    -0.088164871710991, 0.0113414641209698, -0.0945613688087048, 
    -0.0999383636907906, -0.0310899959546775, -0.0447113511326191, 
    -0.156059689266054, -0.0604878564653727, 0.0155286469850242, 
    -0.129856949970678, -0.0808026589221384, -0.0216451360456972, 
    -0.0601832528044585, -0.130063260907349, -0.052650788056375, 
    -0.00133406817651547, -0.154873107063183, -0.0692880126454172, 
    0.0136993377795594, -0.0952771596858022, -0.066521104730452, 
    -0.0243763703214763, -0.0588211085537743, -0.143493163750598, 
    -0.0574373947706396, 0.00750756354198772, -0.116672279821419, 
    -0.0684350103136412, -0.0154585658831343, -0.071459339888226, 
    -0.0913746735052436, -0.0407878567659959, -0.0298455093556456, 
    -0.150254112740138, -0.0503358744081328, 0.00244499830338362, 
    -0.0847340874414644, -0.0255602361433535, -0.0744950814177398, 
    -0.13499736889067, -0.0445358588571562, -0.00906417446079648, 
    -0.112319396125683, -0.0911851429041826, -0.0148164655108956, 
    -0.0769575170512615, -0.0552895678652178, -0.0390720922941164, 
    -0.0656406592472309, -0.148151140145609, -0.0345383548174773, 
    -0.0103348436845749, -0.0760286115906381, -0.0220494472307906, 
    -0.086679829390179, -0.105920942126029, -0.0340396573031053, 
    -0.0370121869010767, -0.119055992622951, -0.0580699492469764, 
    -0.0186944368465569, -0.0772588231791748, -0.0351026057741413, 
    -0.103241497543151, -0.131093813716077, -0.0136852932346342, 
    -0.0256698568338434, -0.0818730014623406, -0.125240380221514, 
    -0.0146080304523018, -0.0913186315532146, -0.0736159553687818, 
    -0.0309754736417727, -0.0740213260504744, -0.12460652344639, 
    -0.0266134025567114, -0.0284615378207398, -0.0768928398235867, 
    -0.0263146988440646, -0.126733447620655, -0.0854163328201741, 
    0.00140215111451796, -0.0511859234733423, -0.101023918812267, 
    -0.0872945804748655, -0.00890378743249437, -0.090441959165503, 
    -0.029349889709688, -0.113083215270805, -0.104171664057874, 
    0.00118271322535027, -0.0462346137609926, -0.0886396344803627, 
    -0.0168288437579826, -0.124208270447901, -0.0417727979012361, 
    0.000162298925750664, -0.086022668823912, -0.111129968170324, 
    -0.0488647607270571, -0.0197739462680056, -0.0899918998821803, 
    -0.0281510941077366, -0.137440362316942, -0.0506873289139241, 
    0.0124512289771245, -0.0787666008340579, -0.116527666260296, 
    -0.0117794815918224, -0.105987287511847, -0.0200340176209913, 
    -0.0112219167767725, -0.12296236566143, -0.0875664313468761, 
    -0.0231964016216429, -0.0473056281652895, -0.0961197980545814, 
    -0.0283895127032951, -0.134815087487938, 0.00307110468665448, 
    -6.38382296024986e-05, -0.120124736738472, -0.140661408251265, 
    -0.022421874151389, -0.099709955161841, -0.0221447829920016, 
    -0.146126122814989, -0.0258213128493742, -0.0204647490592673, 
    -0.0853072807656986, -0.113473314453655, -0.0294917313476817, 
    -0.115254840635868, 0.010337839068462, -0.0155624338149381, 
    -0.155738202372373, -0.130892252932326, -0.0464535723222468, 
    -0.107731750791379, -0.031348766611388, -0.14495974080825, 
    0.0391899494469559, -0.0342786849511613, -0.124083324384956, 
    -0.137568299120406, -0.0364962760068579, -0.108259138461534, 
    -0.0209888553279368, -0.168811079627367, -0.0797371918078711, 
    -0.0770381260090228, -0.11271204615583, -0.0385519236532721, 
    -0.126914386534306, 0.0508284220333479, -0.0407805328303598, 
    -0.155846844950498, -0.146052470217482, -0.0484308062089656, 
    -0.116870043172654, -0.0235180431746326, -0.158780279162097, 
    -0.0132875828278238, -0.106076048836427, -0.119052149326779, 
    -0.0402897639227401, -0.118296827670518, -0.0361563395141977, 
    -0.165860945350023, -0.122886148106699, -0.0630261326008196, 
    -0.122550360673447, -0.0310896999723763, -0.131253204751859, 
    0.0184919349798425, -0.127087945537322, -0.125539427641385, 
    -0.036624870515175, -0.125029985799608, -0.0355699213182895, 
    -0.15310721397655, -0.0754947666657144, -0.0796002187583019, 
    -0.124808513011374, -0.0346357830396959, -0.106966981939024, 
    -0.135210468481689, -0.118982365206712, -0.0321226510578052, 
    -0.132410132401963, -0.0462963693333188, -0.122498169351468, 
    -0.0450098045221106, -0.0975823303029465, -0.126621566472464, 
    -0.0305199924153339, -0.101269931489404, -0.127324080293082, 
    -0.0919071751430006, -0.0389361603751569, -0.137736674632467, 
    -0.0569469865842275, -0.094687166265196, -0.0743182818509778, 
    -0.113376514624267, -0.120128285776072, -0.027154781624956, 
    -0.110837895586576, -0.104015029160364, -0.0599775108510164, 
    -0.0608907817070922, -0.140742660222464, -0.0603201279676582, 
    -0.0871430393995601, -0.119163985078238, -0.0953484145035084, 
    -0.0360702744969016, -0.122156347964998, -0.0864705959475676, 
    -0.0604223024500774, -0.0929704488153946, -0.135983693490916, 
    -0.0601844097446401, -0.0997288867975137, -0.111282332627161, 
    -0.0582630921513004, -0.0641817973697749, -0.122136860706985, 
    -0.0914323745641206, -0.12141493806665, -0.112537440382415, 
    -0.0675180976496035, -0.117168097232576, -0.106919204346005, 
    -0.0450502336848722, -0.10556512963921, -0.115464767968473, 
    -0.122155584451712, -0.139564685563659, -0.0711795045048161, 
    -0.0908263502255499, -0.117835865833938, -0.119122041312167, 
    -0.146236334223229, -0.106556749235665, -0.157312540677194, 
    -0.155190689640931, -0.0487530840266691, -0.127009511248762, 
    -0.106708664452848, -0.150703558084525, -0.177301839693579, 
    -0.0894004394874331, -0.169370220994206, -0.170146985466184, 
    -0.158204311414673, -0.0975092028489468, -0.180599283841257, 
    -0.196444079122413, -0.0785797192791569, -0.157804017935279, 
    -0.182180874009614, -0.174968543621036, -0.0882862427100893, 
    -0.184992016648503, -0.202810439644986, -0.133105488497221, 
    -0.183275144499571, -0.185725161691657, -0.0876727368572819, 
    -0.167546754751685, -0.191447358450373, -0.107570014479312, 
    -0.172513107006255, -0.18741050096419, -0.0983527185533028, 
    -0.137693501192534, -0.170734301669822, -0.100561052127719, 
    -0.154384726215119, -0.173844664808549, -0.108596930983218, 
    -0.162051741830596, -0.11261825304721, -0.12164132467203, 
    -0.162515140945505, -0.103719468875766, -0.154917165971101, 
    -0.0864605932026787, -0.168344277971129, -0.118757474238616, 
    -0.11834502907645, -0.0832122670212821, -0.170947922932055, 
    -0.0666492869762032, -0.128208841447852, -0.058881078592658, 
    -0.0600248899686703, -0.0955820169376288, -0.0415603455434485 ;

 obs_time = 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 13008.5, 
    13008.5979166667, 13008.5979166667, 13008.5979166667, 13008.5979166667, 
    13008.5979166667, 13008.5979166667, 13008.5979166667, 13008.5979166667, 
    13008.5979166667, 13008.5979166667, 13008.5979166667, 13008.5979166667, 
    13008.5979166667, 13008.5979166667, 13008.5979166667, 13008.5979166667, 
    13008.5979166667, 13008.5979166667, 13008.5979166667, 13008.5979166667, 
    13008.5979166667, 13008.5979166667, 13008.5979166667, 13008.5979166667, 
    13008.5979166667, 13008.5979166667, 13008.5979166667, 13008.5979166667, 
    13008.5979166667, 13008.5979166667, 13008.5979166667, 13008.5979166667, 
    13008.5979166667, 13008.5979166667, 13008.5979166667, 13008.5979166667, 
    13008.5979166667, 13008.5979166667, 13009.34375, 13009.34375, 
    13009.34375, 13009.34375, 13009.34375, 13009.34375, 13009.34375, 
    13009.34375, 13009.34375, 13009.34375, 13009.34375, 13009.34375, 
    13009.34375, 13009.34375, 13009.34375, 13009.34375, 13009.34375, 
    13009.34375, 13009.34375, 13009.34375, 13009.34375, 13009.34375, 
    13009.34375, 13009.34375, 13009.34375, 13009.34375, 13009.34375, 
    13009.34375, 13009.34375, 13009.34375, 13009.34375, 13009.34375, 
    13009.34375, 13009.34375, 13009.34375, 13009.34375, 13009.34375, 
    13009.34375, 13009.34375, 13009.34375, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 13009.5, 
    13009.5, 13009.5, 13009.5, 13009.8034722222, 13009.8034722222, 
    13009.8034722222, 13009.8034722222, 13009.8034722222, 13009.8034722222, 
    13009.8034722222, 13009.8034722222, 13009.8034722222, 13009.8034722222, 
    13009.8034722222, 13009.8034722222, 13009.8034722222, 13009.8034722222, 
    13009.8034722222, 13009.8034722222, 13009.8034722222, 13009.8034722222, 
    13009.8034722222, 13009.8034722222, 13009.8034722222, 13009.8034722222, 
    13009.8034722222, 13009.8034722222, 13009.8034722222, 13009.8034722222, 
    13009.8034722222, 13009.8034722222, 13009.8034722222, 13009.8034722222, 
    13009.8034722222, 13009.8034722222, 13009.8034722222, 13009.8034722222, 
    13009.8034722222, 13009.8034722222, 13009.8034722222, 13009.8034722222, 
    13009.8034722222, 13009.8034722222, 13009.8034722222, 13009.8034722222, 
    13009.8034722222, 13009.8034722222, 13009.8034722222, 13009.8034722222, 
    13010.0548611111, 13010.0548611111, 13010.0548611111, 13010.0548611111, 
    13010.0548611111, 13010.0548611111, 13010.0548611111, 13010.0548611111, 
    13010.0548611111, 13010.0548611111, 13010.0548611111, 13010.0548611111, 
    13010.0548611111, 13010.0548611111, 13010.0548611111, 13010.0548611111, 
    13010.0548611111, 13010.0548611111, 13010.0548611111, 13010.0548611111, 
    13010.0548611111, 13010.0548611111, 13010.0548611111, 13010.0548611111, 
    13010.0548611111, 13010.0548611111, 13010.0548611111, 13010.0548611111, 
    13010.0548611111, 13010.0548611111, 13010.0548611111, 13010.0548611111, 
    13010.0548611111, 13010.0548611111, 13010.0548611111, 13010.0548611111, 
    13010.0548611111, 13010.0548611111, 13010.0548611111, 13010.0548611111, 
    13010.0548611111, 13010.0548611111, 13010.0548611111, 13010.0548611111, 
    13010.0548611111, 13010.0548611111, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 
    13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.5, 13010.9763888889, 
    13010.9763888889, 13010.9763888889, 13010.9763888889, 13010.9763888889, 
    13010.9763888889, 13010.9763888889, 13010.9763888889, 13010.9763888889, 
    13010.9763888889, 13010.9763888889, 13010.9763888889, 13010.9763888889, 
    13010.9763888889, 13010.9763888889, 13010.9763888889, 13010.9763888889, 
    13010.9763888889, 13010.9763888889, 13010.9763888889, 13010.9763888889, 
    13010.9763888889, 13010.9763888889, 13010.9763888889, 13010.9763888889, 
    13010.9763888889, 13010.9763888889, 13011.0388888889, 13011.0388888889, 
    13011.0388888889, 13011.0388888889, 13011.0388888889, 13011.0388888889, 
    13011.0388888889, 13011.0388888889, 13011.0388888889, 13011.0388888889, 
    13011.0388888889, 13011.0388888889, 13011.0388888889, 13011.0388888889, 
    13011.28125, 13011.28125, 13011.28125, 13011.28125, 13011.28125, 
    13011.28125, 13011.28125, 13011.28125, 13011.28125, 13011.28125, 
    13011.28125, 13011.28125, 13011.28125, 13011.28125, 13011.28125, 
    13011.28125, 13011.28125, 13011.28125, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 13011.5, 
    13011.5, 13011.875, 13011.875, 13011.875, 13011.875, 13011.875, 
    13011.875, 13011.875, 13011.875, 13011.875, 13011.875, 13011.875, 
    13011.875, 13011.875, 13011.875, 13011.875, 13011.875, 13011.875, 
    13011.875, 13011.875, 13011.875, 13011.875, 13011.875, 13011.875, 
    13011.875, 13011.875, 13011.875, 13011.875, 13011.875, 13011.875, 
    13011.875, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 13012, 
    13012 ;

 obs_provenance = 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 7, 7, 7, 
    7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 
    7, 7, 7, 7, 7, 7, 7, 7, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 
    7, 7, 7, 7, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 
    6, 6, 6, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 
    7, 7, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 
    3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 4, 4, 4, 4, 4, 4, 4, 5, 5, 
    5, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 5, 5, 5, 5, 5, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 4, 4, 4, 4, 4, 4, 4, 
    4, 4, 5, 5, 5, 5, 5, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 
    4, 4, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1 ;
}
