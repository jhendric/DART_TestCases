netcdf \2011060311_profiler {
dimensions:
	recNum = UNLIMITED ; // (26 currently)
	beam = 3 ;
	beamNameLen = 8 ;
	level = 72 ;
	staNamLen = 6 ;
	QCcheckNum = 10 ;
	QCcheckNameLen = 60 ;
	ICcheckNum = 3 ;
	ICcheckNameLen = 72 ;
	station = 50 ;
	maxStaticIds = 50 ;
	totalIdLen = 6 ;
	nInventoryBins = 1 ;
variables:
	int nStaticIds ;
		nStaticIds:_FillValue = 0 ;
	char staticIds(maxStaticIds, totalIdLen) ;
		staticIds:_FillValue = "" ;
	int lastRecord(maxStaticIds) ;
		lastRecord:_FillValue = -1 ;
	int invTime(recNum) ;
		invTime:_FillValue = 0 ;
	int prevRecord(recNum) ;
		prevRecord:_FillValue = -1 ;
	int inventory(maxStaticIds) ;
		inventory:_FillValue = 0 ;
	int globalInventory ;
		globalInventory:_FillValue = 0 ;
	int firstOverflow ;
		firstOverflow:_FillValue = -1 ;
	int isOverflow(recNum) ;
		isOverflow:_FillValue = 0 ;
	int firstInBin(nInventoryBins) ;
		firstInBin:_FillValue = -1 ;
	int lastInBin(nInventoryBins) ;
		lastInBin:_FillValue = -1 ;
	int wmoStaNum(recNum) ;
		wmoStaNum:long_name = "WMO numeric station ID" ;
	char staName(recNum, staNamLen) ;
		staName:long_name = "Alphanumeric station name" ;
	char QCT(QCcheckNum, QCcheckNameLen) ;
		QCT:long_name = "list of possible QC checks" ;
		QCT:reference = "Data statement definitions" ;
	char ICT(ICcheckNum, ICcheckNameLen) ;
		ICT:long_name = "list of possible IC checks" ;
		ICT:reference = "Data statement definitions" ;
	float staLat(recNum) ;
		staLat:long_name = "Station latitude" ;
		staLat:units = "degree_N" ;
		staLat:_FillValue = 1.e+38f ;
		staLat:valid_range = -90.f, 90.f ;
	float staLon(recNum) ;
		staLon:long_name = "Station longitude" ;
		staLon:units = "degree_E" ;
		staLon:_FillValue = 1.e+38f ;
		staLon:valid_range = -180.f, 180.f ;
	float staElev(recNum) ;
		staElev:long_name = "Elevation above MSL" ;
		staElev:units = "meter" ;
		staElev:_FillValue = 1.e+38f ;
		staElev:valid_range = 0.f, 8000.f ;
	double timeObs(recNum) ;
		timeObs:long_name = "Time of observation" ;
		timeObs:units = "seconds since 1970-1-1 00:00:00.0" ;
		timeObs:_FillValue = 1.7e+308 ;
	float pressure(recNum) ;
		pressure:long_name = "Pressure reduced to MSL" ;
		pressure:units = "hectopascal" ;
		pressure:_FillValue = 1.e+38f ;
	float temperature(recNum) ;
		temperature:long_name = "Surface temperature" ;
		temperature:units = "kelvin" ;
		temperature:_FillValue = 1.e+38f ;
	int relHumidity(recNum) ;
		relHumidity:long_name = "Surface relative humidity" ;
		relHumidity:units = "percent" ;
		relHumidity:_FillValue = -1 ;
	float windSpeedSfc(recNum) ;
		windSpeedSfc:long_name = "Surface wind speed" ;
		windSpeedSfc:units = "meter/sec" ;
		windSpeedSfc:_FillValue = 1.e+38f ;
		windSpeedSfc:valid_range = -150.f, 150.f ;
	int windDirSfc(recNum) ;
		windDirSfc:long_name = "Surface wind direction" ;
		windDirSfc:units = "degree" ;
		windDirSfc:_FillValue = -1 ;
		windDirSfc:valid_range = 0, 360 ;
	float rainRate(recNum) ;
		rainRate:long_name = "Rainfall rate - surface" ;
		rainRate:units = "kg/meter2/sec" ;
		rainRate:_FillValue = 1.e+38f ;
	int submode(recNum) ;
		submode:long_name = "NOAA wind profiler submode information" ;
		submode:units = "in code" ;
		submode:_FillValue = -1 ;
	float levels(recNum, level) ;
		levels:long_name = "Height above station" ;
		levels:units = "meter" ;
		levels:_FillValue = 1.e+38f ;
		levels:valid_range = 0.f, 16250.f ;
	int levelMode(recNum, level) ;
		levelMode:long_name = "Wind profiler mode information" ;
		levelMode:value1 = "Data from low mode" ;
		levelMode:value2 = "Data from high mode" ;
		levelMode:value-1 = "Missing" ;
		levelMode:level = "levels" ;
		levelMode:_FillValue = -1 ;
	float uComponent(recNum, level) ;
		uComponent:long_name = "u (eastward) component" ;
		uComponent:level = "levels" ;
		uComponent:_FillValue = 1.e+38f ;
	char uComponentDD(recNum, level) ;
		uComponentDD:long_name = "U component QC summary value" ;
		uComponentDD:values = "Z,S,X,Q,G, or B" ;
		uComponentDD:reference = "Global Attributes Section" ;
	int uComponentQCA(recNum, level) ;
		uComponentQCA:long_name = "U component QC applied word" ;
		uComponentQCA:NoBitsSet = "No QC applied" ;
		uComponentQCA:Bit1Set = "Master bit - at least 1 check applied" ;
		uComponentQCA:Bit2Set = "Validity check applied" ;
		uComponentQCA:Bit3Set = "Reserved" ;
		uComponentQCA:Bit4Set = "Internal Consistency check applied" ;
		uComponentQCA:Bit5Set = "Reserved" ;
		uComponentQCA:Bit6Set = "Reserved" ;
		uComponentQCA:Bit7Set = "Reserved" ;
		uComponentQCA:Bit8Set = "Reserved" ;
		uComponentQCA:Bit9Set = "Reserved" ;
		uComponentQCA:Bit10Set = "Time-Height Consistency applied" ;
		uComponentQCA:reference = "Global Attributes Section" ;
	int uComponentQCR(recNum, level) ;
		uComponentQCR:long_name = "U component QC results word" ;
		uComponentQCR:NoBitsSet = "No QC applied" ;
		uComponentQCR:Bit1Set = "Master bit - at least 1 check failed" ;
		uComponentQCR:Bit2Set = "Validity check failed" ;
		uComponentQCR:Bit3Set = "Reserved" ;
		uComponentQCR:Bit4Set = "Internal Consistency check failed" ;
		uComponentQCR:Bit5Set = "Reserved" ;
		uComponentQCR:Bit6Set = "Reserved" ;
		uComponentQCR:Bit7Set = "Reserved" ;
		uComponentQCR:Bit8Set = "Reserved" ;
		uComponentQCR:Bit9Set = "Reserved" ;
		uComponentQCR:Bit10Set = "Time-Height Consistency failed" ;
		uComponentQCR:reference = "Global Attributes Section" ;
	int uComponentICA(recNum, level) ;
		uComponentICA:long_name = "U component IC applied word" ;
		uComponentICA:NoBitsSet = "No IC check applied" ;
		uComponentICA:Bit1Set = "Master bit - at least 1 check applied" ;
		uComponentICA:Bit2Set = "IC check 1 applied" ;
		uComponentICA:Bit3Set = "IC check 3 applied" ;
		uComponentICA:reference = "Global Attributes Section" ;
	int uComponentICR(recNum, level) ;
		uComponentICR:long_name = "U component IC results word" ;
		uComponentICR:NoBitsSet = "No IC check failures" ;
		uComponentICR:Bit1Set = "Master bit - at least 1 check failed" ;
		uComponentICR:Bit2Set = "IC check 1 failed" ;
		uComponentICR:Bit3Set = "IC check 3 failed" ;
		uComponentICR:reference = "Global Attributes Section" ;
	float vComponent(recNum, level) ;
		vComponent:long_name = "v (northward) component" ;
		vComponent:level = "levels" ;
		vComponent:_FillValue = 1.e+38f ;
	char vComponentDD(recNum, level) ;
		vComponentDD:long_name = "V component QC summary value" ;
		vComponentDD:values = "Z,S,X,Q,G, or B" ;
		vComponentDD:reference = "Global Attributes Section" ;
	int vComponentQCA(recNum, level) ;
		vComponentQCA:long_name = "V component QC applied word" ;
		vComponentQCA:NoBitsSet = "No QC applied" ;
		vComponentQCA:Bit1Set = "Master bit - at least 1 check applied" ;
		vComponentQCA:Bit2Set = "Validity check applied" ;
		vComponentQCA:Bit3Set = "Reserved" ;
		vComponentQCA:Bit4Set = "Internal Consistency check applied" ;
		vComponentQCA:Bit5Set = "Reserved" ;
		vComponentQCA:Bit6Set = "Reserved" ;
		vComponentQCA:Bit7Set = "Reserved" ;
		vComponentQCA:Bit8Set = "Reserved" ;
		vComponentQCA:Bit9Set = "Reserved" ;
		vComponentQCA:Bit10Set = "Time-Height Consistency applied" ;
		vComponentQCA:reference = "Global Attributes Section" ;
	int vComponentQCR(recNum, level) ;
		vComponentQCR:long_name = "V component QC results word" ;
		vComponentQCR:NoBitsSet = "No QC applied" ;
		vComponentQCR:Bit1Set = "Master bit - at least 1 check failed" ;
		vComponentQCR:Bit2Set = "Validity check failed" ;
		vComponentQCR:Bit3Set = "Reserved" ;
		vComponentQCR:Bit4Set = "Internal Consistency check failed" ;
		vComponentQCR:Bit5Set = "Reserved" ;
		vComponentQCR:Bit6Set = "Reserved" ;
		vComponentQCR:Bit7Set = "Reserved" ;
		vComponentQCR:Bit8Set = "Reserved" ;
		vComponentQCR:Bit9Set = "Reserved" ;
		vComponentQCR:Bit10Set = "Time-Height Consistency failed" ;
		vComponentQCR:reference = "Global Attributes Section" ;
	int vComponentICA(recNum, level) ;
		vComponentICA:long_name = "V component IC applied word" ;
		vComponentICA:NoBitsSet = "No IC check applied" ;
		vComponentICA:Bit1Set = "Master bit - at least 1 check applied" ;
		vComponentICA:Bit2Set = "IC check 1 applied" ;
		vComponentICA:Bit3Set = "IC check 3 applied" ;
		vComponentICA:reference = "Global Attributes Section" ;
	int vComponentICR(recNum, level) ;
		vComponentICR:long_name = "V component IC results word" ;
		vComponentICR:NoBitsSet = "No IC check failures" ;
		vComponentICR:Bit1Set = "Master bit - at least 1 check failed" ;
		vComponentICR:Bit2Set = "IC check 1 failed" ;
		vComponentICR:Bit3Set = "IC check 3 failed" ;
		vComponentICR:reference = "Global Attributes Section" ;
	float wComponent(recNum, level) ;
		wComponent:long_name = "w (upward) component" ;
		wComponent:level = "levels" ;
		wComponent:_FillValue = 1.e+38f ;
	int uvQualityCode(recNum, level) ;
		uvQualityCode:long_name = "NOAA wind profiler quality control test results for U and V" ;
		uvQualityCode:level = "levels" ;
		uvQualityCode:_FillValue = -1 ;
		uvQualityCode:reference = "Quality code bit table in global attributes section" ;
	byte wQualityCode(recNum, level) ;
		wQualityCode:long_name = "NOAA wind profiler quality control test results for W" ;
		wQualityCode:level = "levels" ;
		wQualityCode:_FillValue = -1b ;
		wQualityCode:reference = "Quality code bit table in global attributes section" ;
	float HorizSpStdDev(recNum, level) ;
		HorizSpStdDev:long_name = "Horizontal wind speed standard deviation" ;
		HorizSpStdDev:units = "meter/sec" ;
		HorizSpStdDev:level = "levels" ;
		HorizSpStdDev:_FillValue = 1.e+38f ;
	float VertSpStdDev(recNum, level) ;
		VertSpStdDev:long_name = "Vertical wind speed standard deviation" ;
		VertSpStdDev:units = "meter/sec" ;
		VertSpStdDev:level = "levels" ;
		VertSpStdDev:_FillValue = 1.e+38f ;
	char beamNames(beam, beamNameLen) ;
		beamNames:long_name = "Beam direction names" ;
	float azimBeam(recNum, beam) ;
		azimBeam:long_name = "Azimuth of beam" ;
		azimBeam:units = "degree" ;
		azimBeam:beam = "beamNames" ;
		azimBeam:_FillValue = 1.e+38f ;
		azimBeam:valid_range = 0.f, 360.f ;
	float elevBeam(recNum, beam) ;
		elevBeam:long_name = "Elevation of beam" ;
		elevBeam:units = "degree" ;
		elevBeam:beam = "beamNames" ;
		elevBeam:_FillValue = 1.e+38f ;
		elevBeam:valid_range = 0.f, 90.f ;
	byte momentsQualityCode(recNum, level, beam) ;
		momentsQualityCode:long_name = "NOAA wind profiler data quality control test results for moments" ;
		momentsQualityCode:level = "levels" ;
		momentsQualityCode:beam = "beamNames" ;
		momentsQualityCode:_FillValue = -1b ;
		momentsQualityCode:reference = "Quality code bit table in global attributes section" ;
	int consensusNum(recNum, level) ;
		consensusNum:long_name = "Consensus number" ;
		consensusNum:level = "levels" ;
		consensusNum:_FillValue = 2147483647 ;
	int consensusNumBeam(recNum, level, beam) ;
		consensusNumBeam:long_name = "Consensus number" ;
		consensusNumBeam:level = "levels" ;
		consensusNumBeam:beam = "beamNames" ;
		consensusNumBeam:_FillValue = 2147483647 ;
	int peakPower(recNum, level) ;
		peakPower:long_name = "Spectral peak power" ;
		peakPower:units = "dB" ;
		peakPower:level = "levels" ;
		peakPower:_FillValue = 2147483647 ;
	float peakPowerBeam(recNum, level, beam) ;
		peakPowerBeam:long_name = "Spectral peak power" ;
		peakPowerBeam:units = "dB" ;
		peakPowerBeam:level = "levels" ;
		peakPowerBeam:beam = "beamNames" ;
		peakPowerBeam:_FillValue = 1.e+38f ;
	float radVelocity(recNum, level, beam) ;
		radVelocity:long_name = "Radial velocity" ;
		radVelocity:units = "meter/sec" ;
		radVelocity:level = "levels" ;
		radVelocity:beam = "beamNames" ;
		radVelocity:_FillValue = 1.e+38f ;
	float specWidth(recNum, level, beam) ;
		specWidth:long_name = "Spectral width" ;
		specWidth:units = "meter2/sec2" ;
		specWidth:level = "levels" ;
		specWidth:beam = "beamNames" ;
		specWidth:_FillValue = 1.e+38f ;

// global attributes:
		:avgTimePeriod = "60 minutes" ;
		:staVarNum = 13 ;
		:levVarNum = 10 ;
		:nonStaticLevVar = 8 ;
		:cdlDate = "20020503" ;
		:idVariables = "staName" ;
		:timeVariables = "timeObs" ;
		:filePeriod = 3600 ;
		:fileEndOffset = 0 ;
		:qualityCodeNoBitsSet = "Good" ;
		:qualityCodeBit1Set = "Reserved" ;
		:qualityCodeBit2Set = "Test results inconclusive" ;
		:qualityCodeBit3Set = "Test B performed and failed" ;
		:qualityCodeBit4Set = "Test A performed and failed" ;
		:qualityCodeBit5Set = "Reserved" ;
		:qualityCodeBit6Set = "Reserved" ;
		:qualityCodeBit7Set = "Reserved" ;
		:qualityCodeBit8Set = "Reserved" ;
		:qualityCodeBits1To8Set = "Missing" ;
		:qualityCodeLeastSignificantBit = "bit1" ;
		:DD_long_name = "QC data descriptor model:  QC summary values" ;
		:DD_reference = "AWIPS Technique Specification Package (TSP) 88-21-R2" ;
		:DD_values = "Z,C,S,V,X,Q,G, or B" ;
		:DD_value_Z = "No QC applied" ;
		:DD_value_C = "Passed QC stage 1" ;
		:DD_value_S = "Passed QC stages 1 and 2" ;
		:DD_value_V = "Passed QC stages 1, 2 and 3" ;
		:DD_value_X = "Failed QC stage 1" ;
		:DD_value_Q = "Passed QC stage 1, but failed stages 2 or 3 " ;
		:DD_value_G = "Included in accept list" ;
		:DD_value_B = "Included in reject list" ;
		:QCStage_long_name = "automated QC checks contained in each stage" ;
		:QCStage_values = "1, 2, or 3" ;
		:QCStage_value_1 = "Validity and Position Consistency Check" ;
		:QCStage_value_2 = "Internal, Temporal, Time-Height, Vertical and Model Consistency Checks" ;
		:QCStage_value_3 = "Spatial Consistency Check" ;
		:QCStage_reference = "AWIPS TSP 88-21_R2" ;
		:QCA_long_name = "QC applied model:  applied word definition" ;
		:QCA_NoBitsSet = "No QC applied" ;
		:QCA_Bit1Set = "Master bit - at least 1 check applied" ;
		:QCA_Bit2Set = "Validity check applied" ;
		:QCA_Bit3Set = "Position Consistency check applied" ;
		:QCA_Bit4Set = "Internal Consistency check applied" ;
		:QCA_Bit5Set = "Temporal Consistency check applied" ;
		:QCA_Bit6Set = "Hydrostatic check applied" ;
		:QCA_Bit7Set = "Spatial Consistency check applied" ;
		:QCA_Bit8Set = "Super Adiabatic Lapse Rate check applied" ;
		:QCA_Bit9Set = "Wind Shear check applied" ;
		:QCA_Bit10Set = "Time-Height Consistency check applied" ;
		:QCA_LeastSignificantBit = "bit1" ;
		:QCA_reference1 = "AWIPS TSP 88-21_R2" ;
		:QCA_reference2 = "10th Met Obs and Inst, Paper FA5.7, Phoenix, 1998" ;
		:QCA_reference3 = "Ann. Geophysicae 12, 711-724 (1994)" ;
		:QCA_reference4 = "1st Int Obs Sys, Paper FA8.4, Long Beach, 1997" ;
		:QCR_long_name = "QC results model:  results word definition" ;
		:QCR_NoBitsSet = "No QC failures" ;
		:QCR_Bit1Set = "Master bit - at least 1 check failed" ;
		:QCR_Bit2Set = "Validity check failed" ;
		:QCR_Bit3Set = "Position Consistency check failed" ;
		:QCR_Bit4Set = "Internal Consistency check failed" ;
		:QCR_Bit5Set = "Temporal Consistency check failed" ;
		:QCR_Bit6Set = "Hydrostatic check failed" ;
		:QCR_Bit7Set = "Spatial Consistency check failed" ;
		:QCR_Bit8Set = "Super Adiabatic Lapse Rate check failed" ;
		:QCR_Bit9Set = "Wind Shear check failed" ;
		:QCR_Bit10Set = "Time-Height Consistency check failed" ;
		:QCR_LeastSignificantBit = "bit1" ;
		:QCR_reference1 = "AWIPS TSP 88-21_R2" ;
		:QCR_reference2 = "10th Met Obs and Inst, Paper FA5.7, Phoenix, 1998" ;
		:QCR_reference3 = "Ann. Geophysicae 12, 711-724 (1994)" ;
		:QCR_reference4 = "1st Int Obs Sys, Paper FA8.4, Long Beach, 1997" ;
		:ICA_long_name = "IC applied model:  applied word definition" ;
		:ICA_NoBitsSet = "No IC applied" ;
		:ICA_Bit1Set = "Master bit - at least 1 check applied" ;
		:ICA_BitiSet = "IC check # applied" ;
		:ICA_LeastSignificantBit = "bit1" ;
		:ICA_reference = "IC check #\'s defined in IC check table" ;
		:ICR_long_name = "IC results Model:  results word definition" ;
		:ICR_NoBitsSet = "No IC applied" ;
		:ICR_Bit1Set = "Master bit - at least 1 check applied" ;
		:ICR_BitiSet = "IC check # applied" ;
		:ICR_LeastSignificantBit = "bit1" ;
		:ICR_reference = "IC check #\'s defined in IC check table" ;
data:

 nStaticIds = 26 ;

 staticIds =
  "BLRW3",
  "CENA2",
  "CNWM7",
  "DQUA4",
  "FBYN1",
  "GDAC2",
  "GNAA2",
  "HBRK1",
  "HKLO2",
  "HVLK1",
  "LDBT2",
  "LMNO2",
  "LTHM7",
  "MBWW4",
  "NDSK1",
  "NLGN1",
  "OKOM6",
  "PLTC2",
  "PRCO2",
  "SLAI4",
  "TCUN5",
  "TLKA2",
  "WDLM5",
  "WLCI3",
  "WNFL1",
  "WSMN5",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "",
  "" ;

 lastRecord = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 
    18, 19, 20, 21, 22, 23, 24, 25, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _ ;

 invTime = 1307098800, 1307098800, 1307098800, 1307098800, 1307098800, 
    1307098800, 1307098800, 1307098800, 1307098800, 1307098800, 1307098800, 
    1307098800, 1307098800, 1307098800, 1307098800, 1307098800, 1307098800, 
    1307098800, 1307098800, 1307098800, 1307098800, 1307098800, 1307098800, 
    1307098800, 1307098800, 1307098800 ;

 prevRecord = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _ ;

 inventory = 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _ ;

 globalInventory = 1 ;

 firstOverflow = _ ;

 isOverflow = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _ ;

 firstInBin = 0 ;

 lastInBin = 25 ;

 wmoStaNum = 74357, 70197, 74550, 74752, 74440, 74530, 70268, 74546, 74648, 
    74541, 72246, 74647, 74551, 74431, 74542, 74445, 74769, 74533, 74649, 
    74449, 74731, 70252, 74341, 74466, 74753, 74629 ;

 staName =
  "BLRW3",
  "CENA2",
  "CNWM7",
  "DQUA4",
  "FBYN1",
  "GDAC2",
  "GNAA2",
  "HBRK1",
  "HKLO2",
  "HVLK1",
  "LDBT2",
  "LMNO2",
  "LTHM7",
  "MBWW4",
  "NDSK1",
  "NLGN1",
  "OKOM6",
  "PLTC2",
  "PRCO2",
  "SLAI4",
  "TCUN5",
  "TLKA2",
  "WDLM5",
  "WLCI3",
  "WNFL1",
  "WSMN5" ;

 QCT =
  "1- Validity Check",
  "2- Position Consistency Check",
  "3- Internal Consistency Check",
  "4- Temporal Consistency Check",
  "5- Hydrostatic Check",
  "6- Spatial Consistency Check",
  "7- Super Adiabatic Lapse Rate Check",
  "8- Wind Shear Check",
  "9- Time-Height Consistency Check",
  "" ;

 ICT =
  "1-Bird contamination check",
  "2-Signal strength check",
  "3-Alaska interference check" ;

 staLat = 43.22, 65.5, 37.52, 34.11, 40.08, 37.77, 62.11, 38.3, 35.68, 37.65, 
    30.09, 36.69, 39.57, 41.9, 37.3, 42.2, 34.08, 40.18, 34.97, 41.9, 35.08, 
    62.31, 44.67, 40.81, 31.89, 32.4 ;

 staLon = -90.53, -144.68, -92.7, -94.29, -97.31, -102.17, -145.97, -97.29, 
    -95.86, -99.11, -96.78, -97.48, -94.18, -106.18, -95.6, -97.79, -88.86, 
    -104.73, -97.51, -93.69, -103.6, -150.42, -95.44, -87.05, -92.78, -106.34 ;

 staElev = 226, 259, 390, 195, 433, 1155, 564, 447, 219, 648, 122, 306, 297, 
    1997, 265, 524, 125, 1524, 331, 315, 1241, 137, 319, 212, 93, 1224 ;

 timeObs = 1307098800, 1307098800, 1307098800, 1307098800, 1307098800, 
    1307098800, 1307098800, 1307098800, 1307098800, 1307098800, 1307098800, 
    1307098800, 1307098800, 1307098800, 1307098800, 1307098800, 1307098800, 
    1307098800, 1307098800, 1307098800, 1307098800, 1307098800, 1307098800, 
    1307098800, 1307098800, 1307098800 ;

 pressure = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _ ;

 temperature = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _ ;

 relHumidity = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _ ;

 windSpeedSfc = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _ ;

 windDirSfc = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _ ;

 rainRate = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _ ;

 submode = _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _ ;

 levels =
  500, 750, 1000, 1250, 1500, 1750, 2000, 2250, 2500, 2750, 3000, 3250, 3500, 
    3750, 4000, 4250, 4500, 4750, 5000, 5250, 5500, 5750, 6000, 6250, 6500, 
    6750, 7000, 7250, 7500, 7750, 8000, 8250, 8500, 8750, 9000, 9250, 7500, 
    7750, 8000, 8250, 8500, 8750, 9000, 9250, 9500, 9750, 10000, 10250, 
    10500, 10750, 11000, 11250, 11500, 11750, 12000, 12250, 12500, 12750, 
    13000, 13250, 13500, 13750, 14000, 14250, 14500, 14750, 15000, 15250, 
    15500, 15750, 16000, 16250,
  500, 750, 1000, 1250, 1500, 1750, 2000, 2250, 2500, 2750, 3000, 3250, 3500, 
    3750, 4000, 4250, 4500, 4750, 5000, 5250, 5500, 5750, 6000, 6250, 6500, 
    6750, 7000, 7250, 7500, 7750, 8000, 8250, 8500, 8750, 9000, 9250, 7500, 
    7750, 8000, 8250, 8500, 8750, 9000, 9250, 9500, 9750, 10000, 10250, 
    10500, 10750, 11000, 11250, 11500, 11750, 12000, 12250, 12500, 12750, 
    13000, 13250, 13500, 13750, 14000, 14250, 14500, 14750, 15000, 15250, 
    15500, 15750, 16000, 16250,
  500, 750, 1000, 1250, 1500, 1750, 2000, 2250, 2500, 2750, 3000, 3250, 3500, 
    3750, 4000, 4250, 4500, 4750, 5000, 5250, 5500, 5750, 6000, 6250, 6500, 
    6750, 7000, 7250, 7500, 7750, 8000, 8250, 8500, 8750, 9000, 9250, 7500, 
    7750, 8000, 8250, 8500, 8750, 9000, 9250, 9500, 9750, 10000, 10250, 
    10500, 10750, 11000, 11250, 11500, 11750, 12000, 12250, 12500, 12750, 
    13000, 13250, 13500, 13750, 14000, 14250, 14500, 14750, 15000, 15250, 
    15500, 15750, 16000, 16250,
  500, 750, 1000, 1250, 1500, 1750, 2000, 2250, 2500, 2750, 3000, 3250, 3500, 
    3750, 4000, 4250, 4500, 4750, 5000, 5250, 5500, 5750, 6000, 6250, 6500, 
    6750, 7000, 7250, 7500, 7750, 8000, 8250, 8500, 8750, 9000, 9250, 7500, 
    7750, 8000, 8250, 8500, 8750, 9000, 9250, 9500, 9750, 10000, 10250, 
    10500, 10750, 11000, 11250, 11500, 11750, 12000, 12250, 12500, 12750, 
    13000, 13250, 13500, 13750, 14000, 14250, 14500, 14750, 15000, 15250, 
    15500, 15750, 16000, 16250,
  500, 750, 1000, 1250, 1500, 1750, 2000, 2250, 2500, 2750, 3000, 3250, 3500, 
    3750, 4000, 4250, 4500, 4750, 5000, 5250, 5500, 5750, 6000, 6250, 6500, 
    6750, 7000, 7250, 7500, 7750, 8000, 8250, 8500, 8750, 9000, 9250, 7500, 
    7750, 8000, 8250, 8500, 8750, 9000, 9250, 9500, 9750, 10000, 10250, 
    10500, 10750, 11000, 11250, 11500, 11750, 12000, 12250, 12500, 12750, 
    13000, 13250, 13500, 13750, 14000, 14250, 14500, 14750, 15000, 15250, 
    15500, 15750, 16000, 16250,
  500, 750, 1000, 1250, 1500, 1750, 2000, 2250, 2500, 2750, 3000, 3250, 3500, 
    3750, 4000, 4250, 4500, 4750, 5000, 5250, 5500, 5750, 6000, 6250, 6500, 
    6750, 7000, 7250, 7500, 7750, 8000, 8250, 8500, 8750, 9000, 9250, 7500, 
    7750, 8000, 8250, 8500, 8750, 9000, 9250, 9500, 9750, 10000, 10250, 
    10500, 10750, 11000, 11250, 11500, 11750, 12000, 12250, 12500, 12750, 
    13000, 13250, 13500, 13750, 14000, 14250, 14500, 14750, 15000, 15250, 
    15500, 15750, 16000, 16250,
  500, 750, 1000, 1250, 1500, 1750, 2000, 2250, 2500, 2750, 3000, 3250, 3500, 
    3750, 4000, 4250, 4500, 4750, 5000, 5250, 5500, 5750, 6000, 6250, 6500, 
    6750, 7000, 7250, 7500, 7750, 8000, 8250, 8500, 8750, 9000, 9250, 7500, 
    7750, 8000, 8250, 8500, 8750, 9000, 9250, 9500, 9750, 10000, 10250, 
    10500, 10750, 11000, 11250, 11500, 11750, 12000, 12250, 12500, 12750, 
    13000, 13250, 13500, 13750, 14000, 14250, 14500, 14750, 15000, 15250, 
    15500, 15750, 16000, 16250,
  500, 750, 1000, 1250, 1500, 1750, 2000, 2250, 2500, 2750, 3000, 3250, 3500, 
    3750, 4000, 4250, 4500, 4750, 5000, 5250, 5500, 5750, 6000, 6250, 6500, 
    6750, 7000, 7250, 7500, 7750, 8000, 8250, 8500, 8750, 9000, 9250, 7500, 
    7750, 8000, 8250, 8500, 8750, 9000, 9250, 9500, 9750, 10000, 10250, 
    10500, 10750, 11000, 11250, 11500, 11750, 12000, 12250, 12500, 12750, 
    13000, 13250, 13500, 13750, 14000, 14250, 14500, 14750, 15000, 15250, 
    15500, 15750, 16000, 16250,
  500, 750, 1000, 1250, 1500, 1750, 2000, 2250, 2500, 2750, 3000, 3250, 3500, 
    3750, 4000, 4250, 4500, 4750, 5000, 5250, 5500, 5750, 6000, 6250, 6500, 
    6750, 7000, 7250, 7500, 7750, 8000, 8250, 8500, 8750, 9000, 9250, 7500, 
    7750, 8000, 8250, 8500, 8750, 9000, 9250, 9500, 9750, 10000, 10250, 
    10500, 10750, 11000, 11250, 11500, 11750, 12000, 12250, 12500, 12750, 
    13000, 13250, 13500, 13750, 14000, 14250, 14500, 14750, 15000, 15250, 
    15500, 15750, 16000, 16250,
  500, 750, 1000, 1250, 1500, 1750, 2000, 2250, 2500, 2750, 3000, 3250, 3500, 
    3750, 4000, 4250, 4500, 4750, 5000, 5250, 5500, 5750, 6000, 6250, 6500, 
    6750, 7000, 7250, 7500, 7750, 8000, 8250, 8500, 8750, 9000, 9250, 7500, 
    7750, 8000, 8250, 8500, 8750, 9000, 9250, 9500, 9750, 10000, 10250, 
    10500, 10750, 11000, 11250, 11500, 11750, 12000, 12250, 12500, 12750, 
    13000, 13250, 13500, 13750, 14000, 14250, 14500, 14750, 15000, 15250, 
    15500, 15750, 16000, 16250,
  500, 750, 1000, 1250, 1500, 1750, 2000, 2250, 2500, 2750, 3000, 3250, 3500, 
    3750, 4000, 4250, 4500, 4750, 5000, 5250, 5500, 5750, 6000, 6250, 6500, 
    6750, 7000, 7250, 7500, 7750, 8000, 8250, 8500, 8750, 9000, 9250, 7500, 
    7750, 8000, 8250, 8500, 8750, 9000, 9250, 9500, 9750, 10000, 10250, 
    10500, 10750, 11000, 11250, 11500, 11750, 12000, 12250, 12500, 12750, 
    13000, 13250, 13500, 13750, 14000, 14250, 14500, 14750, 15000, 15250, 
    15500, 15750, 16000, 16250,
  500, 750, 1000, 1250, 1500, 1750, 2000, 2250, 2500, 2750, 3000, 3250, 3500, 
    3750, 4000, 4250, 4500, 4750, 5000, 5250, 5500, 5750, 6000, 6250, 6500, 
    6750, 7000, 7250, 7500, 7750, 8000, 8250, 8500, 8750, 9000, 9250, 7500, 
    7750, 8000, 8250, 8500, 8750, 9000, 9250, 9500, 9750, 10000, 10250, 
    10500, 10750, 11000, 11250, 11500, 11750, 12000, 12250, 12500, 12750, 
    13000, 13250, 13500, 13750, 14000, 14250, 14500, 14750, 15000, 15250, 
    15500, 15750, 16000, 16250,
  500, 750, 1000, 1250, 1500, 1750, 2000, 2250, 2500, 2750, 3000, 3250, 3500, 
    3750, 4000, 4250, 4500, 4750, 5000, 5250, 5500, 5750, 6000, 6250, 6500, 
    6750, 7000, 7250, 7500, 7750, 8000, 8250, 8500, 8750, 9000, 9250, 7500, 
    7750, 8000, 8250, 8500, 8750, 9000, 9250, 9500, 9750, 10000, 10250, 
    10500, 10750, 11000, 11250, 11500, 11750, 12000, 12250, 12500, 12750, 
    13000, 13250, 13500, 13750, 14000, 14250, 14500, 14750, 15000, 15250, 
    15500, 15750, 16000, 16250,
  500, 750, 1000, 1250, 1500, 1750, 2000, 2250, 2500, 2750, 3000, 3250, 3500, 
    3750, 4000, 4250, 4500, 4750, 5000, 5250, 5500, 5750, 6000, 6250, 6500, 
    6750, 7000, 7250, 7500, 7750, 8000, 8250, 8500, 8750, 9000, 9250, 7500, 
    7750, 8000, 8250, 8500, 8750, 9000, 9250, 9500, 9750, 10000, 10250, 
    10500, 10750, 11000, 11250, 11500, 11750, 12000, 12250, 12500, 12750, 
    13000, 13250, 13500, 13750, 14000, 14250, 14500, 14750, 15000, 15250, 
    15500, 15750, 16000, 16250,
  500, 750, 1000, 1250, 1500, 1750, 2000, 2250, 2500, 2750, 3000, 3250, 3500, 
    3750, 4000, 4250, 4500, 4750, 5000, 5250, 5500, 5750, 6000, 6250, 6500, 
    6750, 7000, 7250, 7500, 7750, 8000, 8250, 8500, 8750, 9000, 9250, 7500, 
    7750, 8000, 8250, 8500, 8750, 9000, 9250, 9500, 9750, 10000, 10250, 
    10500, 10750, 11000, 11250, 11500, 11750, 12000, 12250, 12500, 12750, 
    13000, 13250, 13500, 13750, 14000, 14250, 14500, 14750, 15000, 15250, 
    15500, 15750, 16000, 16250,
  500, 750, 1000, 1250, 1500, 1750, 2000, 2250, 2500, 2750, 3000, 3250, 3500, 
    3750, 4000, 4250, 4500, 4750, 5000, 5250, 5500, 5750, 6000, 6250, 6500, 
    6750, 7000, 7250, 7500, 7750, 8000, 8250, 8500, 8750, 9000, 9250, 7500, 
    7750, 8000, 8250, 8500, 8750, 9000, 9250, 9500, 9750, 10000, 10250, 
    10500, 10750, 11000, 11250, 11500, 11750, 12000, 12250, 12500, 12750, 
    13000, 13250, 13500, 13750, 14000, 14250, 14500, 14750, 15000, 15250, 
    15500, 15750, 16000, 16250,
  500, 750, 1000, 1250, 1500, 1750, 2000, 2250, 2500, 2750, 3000, 3250, 3500, 
    3750, 4000, 4250, 4500, 4750, 5000, 5250, 5500, 5750, 6000, 6250, 6500, 
    6750, 7000, 7250, 7500, 7750, 8000, 8250, 8500, 8750, 9000, 9250, 7500, 
    7750, 8000, 8250, 8500, 8750, 9000, 9250, 9500, 9750, 10000, 10250, 
    10500, 10750, 11000, 11250, 11500, 11750, 12000, 12250, 12500, 12750, 
    13000, 13250, 13500, 13750, 14000, 14250, 14500, 14750, 15000, 15250, 
    15500, 15750, 16000, 16250,
  500, 750, 1000, 1250, 1500, 1750, 2000, 2250, 2500, 2750, 3000, 3250, 3500, 
    3750, 4000, 4250, 4500, 4750, 5000, 5250, 5500, 5750, 6000, 6250, 6500, 
    6750, 7000, 7250, 7500, 7750, 8000, 8250, 8500, 8750, 9000, 9250, 7500, 
    7750, 8000, 8250, 8500, 8750, 9000, 9250, 9500, 9750, 10000, 10250, 
    10500, 10750, 11000, 11250, 11500, 11750, 12000, 12250, 12500, 12750, 
    13000, 13250, 13500, 13750, 14000, 14250, 14500, 14750, 15000, 15250, 
    15500, 15750, 16000, 16250,
  500, 750, 1000, 1250, 1500, 1750, 2000, 2250, 2500, 2750, 3000, 3250, 3500, 
    3750, 4000, 4250, 4500, 4750, 5000, 5250, 5500, 5750, 6000, 6250, 6500, 
    6750, 7000, 7250, 7500, 7750, 8000, 8250, 8500, 8750, 9000, 9250, 7500, 
    7750, 8000, 8250, 8500, 8750, 9000, 9250, 9500, 9750, 10000, 10250, 
    10500, 10750, 11000, 11250, 11500, 11750, 12000, 12250, 12500, 12750, 
    13000, 13250, 13500, 13750, 14000, 14250, 14500, 14750, 15000, 15250, 
    15500, 15750, 16000, 16250,
  500, 750, 1000, 1250, 1500, 1750, 2000, 2250, 2500, 2750, 3000, 3250, 3500, 
    3750, 4000, 4250, 4500, 4750, 5000, 5250, 5500, 5750, 6000, 6250, 6500, 
    6750, 7000, 7250, 7500, 7750, 8000, 8250, 8500, 8750, 9000, 9250, 7500, 
    7750, 8000, 8250, 8500, 8750, 9000, 9250, 9500, 9750, 10000, 10250, 
    10500, 10750, 11000, 11250, 11500, 11750, 12000, 12250, 12500, 12750, 
    13000, 13250, 13500, 13750, 14000, 14250, 14500, 14750, 15000, 15250, 
    15500, 15750, 16000, 16250,
  500, 750, 1000, 1250, 1500, 1750, 2000, 2250, 2500, 2750, 3000, 3250, 3500, 
    3750, 4000, 4250, 4500, 4750, 5000, 5250, 5500, 5750, 6000, 6250, 6500, 
    6750, 7000, 7250, 7500, 7750, 8000, 8250, 8500, 8750, 9000, 9250, 7500, 
    7750, 8000, 8250, 8500, 8750, 9000, 9250, 9500, 9750, 10000, 10250, 
    10500, 10750, 11000, 11250, 11500, 11750, 12000, 12250, 12500, 12750, 
    13000, 13250, 13500, 13750, 14000, 14250, 14500, 14750, 15000, 15250, 
    15500, 15750, 16000, 16250,
  500, 750, 1000, 1250, 1500, 1750, 2000, 2250, 2500, 2750, 3000, 3250, 3500, 
    3750, 4000, 4250, 4500, 4750, 5000, 5250, 5500, 5750, 6000, 6250, 6500, 
    6750, 7000, 7250, 7500, 7750, 8000, 8250, 8500, 8750, 9000, 9250, 7500, 
    7750, 8000, 8250, 8500, 8750, 9000, 9250, 9500, 9750, 10000, 10250, 
    10500, 10750, 11000, 11250, 11500, 11750, 12000, 12250, 12500, 12750, 
    13000, 13250, 13500, 13750, 14000, 14250, 14500, 14750, 15000, 15250, 
    15500, 15750, 16000, 16250,
  500, 750, 1000, 1250, 1500, 1750, 2000, 2250, 2500, 2750, 3000, 3250, 3500, 
    3750, 4000, 4250, 4500, 4750, 5000, 5250, 5500, 5750, 6000, 6250, 6500, 
    6750, 7000, 7250, 7500, 7750, 8000, 8250, 8500, 8750, 9000, 9250, 7500, 
    7750, 8000, 8250, 8500, 8750, 9000, 9250, 9500, 9750, 10000, 10250, 
    10500, 10750, 11000, 11250, 11500, 11750, 12000, 12250, 12500, 12750, 
    13000, 13250, 13500, 13750, 14000, 14250, 14500, 14750, 15000, 15250, 
    15500, 15750, 16000, 16250,
  500, 750, 1000, 1250, 1500, 1750, 2000, 2250, 2500, 2750, 3000, 3250, 3500, 
    3750, 4000, 4250, 4500, 4750, 5000, 5250, 5500, 5750, 6000, 6250, 6500, 
    6750, 7000, 7250, 7500, 7750, 8000, 8250, 8500, 8750, 9000, 9250, 7500, 
    7750, 8000, 8250, 8500, 8750, 9000, 9250, 9500, 9750, 10000, 10250, 
    10500, 10750, 11000, 11250, 11500, 11750, 12000, 12250, 12500, 12750, 
    13000, 13250, 13500, 13750, 14000, 14250, 14500, 14750, 15000, 15250, 
    15500, 15750, 16000, 16250,
  500, 750, 1000, 1250, 1500, 1750, 2000, 2250, 2500, 2750, 3000, 3250, 3500, 
    3750, 4000, 4250, 4500, 4750, 5000, 5250, 5500, 5750, 6000, 6250, 6500, 
    6750, 7000, 7250, 7500, 7750, 8000, 8250, 8500, 8750, 9000, 9250, 7500, 
    7750, 8000, 8250, 8500, 8750, 9000, 9250, 9500, 9750, 10000, 10250, 
    10500, 10750, 11000, 11250, 11500, 11750, 12000, 12250, 12500, 12750, 
    13000, 13250, 13500, 13750, 14000, 14250, 14500, 14750, 15000, 15250, 
    15500, 15750, 16000, 16250,
  500, 750, 1000, 1250, 1500, 1750, 2000, 2250, 2500, 2750, 3000, 3250, 3500, 
    3750, 4000, 4250, 4500, 4750, 5000, 5250, 5500, 5750, 6000, 6250, 6500, 
    6750, 7000, 7250, 7500, 7750, 8000, 8250, 8500, 8750, 9000, 9250, 7500, 
    7750, 8000, 8250, 8500, 8750, 9000, 9250, 9500, 9750, 10000, 10250, 
    10500, 10750, 11000, 11250, 11500, 11750, 12000, 12250, 12500, 12750, 
    13000, 13250, 13500, 13750, 14000, 14250, 14500, 14750, 15000, 15250, 
    15500, 15750, 16000, 16250 ;

 levelMode =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 2, 2, 2, 2, 2, 
    2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2 ;

 uComponent =
  4.499745, 9.899999, 10.52135, 11.86677, 12.28674, 10.03696, 8.485592, 
    6.768201, 7.094131, 9.800718, 11.51067, 12.22991, 11.38968, 10.30615, 
    9.420365, 9.03586, 7.418241, 6.311611, 6.333405, 6.499732, 6.634796, 
    7.58302, 8.272385, 9.05015, 11.19318, 12.87348, 14.65597, 15.95389, 
    14.09785, 13.98081, 13.74749, 13.46765, 13.53133, 13.82764, 14.42025, 
    14.95305, _, _, _, _, _, _, _, _, 15.73988, 16.78977, 18.52922, 20.39952, 
    22.22299, 23.43842, 24.63884, 25.70348, 26.37128, 27.13334, 27.82653, 
    29.11388, 30.20318, 30.4208, 29.05617, 28.66352, 26.39285, 23.50698, 
    20.77149, 17.7, 16.03873, 16.09755, 16.09755, 15.99756, _, _, 6.153786, _,
  3.95559, -2.688833, _, -2.6963, -2.899559, _, _, 0.6413809, 0.1622415, 
    26.60024, _, _, 0.9811226, 0.9969386, 0.09407578, 0.6363962, 4.30385, 
    8.98311, 9.228113, 3.731411, 8.74972, 8.376595, 9.335805, 8.739141, 
    8.798004, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  9.840886, 10.21463, 12.29756, 12.04228, 11.97953, 13.08326, 13.16359, 
    12.23516, 9.774936, 8.775657, 8.808247, 8.066499, 5.347216, 5.078737, 
    4.853488, 4.476803, 0.4808308, -0.4096326, 0.05584766, 0.4838436, 
    0.3882286, 0.3581249, 0.8965752, 1.213655, 1.485402, 1.649503, 1.538019, 
    1.782483, 2.282856, 2.765527, 3.312858, 4.189792, 5.791601, 6.913818, 
    8.197813, 8.912413, _, _, _, _, _, _, _, _, 9.90268, 10.242, 10.62024, 
    11.31503, _, _, _, 11.05307, 12.70459, _, _, _, _, _, _, _, 15.0908, 
    13.74749, 12.93872, 11.30133, 11.40013, _, _, _, _, _, _, _,
  0.1937216, -0.648967, -1.683995, -0.5704629, 1.194318, 4.305786, 5.558288, 
    4.408389, 3.85892, 4.131314, 3.538608, 1.741837, 3.051565, 4.51528, 
    5.053384, -18.13074, -2.35, _, -3.920849, _, _, _, _, _, _, -4.683896, _, 
    _, -2.617972, -3.599611, -2.4, -1.433472, -0.809824, -1.162869, 
    -2.275044, -2.427051, _, _, _, _, _, _, _, _, -2.621286, -2.810349, 
    -3.940233, _, _, -0.9587147, -0.5285941, -0.2966453, 0.3925199, 
    0.5752283, 0.2059064, 0.3087823, _, _, _, _, _, _, _, 1.367559, _, _, _, 
    _, _, _, _, _,
  9.515009, 16.98699, 19.9367, 20.46356, 18.95395, 14.63995, 12.5865, 
    11.17448, 10.49695, 9.577535, 9.125147, 8.431573, 8.488931, 8.69922, 
    7.828701, 7.549105, 7.733873, 7.8, 7.082253, 6.66324, 6.507784, 8.217229, 
    9.849999, 10.65, 11.91081, 12.22593, 14.25248, 14.24293, 13.12904, 
    12.94812, 12.58845, 12.73232, 13.16392, 13.82259, 14.71684, 15.32089, _, 
    _, _, _, _, _, _, _, 15.78052, 16.24014, 15.62249, 15.06589, 13.84456, 
    12.49793, 11.96673, 12.71806, 14.70525, 16.92821, 18.34671, 19.73358, 
    22.36954, 25.28277, 25.61035, 24.67501, 22.89518, 21.03444, 18.92766, 
    17.17066, 15.12981, 14.2387, 13.67912, 13.28609, 13.1193, 13.41336, 
    12.74416, _,
  7.658329, 15.22956, 20.98093, 20.05037, 17.71747, 15.54292, 12.53858, 
    10.95335, 9.495286, 9.169491, 8.397556, 7.32637, 6.759529, 6.524415, 
    6.078332, 6.683583, 7.3285, 7.454285, 8.456183, 8.120072, 8.416276, 
    9.063683, 9.616652, 9.256141, 10.28155, 11.20504, 12.85876, _, 14.25248, 
    16.32681, 17.92745, 16.4275, 15.0291, 14.93629, 13.9464, 12.69876, _, _, 
    _, _, _, _, _, _, 12.32456, 12.00532, 12.77409, 13.5193, 14.22261, 
    16.43892, 17.16084, 18.16855, 18.23234, _, 17.66615, 15.84459, 17.55866, 
    18.57401, 18.39767, 16.74545, 17.54033, 18.47791, _, _, _, _, _, _, _, _, 
    _, _,
  _, _, -2.831543, -1.427339, -0.3976119, -1.378955, -1.723191, -0.344944, 
    0.7873287, 2.253463, 3.386137, 3.95559, 2.832042, 1.299677, 0.2093439, 
    -0.89402, -0.4115632, 0.6013751, 1.507172, 2.3, 2.181644, 3.866937, 
    5.53802, 4.429327, 5.957969, 7.2635, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  11.85, 11.57529, 15.82773, 13.54084, 11.32817, 10.43457, 7.935099, 
    7.582428, 7.643051, 8.316857, 9.110669, 8.001781, 7.099999, 6.49645, 
    5.494038, 4.093205, 2.205725, 0.9277602, 0.6751342, 0.4257725, 1.377122, 
    2.676917, 4.757504, 8.619259, 9.702394, 10.21148, 10.67776, 11.03104, 
    11.41406, 12.21417, 13.01776, 13.21148, 13.13195, 12.87183, 12.87183, 
    13.2375, _, _, _, _, _, _, _, _, 13.52524, 13.88666, 13.97112, 14.19407, 
    14.24293, 14.18556, 13.69137, 12.93127, 12.2579, 11.78374, 13.47771, 
    15.19362, 16.55211, 17.87391, 18.7694, 19.58937, 20.22358, 19.70876, 
    17.66732, 15.83062, 14.82899, 14.33201, 14.51869, 14.08138, 13.4208, 
    12.83049, 11.32481, 8.952745,
  5.881324, 7.21845, 8.652637, 9.008628, 11.22149, 10.49645, 10.46257, 
    10.09685, 10.30013, 10.67776, 9.886696, 9.896313, 9.857423, 8.638307, 
    0.1186763, -4.738359, -6.490567, -4.082109, -3.223333, -3.169637, 
    -5.140217, -4.900001, -4.189387, -4.195595, -3.16983, -2.04905, 
    -1.924144, -1.720779, -1.097549, 0.1902311, 1.736422, 2.474462, 2.540179, 
    2.298257, 2.122316, 2.365228, _, _, _, _, _, _, _, _, 3.326743, 4.902685, 
    5.586143, 6.342584, 5.663085, _, _, _, _, 8.818283, 9.085973, 9.922162, 
    9.752552, 10.08654, 10.25833, 9.692532, 9.782644, 8.989309, 7.929957, 
    6.64711, 5.859952, 5.435139, 8.118625, 9.287254, 9.1, _, 3.275402, _,
  2.519033, 8.419446, 11.8172, 11.40754, 11.73973, 10.09268, 9.358398, 
    8.202438, 8.058038, 8.661378, 9.577535, 9.72745, 9.394442, 8.704142, 
    7.263849, 9.23458, 9.287005, 9.406652, 8.743668, 7.887121, 7.890679, 
    8.197539, 8.416725, 7.715331, 7.793227, 9.521368, 10.65213, 10.26702, 
    10.20966, 10.28915, 10.28624, 10.87402, 10.83564, 10.95018, 11.07604, 
    11.2019, _, _, _, _, _, _, _, _, 11.2666, 11.43449, 11.57937, 10.81035, 
    10.5, 9.579201, 8.832722, 9.299399, 9.739773, _, _, 35.74871, 16.86943, 
    18.50087, 21.00472, 16.92958, 17.56998, 17.15116, 16.35408, 16.48362, 
    16.40417, 15.00986, 13.25257, _, _, _, _, _,
  -1.273663, -1.023301, -2.490621, -4.82608, -8.437373, -10.64282, -12.59188, 
    -13.90745, -11.99299, -11.42616, -11.42405, -10.95444, -10.03518, 
    -8.09017, -7.609191, -8.100443, -7.975508, -7.65536, -8.296582, -7.51019, 
    -8.036908, -8.74972, -7.502649, -8.41207, -9.897017, -11.05451, 
    -9.866291, -10.67786, -9.960742, -9.774937, -9.355569, -10.06002, 
    -10.06837, -9.582943, -8.40024, -7.505054, _, _, _, _, _, _, _, _, 
    -7.656692, -7.012587, -8.296582, -10.69489, -11.30269, -12.14507, 
    -12.32326, -12.68585, -12.15066, -10.96632, -9.700776, -8.764789, 
    -8.688077, -9.287254, -10.4984, -11.79281, -12.36979, -10.7658, 
    -8.736482, -5.486602, -4.65426, -1.454429, 1.237231, 1.717645, 0.9742116, 
    0.9855365, _, _,
  10.81919, 13.28379, 14.03574, 12.90547, 12.90107, 12.71348, 10.77557, 
    9.033263, 8.266345, 4.585305, 5.398922, 7.100918, 4.840165, 1.26744, 
    9.179391e-07, -1.564344, -2.484664, -2.618555, -3.087138, -3.261121, 
    -3.338522, -2.804893, -1.350916, -0.8164424, 1.464218, 2.424733, 
    3.368171, 7.611512, 8.240607, 9.568859, 10.82498, 12.65721, 13.09123, 
    12.33332, 12.20119, 12.21417, _, _, _, _, _, _, _, _, 12.13536, 11.81262, 
    11.33746, 11.47159, 11.14977, 10.62816, 10.28155, 9.640111, 10.02136, 
    11.01267, 11.18474, 11.63121, 12.33189, 12.47, 11.9, 10.53176, 10.86311, 
    10.73455, 11.10757, 11.04507, 11.11658, 12.17177, 12.13372, 15.42901, 
    13.51331, _, 8.218971, _,
  9.899999, 14.52961, 16.26124, 15.73312, 14.4994, 15.13534, 15.41096, 
    14.99568, 14.84464, 15.1218, 14.11107, 9.61373, 7.070663, 6.232561, 
    6.556433, 4.789231, 0.3976115, -0.3768196, -1.910494, -4.431635, 
    -3.987755, -0.5119476, 2.755448, 3.355201, 4.476373, 6.949851, 7.534421, 
    8.269296, 9.849938, 10.67001, 11.18876, 11.44077, 11.49708, 11.51067, 
    11.69338, 12.15066, _, _, _, _, _, _, _, _, 12.70297, 13.33776, 13.59462, 
    13.75155, 13.3651, 13.90799, 13.25099, 12.61494, 14.49899, 14.74474, _, 
    _, 20.39609, 22.1078, 20.86118, 18.93686, 19.11624, 15.46148, 11.48504, 
    9.816273, 8.638307, 13.67516, 17.72654, 17.58085, 17.66732, 15.59762, 
    7.989036, _,
  9.676371, 9.80487, 10.56399, 9.7, 8.066218, 10.7756, 13.86541, 16.16292, 
    17.32276, 19.02775, 17.87391, 16.82934, 18.0103, 19.70116, 20.27223, 
    20.33783, 22.62741, 22.64234, 24.24358, 25.14664, 26.22992, 23.95224, 
    24.73229, _, _, _, _, _, 26.43146, _, 0.575929, _, _, _, 22, 21.95, _, _, 
    _, _, _, _, _, _, 23.33122, 22.73758, 22.01822, 22.9315, 24.25829, 
    25.21679, 25.2196, 24.71633, 24.66041, 22.30114, 22.73354, _, _, 
    26.58721, 19.50515, 18.33898, 16.66135, 14.22178, 13.75417, 13.66768, _, 
    5.209103, 5.051449, _, _, _, _, 5.542563,
  6.891078, 10.66878, 12.79075, 13.44921, 13.85929, 12.13926, 12.70242, 
    13.03251, 14.95408, 15.7289, 12.62615, 7.971755, 4.473544, 2.222025, 
    1.238641, -0.6975647, -1.419566, -1.328375, -1.544822, -1.850847, 
    -2.602109, -2.425609, -1.755443, -0.7324429, 1.072016, 1.072016, 
    0.6332654, 1.296153, 1.054585, 1.037154, 1.202077, 1.97959, 5.260453, 
    9.100025, 10.86144, 11.65752, _, _, _, _, _, _, _, _, 12.08606, 12.55737, 
    13.03183, 13.8997, 15.16485, 15.64858, 15.64858, 15.25621, 16.01678, 
    17.21985, _, 15.83062, 16.97191, 16.96096, 16.49785, 14.47824, 12.43439, 
    11.54664, 11.50905, 11.53133, 10.81873, 10.95444, 13.24641, 13.97226, 
    13.49844, 12.3461, 8.851245, 5.629823,
  13.33299, 11.60081, 23.24029, 24.90222, 25.3118, 23.81824, 24.94153, 
    24.22697, 21.82384, 18.10326, 16.55321, 14.86569, 12.22593, 10.76429, 
    10.1, 8.762017, 7.192448, 6.498383, 6.9165, 6.667998, 7.013937, 7.323756, 
    7.808638, 8.541467, 9.064961, 9.931529, 11.17342, 11.92759, 13.42063, 
    14.56392, 15.4269, 16.16336, 17.12029, 18.13757, 19.2346, 19.58686, _, _, 
    _, _, _, _, _, _, 19.64155, 19.73935, 20.52815, 21.41475, 22.5764, 
    23.47594, 24.81722, 26.53027, 27.19458, 28.87988, _, 28.6392, 27.27534, 
    25.5389, 24.31443, 22.86307, 21.62523, 20.14561, 17.87927, 13.30229, 
    14.25945, 14.55394, 17.91479, 19.03298, 17.85779, 14.60615, 12.02105, 
    10.70171,
  -0.2756374, 0.0453692, 0.3149315, 2.526692, 3.307387, 2.828652, 2.507952, 
    1.991716, 2.647452, 3.399482, 3.950753, 5.196832, 7.497842, 17.44872, 
    17.94813, 18.64071, -1.99847, -5.143004, -7.190352, 11.94983, 14.18936, 
    _, -0.6691306, -0.848048, -0.2930113, 0.7000002, -21.25326, 0.329932, 
    1.308986, 1.179536, 1.211266, 1.074374, 1.172045, 0.4509169, 0.6487511, 
    1.162869, _, _, _, _, _, _, _, _, 1.254288, 1.66762, 2.113092, -5.819074, 
    -25.69586, -25.61105, -26.28049, -26.71351, -24.43825, -26.19759, 
    -26.13095, _, -27.98783, _, _, _, -25.12626, -23.85838, _, _, -25.71606, 
    -25.79593, -26.21215, -27.19585, -27.19243, _, -29.09248, _,
  -0.4814908, -4.603728, -3.335398, -3.876626, -2.899559, -1.1, 0.1675171, 
    1.110684, 4.337115, 5.915341, 8.431573, 12.07149, 15.9099, 17.62383, 
    19.94009, 17.62097, 16.80756, 18.0615, 18.69082, 18.99711, 18.19723, _, 
    _, _, _, _, _, _, 22.11269, 23.73354, 22.87501, 22.23314, 23.48648, 
    23.07607, 19.57175, 20.75603, _, _, _, _, _, _, _, _, 22, 18.70441, 
    19.77053, 18.18112, 18.70988, _, 20.75056, 23.27087, 23.89936, 23.95235, 
    _, _, _, _, 20.14452, 16.78635, 15.68035, 15.25001, 13.89317, 11.01322, 
    5.253289, 4.796089, 7.167357, 5.643332, _, _, 4.682583, _,
  12.02013, 9.629041, 9.338523, 9.249999, 9.888729, 10.67492, 11.67521, 
    10.43909, 9.338523, 8.891168, 8.849652, 8.160756, 8.947087, 7.733873, 
    0.1902311, -5.817715, -7.523651, -7.141673, -4.607663, -5.328249, 
    -4.788283, -4.35714, _, -2.900297, -2.377804, -2.299586, _, _, -1.442493, 
    -1.18532, -0.6908358, -0.4292633, -0.2094295, 0.3873832, 2.565151, 
    4.266325, _, _, _, _, _, _, _, _, _, _, _, _, 4.557953, 5.431162, 
    4.377858, 2.588191, _, _, _, _, _, 12.73085, 2.04929, 3.597585, _, _, _, 
    _, 14.03575, _, _, _, _, _, _, _,
  7.853695, 14.28334, 13.71718, 12.16224, 13.33721, 15.0735, 15.03508, 
    9.800718, 7.628089, 7.883777, 9.770371, 10.30461, 10.16177, 9.479775, 
    7.018539, 6.481413, 6.538771, 6.524415, 7.193398, 8.143088, 9.522521, 
    10.58981, 11.50778, 12.22573, 12.22573, 13.10718, 14.13543, 15.0053, 
    14.39229, 15.06844, 15.18794, 15.16504, 14.97185, 14.97185, 15.10961, 
    15.31699, _, _, _, _, _, _, _, _, 15.68415, 15.76213, 15.69287, 15.49744, 
    15.48397, 15.81878, 17.57066, 18.4536, 20.49315, 22.73949, 24.14628, 
    28.22855, 29.63627, 29.59887, 30.10051, 25.05624, 21.08506, 18.43761, 
    16.35747, 14.65721, 13.89962, 15.88081, 15.88264, 14.7073, 13.39008, 
    12.22684, 9.03217, 5.192873,
  9.579706, 9.261407, 9.205792, 13.94201, 13.96213, 14.54923, 13.61183, 
    12.51557, 11.84013, 11.2844, 10.38216, 10.23246, 8.587327, 7.434268, 
    5.395049, 4.643503, 4.656971, 7.281151, 11.60203, 14.15995, 15.09974, 
    15.71647, 15.08848, 15.12981, 16.70583, 17.04054, 18.17264, _, 15.53774, 
    15.73312, 14, 13.9, 13.96252, 13.75552, 14.0372, 13.28264, _, _, _, _, _, 
    _, _, _, 12.8476, 11.83915, 11.20074, 11.08836, 12.44614, 11.2382, 
    12.46724, 12.98413, 13.33227, 15.74007, 16.81066, _, _, _, 23.42775, 
    22.69051, 20.56013, 20.04423, 18.81915, 17.31296, 13.37972, 11.50905, 
    11.0161, _, _, 12.41237, 8.723411, 8.144785,
  _, _, 1.102462, -0.9447947, -2.521009, -2.282139, -3.33524, -3.989177, 
    -3.408921, -4.741663, 0.584622, _, _, _, _, _, -0.2024559, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  _, -4.319062, 19.7283, 23.26381, _, 21.46179, 21.52585, 21.13837, 18.72725, 
    17.83963, 17.76116, 17.11368, 17.58473, 17.17066, 16.32007, 15.60261, 
    15.39608, 15.25001, 18.41836, 15.30878, 14.52656, 14.84648, 15.48564, 
    13.98483, 15.81142, 16.04884, 14.68356, 15.35843, 15.01872, 14.47824, 
    15.73312, 18.98179, 15.53172, 22.14679, 24.95857, 15.42142, _, _, _, _, 
    _, _, _, _, 16.39394, 18.20705, 18.05842, 23.32015, 28.09546, 34.0348, 
    35.67108, 37.51137, _, _, 34.57105, 35.33244, 34.38696, 30.98497, 
    29.63787, 28.26398, 25.9762, 25.846, 19.06238, 15.97926, 16.2443, 
    16.26292, 15.28406, 13.44631, 10.39781, _, _, _,
  -1.5802, -0.2233565, 2.210179, 5.374011, 6.685904, 8.376595, 8.075423, 
    6.898949, 6.064515, 5.657513, 7.48173, 2.155704, 1.792298, 9.447958, 
    8.398721, 5.369358, 4.916696, 4.682115, 5.715768, 5.248473, 5.811265, 
    6.171605, 5.870843, 6.868265, 8.146081, 8.82572, 9.202318, 7.863861, 
    8.04758, 9.475232, 10.62697, 12.45886, 14.17353, 15.32865, 16.776, 
    13.73653, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, 10.67731, _, _, _, _, _, _, _, _, -40.60259,
  0.1394493, -1.427339, -3.603451, -4.925292, -4.782836, -5.034564, 
    -4.641302, -2.595743, -4.312911, -14.42068, -15.34119, -11.3043, 
    -5.965195, -4.878617, -4.680664, -4.476373, -5.216, -5.558259, -3.168858, 
    -5.190813, _, _, _, _, _, _, _, _, _, _, -38.88581, -11.87609, -10.32306, 
    -11.06257, -12.00981, -11.89275, _, _, _, _, _, _, _, _, -10.53744, 
    -11.91055, -12.4964, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _,
  4.506927, 6.490567, 7.696936, 8.266435, 7.872709, 7.347862, 7.347862, 
    7.212488, 6.867857, 7.354028, 7.945776, 8.660254, 9.866773, 10.93715, 
    11.18876, 11.87451, 12.49324, 12.66393, 12.07535, 10.7509, 12.43301, 
    11.3924, 11.64287, 11.6008, 13.45092, 14.30996, 15.98061, _, 15.12235, 
    14.89901, 15.25713, 15.15569, 14.011, 13.70857, 13.66162, 13.61467, _, _, 
    _, _, _, _, _, _, 14.15644, 14.25, 15.849, 17.05539, 17.39844, _, _, _, 
    _, _, _, _, _, _, _, _, 26.12346, 26.79561, 27.06284, 25.28599, 24.66573, 
    23.19672, _, _, _, _, 11.56727, 9.448977 ;

 uComponentDD =
  "SSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSZZZZZZZZSSSSSSSSSSSSSSSSSSSSSSSSZZSZ",
  "SQZSSZZSSQZZSSSSSSSSSSSSSZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ",
  "SSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSZZZZZZZZSSSSZZZSSZZZZZZZSSSSSZZZZZZZ",
  "SSSSSSSSSSSSSSSQSZSZZZZZZSZZSSSSSSSSZZZZZZZZSSSZZSSSSSSSZZZZZZZQZZZZZZZZ",
  "QQQSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSZZZZZZZZSSSSSSSSSSSSSSSSSSSSSSSSSSSZ",
  "QQSSSSSSSSSSSSSSSSSSSSSSSSSZSSSSSSSSZZZZZZZZSSSSSSSSSZSSSSSSSSZZZZZZZZZZ",
  "ZZSSSSSSSSSSSSSSSSSSSSSSSSZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ",
  "QQSSQQSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSZZZZZZZZSSSSSSSSSSSSSSSSSSSSSSSSSSSS",
  "SSSSQSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSZZZZZZZZSSSSSZZZZSSSSSSSSSSSSSSSSZSZ",
  "SSSQQSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSZZZZZZZZSSSSSSSSSZZQSSSSSSSSSSSZZZZZ",
  "SSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSZZZZZZZZSSSSSSSSSSSSSSSSSSSSSSSSSSZZ",
  "SSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSZZZZZZZZSSSSSSSSSSSSSSSSSSSSSSSSSZSZ",
  "SSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSZZZZZZZZSSSSSSSSSSZZSSSSSSSSSSSSSSSZ",
  "SSSSSSSSSSSSSSSSSSSSSSSZZZZZSZQZZZSSZZZZZZZZSSSSSSSSSSSZZSSSSSSSZSSZZZZQ",
  "SQSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSZZZZZZZZSSSSSSSSSSZSSSSSSSSSSSSSSSSS",
  "QQQQSQSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSZZZZZZZZSSSSSSSSSSZSSSSSSSSSSSSSSSSS",
  "SSSSSSQQQQSQQSQQSSQQQZSSSSQSSSSSSSSSZZZZZZZZSSSSQQQQQQQZQZZZQQZZQQQQQZQZ",
  "SSSSSSSSSSQQSSSSSSSQQZZZZZZZQSSSSSSSZZZZZZZZSSSSSZSSSSZZZZSSSSSSSSSSZZSZ",
  "SSSSSSSSSSSSSSSSSSSSSSZSSSZZSSSSSSSSZZZZZZZZZZZZSSSSZZZZZQSSZZZZQZZZZZZZ",
  "QSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSZZZZZZZZSSSSSSSSSSSSSSSSSSSSSSSSSSSS",
  "QSSSSSSSSSSSSSSSSSSSSSSSSSSZSSSSSSSSZZZZZZZZSSSSSSSSSSSZZZSSSSSSSSSZZSSS",
  "ZZSSSSSSSSSZZZZZQZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ",
  "ZQQQZSQQSSSSSSSSSSSSSSSSSSSSSSSSSQQSZZZZZZZZSSSSSSSSZZSSSSSSSSSSSSSSSZZZ",
  "SSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSZZZZZZZZZZZZZZZZZZZZZZZZZZQZZZZZZZZQ",
  "QQQSSSSQQQQSSSSSSSSSZZZZZZZZZZQSSSSSZZZZZZZZSSSZZZZZZZZZZZZZZZZZZZZZZZZZ",
  "SSSSSSSSSSSSSSSSSSSSSSSSSSSZSSSSSSSSZZZZZZZZSSSSSZZZZZZZZZZZSSSSSSZZZZQQ" ;

 uComponentQCA =
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 523, 523, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 0, 515, 0,
  523, 523, 0, 523, 523, 0, 0, 523, 523, 523, 0, 0, 523, 523, 523, 523, 523, 
    515, 515, 515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 523, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 
    515, 0, 0, 0, 515, 515, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 515, 515, 0, 
    0, 0, 0, 0, 0, 0,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 523, 0, 515, 0, 0, 0, 0, 0, 0, 515, 0, 0, 515, 515, 515, 515, 515, 
    515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 0, 0, 515, 515, 
    515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 515, 0, 0, 0, 0, 0, 0, 0, 0,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 523, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 0,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 0, 515, 515, 
    515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 0, 515, 515, 515, 515, 515, 515, 515, 515, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 523, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 523, 523, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 
    515, 515, 0, 0, 0, 0, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 0, 515, 0,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 0, 0, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 0, 0, 0, 0, 0,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 523, 523, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 515, 0, 0,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 523, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 0, 515, 0,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 523, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 0, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 515, 0,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 515, 0, 515, 0, 0, 
    0, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 0, 0, 515, 515, 515, 515, 515, 515, 515, 0, 515, 515, 
    0, 0, 0, 0, 515,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 523, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 515, 515,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 515, 515,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 523, 523, 515, 515, 515, 0, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 515, 0, 0, 0, 515, 515, 0, 0, 515, 
    515, 515, 515, 515, 0, 515, 0,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 515, 
    515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 515, 515, 0, 
    515, 515, 515, 515, 0, 0, 0, 0, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 0, 0, 515, 0,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 523, 515, 515, 515, 515, 515, 0, 515, 515, 515, 0, 0, 515, 515, 515, 
    515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 
    515, 515, 0, 0, 0, 0, 0, 515, 515, 515, 0, 0, 0, 0, 515, 0, 0, 0, 0, 0, 
    0, 0,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 523, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 0, 515, 515, 
    515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 0, 0, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 0, 0, 515, 515, 515,
  0, 0, 523, 523, 523, 523, 523, 523, 523, 523, 523, 0, 0, 0, 0, 0, 523, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 523, 523, 523, 0, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 515, 
    515, 515, 515, 515, 0, 0, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 0, 0, 0,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 523, 523, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 523, 523, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 
    515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 0, 515, 515, 
    515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 515, 
    515, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 515, 515, 515, 0, 0, 
    0, 0, 515, 515 ;

 uComponentQCR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 9, 0, 0, 0, 0, 0, 0, 0, 513, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 513, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 513, 0, 0, 0, 0, 0, 0, 0, 0,
  9, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  9, 9, 0, 0, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 513, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 513, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 513,
  0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  9, 9, 9, 9, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 9, 9, 9, 9, 0, 9, 9, 0, 513, 513, 0, 0, 513, 513, 513, 0, 
    0, 0, 0, 0, 513, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 513, 513, 513, 513, 513, 513, 513, 0, 513, 0, 0, 0, 513, 513, 0, 0, 
    513, 513, 513, 513, 513, 0, 513, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 0, 0, 0, 0, 0, 0, 0, 513, 513, 0, 0, 0, 
    0, 0, 0, 0, 513, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 513, 0, 0, 0, 0, 0, 0, 513, 0, 0, 0, 0, 0, 0, 0,
  9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 513, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 513, 9, 9, 0, 0, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 513, 513, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 513, 0, 0, 0, 0, 0, 0, 0, 0, 513,
  9, 9, 9, 0, 0, 0, 0, 9, 9, 513, 513, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 513, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 513, 513 ;

 uComponentICA =
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 0, 3, 3, 0, 0, 3, 3, 3, 0, 0, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 3, 3, 3, 0, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 uComponentICR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 0, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 3, 3, 3, 3, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 3, 3, 0, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 0, 0, 0, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 vComponent =
  18.0475, 17.1473, 14.48141, 12.72556, 11.45757, 11.14717, 11.26076, 
    9.665995, 6.615384, 5.211135, 5.124882, 4.694618, 4.372087, 3.548693, 
    2.701245, 2.59099, 2.410333, 1.929654, 1.462183, 1.146078, 0.9324608, 
    1.337091, 1.458644, 0.9512079, -0.3908723, -1.809253, -2.059764, -2.8131, 
    0.2460774, 0.7327057, 1.202749, 1.892756, 2.143153, 2.190083, 2.283944, 
    2.101516, _, _, _, _, _, _, _, _, 1.37706, 0.586316, -1.621097, 
    -2.866969, -3.519777, -4.132826, -4.789303, -4.532217, -4.176802, 
    -3.813348, -3.910769, -4.091694, -4.244785, -4.818183, -5.647943, 
    -5.57162, -4.65377, -3.723142, -1.088592, -2.110704e-07, 1.403207, 
    0.280982, -0.2809823, 0.2792367, _, _, 0.7555915, _,
  4.241852, 1.086359, _, -0.1413071, -0.05061191, _, _, 4.049522, 3.095751, 
    -3.266093, _, _, -0.8528765, -0.46488, -0.8950697, -0.636396, -0.9148105, 
    -2.407017, -2.646117, -2.331646, -2.842957, -3.555655, -3.583678, 
    -3.180787, -2.689818, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _,
  11.32064, 9.864148, 7.099998, 7.524855, 9.027227, 8.49637, 7.599998, 
    5.705346, 4.352082, 3.368657, 3.558764, 3.259079, 2.493447, 2.587747, 
    2.367203, 3.019642, 4.5748, 4.682115, 3.199513, 1.940591, 1.448889, 
    1.040071, -0.07844016, -0.4658781, -0.2087599, -0.4112673, -0.4410195, 
    0.2505119, 0.2803001, 0.4380167, 0.764834, 0.9672901, 1.125772, 1.095042, 
    1.298407, 1.252559, _, _, _, _, _, _, _, _, 1.391733, 1.805941, 1.304005, 
    1.389313, _, _, _, 2.349405, 1.559931, _, _, _, _, _, _, _, -0.5269796, 
    1.202749, 2.049292, 3.028182, 2.631929, _, _, _, _, _, _, _,
  11.09831, 12.38301, 11.98224, 10.88506, 9.726953, 6.383589, 5.183187, 
    6.067628, 7.573555, 8.10816, 7.947845, 6.986129, 5.73916, 4.675709, 
    4.550089, -1.586236, 4.070319, _, 1.198724, _, _, _, _, _, _, 7.212567, 
    _, _, 4.722947, 4.289849, 4.156922, 3.734322, 3.507732, 3.194955, 
    2.526692, 1.763355, _, _, _, _, _, _, _, _, 1.835445, 3.121208, 5.043269, 
    _, _, 10.95814, 10.08616, 8.494823, 7.489721, 6.574885, 5.896406, 
    5.891914, _, _, _, _, _, _, _, 3.221767, _, _, _, _, _, _, _, _,
  23.55047, 23.38059, 20.64505, 13.28919, 12.30884, 13.18188, 12.5865, 
    12.41052, 12.07535, 11.41406, 11.26862, 12.04154, 12.12345, 11.97345, 
    11.60653, 11.19201, 11.90912, 13.51, 13.8997, 13.66167, 14.61673, 
    16.12722, 17.0607, 18.44634, 17.6585, 16.82755, 15.82898, 13.75423, 
    13.59552, 12.50385, 12.15652, 12.29545, 12.71225, 12.88977, 12.79315, 
    12.85575, _, _, _, _, _, _, _, _, 13.24142, 13.6271, 13.58042, 14.04917, 
    14.84648, 15.99662, 17.7414, 20.35315, 22.64411, 23.29969, 23.48272, 
    23.51757, 23.9884, 21.97798, 20.009, 17.92746, 16.63433, 15.28242, 
    14.26302, 12.93903, 11.8207, 10.34502, 9.226683, 7.983094, 7.272144, 
    6.254749, 4.140829, _,
  18.04189, 18.80693, 18.23844, 16.23646, 12.8725, 12.58641, 9.448498, 
    8.557694, 9.16949, 9.495285, 9.660282, 9.377329, 9.303697, 8.98009, 
    8.066218, 7.167267, 5.725652, 5.219545, 5.703767, 6.813548, 8.127502, 
    8.752695, 9.616653, 11.03104, 13.15978, 14.3418, 14.79231, _, 15.82898, 
    19.45753, 24.67502, 26.28949, 27.11321, 29.31412, 29.90816, 29.91641, _, 
    _, _, _, _, _, _, _, 30.50435, 31.27495, 31.61697, 31.84947, 33.50638, 
    33.70478, 33.68005, 34.17007, 30.34373, _, 25.22988, 25.35664, 26.03178, 
    25.56494, 25.32223, 26.79832, 28.07039, 19.13444, _, _, _, _, _, _, _, _, 
    _, _,
  _, _, 6.072262, 5.724745, 5.686115, 5.530685, 4.265046, 3.281922, 3.410295, 
    4.238149, 4.33406, 4.241852, 3.62485, 3.570832, 3.994518, 4.206035, 
    5.885628, 6.873744, 6.528279, 3.983717, 3.935788, 5.954561, 6.838884, 
    7.37164, 7.906491, 8.656303, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  20.5248, 17.16108, 21.00411, 17.9693, 14.4994, 11.18971, 10.92173, 
    10.43632, 10.14267, 11.8777, 12.53976, 12.80553, 12.29756, 11.7199, 
    11.782, 13.38827, 13.92641, 13.2676, 12.88232, 12.19257, 11.21577, 
    11.595, 11.77523, 11.03215, 10.7756, 10.5743, 9.957176, 9.25614, 
    9.577534, 9.542753, 9.809587, 10.69845, 11.41543, 12.00317, 12.00317, 
    12.34417, _, _, _, _, _, _, _, _, 12.17818, 12.07149, 12.57966, 12.7804, 
    13.75423, 15.21216, 16.31675, 17.79838, 20.40058, 22.16199, 24.31443, 
    25.28644, 24.53951, 23.71947, 22.3685, 20.28538, 16.96959, 12.79902, 
    9.793155, 8.775054, 8.910162, 8.955637, 8.04784, 7.805435, 7.135969, 
    6.537466, 5.523474, 3.986019,
  14.55679, 14.167, 14.40041, 14.41682, 10.10387, 14.99048, 14.4005, 
    12.92338, 11.84894, 9.957176, 8.594374, 6.426742, 5.922941, 5.609783, 
    6.798965, 7.296433, 7.208505, 6.051974, 6.326146, 6.797308, 8.226066, 
    8.487049, 9.409518, 10.38446, 11.05451, 11.62073, 12.14857, 10.86457, 
    10.44248, 10.89834, 10.96334, 10.71807, 10.18811, 9.21781, 7.920591, 
    6.161631, _, _, _, _, _, _, _, _, 4.751082, 4.11384, 5.586144, 6.80159, 
    12.14452, _, _, _, _, 6.406861, 5.459406, 6.200057, 6.094073, 7.880467, 
    8.307028, 7.572637, 6.598476, 5.617146, 4.040517, 3.684553, 3.248224, 
    2.769343, 1.725669, 0.486726, -1.085164e-07, _, -0.4021682, _,
  17.92385, 18.91039, 18.91147, 16.91236, 12.15684, 9.411577, 8.135132, 
    8.202439, 8.344342, 9.288193, 11.41406, 12.45057, 13.92783, 14.48613, 
    14.2561, 13.18835, 12.78247, 13.43409, 13.99279, 14.83352, 16.17829, 
    16.80745, 17.25685, 15.81878, 14.65693, 13.59792, 14.13585, 14.66282, 
    14.58091, 15.25429, 14.1578, 14.96682, 13.86899, 13.52234, 13.67777, 
    13.8332, _, _, _, _, _, _, _, _, 14.4206, 15.17407, 15.93764, 17.30018, 
    18.18653, 18.80024, 18.94183, 21.90801, 24.10678, _, _, 28.94873, 
    23.21879, 21.28281, 20.28402, 14.2056, 13.23993, 12.46105, 10.62046, 
    8.398828, 7.649389, 7.320796, 11.12022, _, _, _, _, _,
  3.152425, 3.347067, 3.985826, 4.049562, 3.40892, 4.085394, 4.583069, 
    5.061898, 7.788339, 8.927091, 9.251009, 9.191863, 8.420518, 5.877852, 
    4.217843, 3.438434, 3.719041, 2.938617, 1.314049, 3.034314, 2.767329, 
    2.842956, 1.732123, 1.78804, 2.467603, 3.16983, 4.392755, 4.532482, 
    3.625413, 4.352081, 4.766899, 4.691063, 5.130092, 5.988089, 5.047373, 
    3.990508, _, _, _, _, _, _, _, _, 1.48831, 1.110685, 1.314049, 1.503069, 
    2.609432, 3.713121, 4.730457, 4.617272, 5.157651, 5.113682, 3.151973, 
    1.545469, 0.4553227, 0.4867243, 0.1832497, 0.4118136, 0.8649803, 
    1.705135, 1.6982, 0.3836606, -0.6541136, -2.623859, -5.359035, -6.8891, 
    -6.931876, -6.222437, _, _,
  24.30031, 23.96458, 20.80884, 18.43092, 15.93149, 14.11975, 11.55539, 
    10.03245, 9.50934, 8.999166, 10.1539, 11.36384, 10.87119, 10.32248, 10.5, 
    9.876884, 9.272888, 9.131986, 10.76613, 12.17067, 13.39008, 14.42992, 
    15.44102, 15.57862, 16.73607, 15.30917, 15.84599, 13.73153, 13.71468, 
    12.6983, 12.45271, 12.65721, 12.20777, 10.34888, 9.880329, 9.542753, _, 
    _, _, _, _, _, _, _, 9.481187, 9.565669, 9.513255, 9.972097, 10.7672, 
    12.2263, 13.15978, 14.84447, 15.43154, 15.72772, 15.97346, 17.24398, 
    17.61177, 18.48754, 20.6114, 13.97612, 12.94615, 12.79294, 12.3362, 
    11.4375, 10.36637, 7.313544, 5.918008, 9.27069, 9.114843, _, 5.337463, _,
  17.1473, 18.59706, 11.81449, 11.85576, 11.32817, 7.057724, 5.609129, 
    4.299941, 5.11142, 4.913372, 6.882424, 7.51107, 8.42649, 7.169741, 
    7.813654, 5.50938, 5.686115, 7.190132, 4.728637, -0.781417, -1.85952, 
    0.4773988, 3.16978, 1.783992, 1.99301, 3.541127, 4.349999, 3.009777, 
    3.011431, 3.059573, 3.420751, 3.939375, 4.645124, 5.124882, 5.206229, 
    5.157652, _, _, _, _, _, _, _, _, 5.392091, 5.938355, 6.339272, 6.707076, 
    6.80986, 8.690678, 8.605298, 8.833076, 10.1523, 10.32437, _, _, 10.8448, 
    9.843027, 7.592846, 5.430053, 6.211244, 2.726276, 2.232464, 1.908088, 
    5.609783, 4.180918, 3.125666, 2.784534, 2.169279, 0.2722558, 0.418689, _,
  -0.6766387, -2.8115, -2.245444, -1.156713e-07, 6.078333, 9.702394, 
    11.63445, 15.07216, 18.57639, 20.40477, 23.71947, 25.91492, 25.72137, 
    25.21635, 23.32052, 23.396, 22.62742, 24.28094, 25.10496, 26.0401, 
    29.13128, 31.78569, 30.54183, _, _, _, _, _, 32.64013, _, 32.99498, _, _, 
    _, 38.10512, 38.01852, _, _, _, _, _, _, _, _, 38.82968, 41.01966, 
    41.41024, 41.36951, 40.37258, 38.83045, 37.38959, 36.64346, 36.56055, 
    37.11535, 36.38126, _, _, 26.58722, 20.91672, 18.99057, 18.5043, 
    18.20305, 18.931, 17.49384, _, 4.370955, 4.090582, _, _, _, _, 3.2,
  21.20856, 20.93865, 18.26709, 15.47155, 13.85929, 9.147591, 5.132113, 
    6.356379, 6.9732, 7.671492, 6.713444, 7.433782, 6.6323, 7.267916, 
    8.813385, 9.975641, 10.10073, 10.81875, 10.99198, 9.521783, 8.511111, 
    8.459103, 9.03097, 10.47442, 12.25319, 12.25319, 12.08342, 12.33207, 
    12.05396, 11.85472, 11.437, 11.22681, 10.78553, 9.423351, 8.184687, 
    7.570483, _, _, _, _, _, _, _, _, 7.262041, 7.249999, 7.223663, 7.082254, 
    6.751828, 6.642431, 6.642431, 6.792502, 6.798723, 8.029745, _, 8.775054, 
    10.19776, 10.59839, 11.12794, 12.14868, 12.87618, 13.28289, 12.78209, 
    11.94104, 10.81873, 9.191861, 5.897681, 3.483676, 2.869184, 1.955431, 
    0.9303021, 0.8916767,
  25.07571, 17.86368, 17.51282, 17.43672, 17.72351, 15.46775, 14.4, 13.42923, 
    12.6, 12.67604, 13.40452, 15.39387, 16.82755, 17.9148, 17.49371, 
    17.19642, 17.80193, 17.85416, 18.0181, 16.50387, 14.38071, 13.77398, 
    15.32531, 19.18446, 21.35571, 21.29823, 21.01415, 18.36689, 19.8969, 
    19.32698, 18.38507, 17.33308, 16.53287, 16.91356, 17.93656, 19.58686, _, 
    _, _, _, _, _, _, _, 21.06299, 21.92277, 22.01375, 22.96451, 23.37854, 
    23.47595, 23.96571, 23.88797, 22.81896, 24.23309, _, 20.80761, 18.39745, 
    14.15644, 13.47771, 13.2, 13.51294, 13.58839, 12.99006, 11.97744, 
    9.618118, 13.57177, 10.7643, 5.457616, 7.580185, 8.096321, 8.108297, 
    8.064323,
  0.9612617, 1.299208, 1.364118, 2.275044, 2.066686, 1.699626, 1.822135, 
    1.671247, 0.9115909, 0.05933781, -0.6257381, 0.1814788, 2.14997, 7.76867, 
    6.532583, 6.056735, -2.750658, -3.090229, -3.506969, 4.587108, 5.164503, 
    _, 0.7431448, 0.5299193, -0.8509667, -1.212435, -11.78087, -1.871135, 
    -2.361474, -2.649282, -2.853565, -3.120211, -3.403867, -3.672421, 
    -3.337533, -3.194955, _, _, _, _, _, _, _, _, -3.267531, -3.745537, 
    -4.531538, -8.009268, -16.05655, -16.00356, -17.72642, -16.69246, 
    -18.41554, -17.6705, -18.29709, _, -15.51391, _, _, _, -21.08343, 
    -19.32014, _, _, -19.37844, -19.43863, -19.04424, -19.04274, -18.34153, 
    _, -13.56604, _,
  -9.187391, -4.00196, -4.118874, -1.334829, 0.05061182, 1.905256, 4.797076, 
    7.012587, 10.2176, 11.12514, 12.04154, 13.88665, 15.9099, 17.01913, 
    22.14572, 21.76009, 21.5127, 22.30409, 23.08123, 0.3315936, -0.3176322, 
    _, _, _, _, _, _, _, 95.78058, 25.45111, 22.09014, 23.84213, 26.08438, 
    27.501, 29.01631, 34.54384, _, _, _, _, _, _, _, _, 38.10512, 36.70947, 
    40.53561, 40.83548, 42.02309, _, 44.49971, 41.98174, 38.24697, 38.33178, 
    _, _, _, _, 14.63586, 13.59332, 14.11866, 14.72676, 14.3868, 14.61503, 
    16.16796, 16.72595, 18.67161, 15.50493, _, _, 11.5898, _,
  14.32503, 12.77817, 13.84493, 16.02147, 16.45761, 16.43794, 15.49353, 
    14.90857, 13.84493, 13.1817, 14.1624, 13.05994, 13.2646, 11.90912, 
    10.89834, 10.49544, 10.35542, 9.140925, 11.40436, 11.96745, 13.1557, 
    13.4099, _, 14.92073, 15.01286, 14.51902, _, _, 13.7244, 13.54825, 
    13.18191, 12.29251, 11.99817, 11.09324, 7.047695, 7.696653, _, _, _, _, 
    _, _, _, _, _, _, _, _, 13.23726, 12.79502, 12.02807, 9.659258, _, _, _, 
    _, _, -28.59398, 12.93872, 13.42637, _, _, _, _, -20.80884, _, _, _, _, 
    _, _, _,
  18.50215, 18.28185, 15.23447, 12.16224, 10.05031, 6.711154, 5.472321, 
    5.211135, 8.47185, 10.46212, 11.64388, 11.44443, 10.89717, 10.16582, 
    8.983323, 9.256418, 9.338333, 8.98009, 6.946583, 4.892864, 3.655351, 
    3.646363, 3.739107, 3.048216, 3.048216, 2.78602, 2.747647, 3.464248, 
    3.856403, 4.037576, 4.355068, 4.063458, 4.011694, 4.011694, 4.619476, 
    5.574927, _, _, _, _, _, _, _, _, 6.020578, 6.368315, 5.711735, 5.948905, 
    6.255934, 7.715329, 9.342485, 9.811957, 10.44179, 11.09079, 12.30315, 
    12.56816, 13.81961, 13.17827, 12.77691, 8.627557, 7.26017, 6.348579, 
    5.632329, 5.626374, 5.900042, 5.780139, 5.160586, 4.217249, 3.338523, 
    2.598899, 1.109013, 0.2721478,
  15.94331, 18.17653, 18.87468, 11.69873, 12.13709, 8.399998, 6.060376, 
    5.572292, 4.309453, 3.449988, 2.588565, 3.128379, 3.823324, 4.120882, 
    5.209938, 6.391235, 5.75088, 5.290069, 5.165555, 6.304418, 7.364632, 
    8.356595, 10.17731, 11.8207, 13.05202, 15.89056, 18.17265, _, 15.00462, 
    11.85576, 24.24871, 24.0755, 25.18904, 25.87037, 26.40013, 27.23346, _, 
    _, _, _, _, _, _, _, 27.55176, 27.8913, 27.7228, 27.44464, 27.95449, 
    27.81551, 26.73608, 25.48279, 24.05204, 24.23758, 23.13789, _, _, _, 
    16.40428, 15.88806, 13.86798, 13.01687, 12.69368, 12.57861, 12.92065, 
    12.78209, 16.33204, _, _, 13.31064, 12.93299, 11.63196,
  _, _, 0.6888952, 4.092354, 4.548023, 4.894062, 7.491073, 8.179027, 
    8.437373, 8.91777, -0.1349707, _, _, _, _, _, -0.876933, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _,
  _, 18.70791, 20.42925, 23.26381, _, 15.0277, 18.06233, 17.11751, 16.86209, 
    17.22753, 15.99222, 15.95876, 15.28617, 12.93903, 13.21573, 12.1901, 
    13.3836, 14.72676, 14.91489, 13.78409, 15.57783, 13.84457, 15.48564, 
    15.53173, 21.76256, 23.79338, 20.97029, 14.32197, 13.05557, 12.14868, 
    11.85576, 6.908805, 13.98483, -29.38979, -27.7193, 15.96934, _, _, _, _, 
    _, _, _, _, 16.97642, 16.3937, 16.25987, 17.573, 18.24541, 19.65, 
    18.96665, 19.11301, _, _, 17.61484, 12.85995, 9.213956, 7.153447, 
    6.299731, 4.983702, 4.114228, 3.632422, 3.019186, 5.502102, 6.235599, 
    5.599773, 4.382631, 3.104326, 1.461319, _, _, _,
  8.961751, 6.396101, 5.470385, 5.374012, 4.017299, 3.555654, 1.423915, 
    0.1204208, -1.289051, -0.694654, 0.5231741, -4.841792, -5.516128, 
    0.9930192, 0.1465993, -3.099999, -1.692955, -0.4096319, -3.299999, 
    -6.037676, -5.051653, -3.708273, -5.286133, -5.175611, -6.138515, 
    -6.895409, -6.207041, -5.506333, -8.629975, -9.475229, -9.56857, 
    -9.051889, -9.204401, -8.849998, -8.919962, -10.35122, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, -10.67731, _, 
    _, _, _, _, _, _, _, -18.9333,
  1.593912, 5.724745, 5.766727, 6.304086, 5.906309, 6.217167, 6.881011, 
    7.988874, 8.464561, 3.329275, 21.11535, 7.915355, 8.519181, 6.714842, 
    4.364789, 1.993009, 1.397623, 0.682468, -0.445354, -1.488442, _, _, _, _, 
    _, _, _, _, _, _, -4.087061, 5.287576, 4.596124, 3.809147, 1.474618, 
    0.4153036, _, _, _, _, _, _, _, _, 1.858036, 1.462431, 3.583286, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  8.476297, 7.208505, 7.432844, 8.560143, 9.056515, 8.452746, 8.452746, 
    7.21249, 5.970138, 6.170761, 5.56369, 4.999999, 3.591211, 3.553697, 
    3.420751, 5.040432, 6.093356, 8.224051, 10.49694, 10.02538, 11.59397, 
    11.79717, 12.93072, 12.01297, 12.11127, 14.8184, 15.98061, _, 16.79507, 
    19.06986, 21.78945, 24.25418, 25.27651, 25.78207, 25.69378, 25.60548, _, 
    _, _, _, _, _, _, _, 25.53889, 24.68172, 24.40532, 25.28564, 23.94691, _, 
    _, _, _, _, _, _, _, _, _, _, 9.508158, 10.82614, 11.4875, 11.79105, 
    10.98189, 9.846427, _, _, _, _, 9.706092, 11.26085 ;

 vComponentDD =
  "SSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSZZZZZZZZSSSSSSSSSSSSSSSSSSSSSSSSZZSZ",
  "SQZSSZZSSQZZSSSSSSSSSSSSSZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ",
  "SSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSZZZZZZZZSSSSZZZSSZZZZZZZSSSSSZZZZZZZ",
  "SSSSSSSSSSSSSSSQSZSZZZZZZSZZSSSSSSSSZZZZZZZZSSSZZSSSSSSSZZZZZZZQZZZZZZZZ",
  "QQQSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSZZZZZZZZSSSSSSSSSSSSSSSSSSSSSSSSSSSZ",
  "QQSSSSSSSSSSSSSSSSSSSSSSSSSZSSSSSSSSZZZZZZZZSSSSSSSSSZSSSSSSSSZZZZZZZZZZ",
  "ZZSSSSSSSSSSSSSSSSSSSSSSSSZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ",
  "QQSSQQSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSZZZZZZZZSSSSSSSSSSSSSSSSSSSSSSSSSSSS",
  "SSSSQSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSZZZZZZZZSSSSSZZZZSSSSSSSSSSSSSSSSZSZ",
  "SSSQQSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSZZZZZZZZSSSSSSSSSZZQSSSSSSSSSSSZZZZZ",
  "SSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSZZZZZZZZSSSSSSSSSSSSSSSSSSSSSSSSSSZZ",
  "SSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSZZZZZZZZSSSSSSSSSSSSSSSSSSSSSSSSSZSZ",
  "SSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSZZZZZZZZSSSSSSSSSSZZSSSSSSSSSSSSSSSZ",
  "SSSSSSSSSSSSSSSSSSSSSSSZZZZZSZQZZZSSZZZZZZZZSSSSSSSSSSSZZSSSSSSSZSSZZZZQ",
  "SQSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSZZZZZZZZSSSSSSSSSSZSSSSSSSSSSSSSSSSS",
  "QQQQSQSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSZZZZZZZZSSSSSSSSSSZSSSSSSSSSSSSSSSSS",
  "SSSSSSQQQQSQQSQQSSQQQZSSSSQSSSSSSSSSZZZZZZZZSSSSQQQQQQQZQZZZQQZZQQQQQZQZ",
  "SSSSSSSSSSQQSSSSSSSQQZZZZZZZQSSSSSSSZZZZZZZZSSSSSZSSSSZZZZSSSSSSSSSSZZSZ",
  "SSSSSSSSSSSSSSSSSSSSSSZSSSZZSSSSSSSSZZZZZZZZZZZZSSSSZZZZZQSSZZZZQZZZZZZZ",
  "QSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSZZZZZZZZSSSSSSSSSSSSSSSSSSSSSSSSSSSS",
  "QSSSSSSSSSSSSSSSSSSSSSSSSSSZSSSSSSSSZZZZZZZZSSSSSSSSSSSZZZSSSSSSSSSZZSSS",
  "ZZSSSSSSSSSZZZZZQZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ",
  "ZQQQZSQQSSSSSSSSSSSSSSSSSSSSSSSSSQQSZZZZZZZZSSSSSSSSZZSSSSSSSSSSSSSSSZZZ",
  "SSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSSZZZZZZZZZZZZZZZZZZZZZZZZZZQZZZZZZZZQ",
  "QQQSSSSQQQQSSSSSSSSSZZZZZZZZZZQSSSSSZZZZZZZZSSSZZZZZZZZZZZZZZZZZZZZZZZZZ",
  "SSSSSSSSSSSSSSSSSSSSSSSSSSSZSSSSSSSSZZZZZZZZSSSSSZZZZZZZZZZZSSSSSSZZZZQQ" ;

 vComponentQCA =
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 523, 523, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 0, 515, 0,
  523, 523, 0, 523, 523, 0, 0, 523, 523, 523, 0, 0, 523, 523, 523, 523, 523, 
    515, 515, 515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 523, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 
    515, 0, 0, 0, 515, 515, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 515, 515, 0, 
    0, 0, 0, 0, 0, 0,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 523, 0, 515, 0, 0, 0, 0, 0, 0, 515, 0, 0, 515, 515, 515, 515, 515, 
    515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 0, 0, 515, 515, 
    515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 515, 0, 0, 0, 0, 0, 0, 0, 0,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 523, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 0,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 0, 515, 515, 
    515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 0, 515, 515, 515, 515, 515, 515, 515, 515, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 523, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 523, 523, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 
    515, 515, 0, 0, 0, 0, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 0, 515, 0,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 0, 0, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 0, 0, 0, 0, 0,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 523, 523, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 515, 0, 0,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 523, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 0, 515, 0,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 523, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 0, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 515, 0,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 515, 0, 515, 0, 0, 
    0, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 0, 0, 515, 515, 515, 515, 515, 515, 515, 0, 515, 515, 
    0, 0, 0, 0, 515,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 523, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 515, 515,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 515, 515,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 523, 523, 515, 515, 515, 0, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 515, 0, 0, 0, 515, 515, 0, 0, 515, 
    515, 515, 515, 515, 0, 515, 0,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 515, 
    515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 515, 515, 0, 
    515, 515, 515, 515, 0, 0, 0, 0, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 0, 0, 515, 0,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 523, 515, 515, 515, 515, 515, 0, 515, 515, 515, 0, 0, 515, 515, 515, 
    515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 
    515, 515, 0, 0, 0, 0, 0, 515, 515, 515, 0, 0, 0, 0, 515, 0, 0, 0, 0, 0, 
    0, 0,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 523, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 0, 515, 515, 
    515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 0, 0, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 0, 0, 515, 515, 515,
  0, 0, 523, 523, 523, 523, 523, 523, 523, 523, 523, 0, 0, 0, 0, 0, 523, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 523, 523, 523, 0, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 515, 
    515, 515, 515, 515, 0, 0, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 0, 0, 0,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 523, 523, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 
    515, 515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 
    523, 523, 523, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 
    515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 523, 515, 
    515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 515, 0, 515, 515, 
    515, 515, 515, 515, 515, 515, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 515, 
    515, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 515, 515, 515, 515, 515, 515, 0, 0, 
    0, 0, 515, 515 ;

 vComponentQCR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 9, 0, 0, 0, 0, 0, 0, 0, 513, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 513, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 513, 0, 0, 0, 0, 0, 0, 0, 0,
  9, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  9, 9, 0, 0, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 513, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 513, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 513,
  0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  9, 9, 9, 9, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 9, 9, 9, 9, 0, 9, 9, 0, 513, 513, 0, 0, 513, 513, 513, 0, 
    0, 0, 0, 0, 513, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 513, 513, 513, 513, 513, 513, 513, 0, 513, 0, 0, 0, 513, 513, 0, 0, 
    513, 513, 513, 513, 513, 0, 513, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 9, 0, 0, 0, 0, 0, 0, 0, 513, 513, 0, 0, 0, 
    0, 0, 0, 0, 513, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 513, 0, 0, 0, 0, 0, 0, 513, 0, 0, 0, 0, 0, 0, 0,
  9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 513, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 513, 9, 9, 0, 0, 9, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 513, 513, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 513, 0, 0, 0, 0, 0, 0, 0, 0, 513,
  9, 9, 9, 0, 0, 0, 0, 9, 9, 513, 513, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 513, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 513, 513 ;

 vComponentICA =
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 0, 3, 3, 0, 0, 3, 3, 3, 0, 0, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 3, 3, 3, 0, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 vComponentICR =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 0, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 3, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 3, 3, 3, 3, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 3, 3, 0, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  3, 3, 3, 0, 0, 0, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 wComponent =
  0, -0.01, 0, 0.01, 0, -0.02, -0.02, -0.03, -0.05, -0.08, -0.06, -0.05, 
    -0.03, 0.02, 0.04, 0.02, -0.02, -0.04, -0.05, -0.05, 0, 0.02, 0.04, 0.03, 
    0.04, 0.02, 0, 0.01, 0.03, 0.02, 0.04, 0.07, 0.08, 0.07, 0.06, 0.05, _, 
    _, _, _, _, _, _, _, 0.05, 0.06, 0.08, 0.04, 0.04, 0.03, 0.03, -0.01, 
    0.02, 0.03, 0.1, 0.08, 0.11, 0.22, 0.14, 0.15, 0.06, 0.07, 0.07, 0.08, 
    0.11, 0.08, 0.07, -0.01, _, _, -0.17, _,
  -1.37, -0.07, _, -0.06, -0.09, _, _, -0.16, 0.03, 0, _, _, -0.05, 0.03, 
    -0.13, -0.26, -0.37, -0.36, -0.2, -0.13, -0.2, -0.16, -0.04, -0.02, 
    -0.03, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  -0.04, -0.04, -0.04, -0.06, -0.07, -0.09, -0.09, 0.03, 0.08, 0.18, 0.1, 
    0.11, 0.11, 0.13, 0.11, 0.13, -0.07, -0.07, -0.11, -0.11, -0.07, -0.01, 
    -0.02, 0.02, -0.12, 0.01, 0.09, -0.06, 0.02, 0.03, 0.03, 0.03, 0.02, 
    0.01, -0.01, 0, _, _, _, _, _, _, _, _, -0.02, -0.01, 0.01, 0.04, _, _, 
    _, 0.18, 0.38, _, _, _, _, _, _, _, 0.05, 0.09, 0.1, 0.05, -0.11, _, _, 
    _, _, _, _, _,
  0, 0, 0.03, -0.03, -0.06, -0.06, -0.02, -0.01, 0, -0.01, -0.02, -0.06, 
    -0.08, -0.11, -0.09, -0.04, 0, _, 0.07, _, _, _, _, _, _, -0.05, _, _, 
    -0.03, -0.04, -0.04, -0.01, -0.02, 0.02, 0.04, 0.04, _, _, _, _, _, _, _, 
    _, 0.02, 0.01, 0.01, _, _, -0.07, -0.06, -0.05, -0.04, -0.04, -0.07, 
    -0.03, _, _, _, _, _, _, _, -0.02, _, _, _, _, _, _, _, _,
  0.14, 0.2, 0.15, 0.1, 0.14, 0.11, 0.13, 0.13, 0.14, 0.21, 0.21, 0.16, 0.12, 
    -0.02, 0.19, 0.24, 0.38, -0.05, -0.25, -0.21, -0.28, -0.52, -0.59, -0.54, 
    -0.57, -0.51, -0.49, -0.49, -0.46, -0.42, -0.41, -0.39, -0.35, -0.32, 
    -0.29, -0.25, _, _, _, _, _, _, _, _, -0.19, -0.15, -0.13, -0.13, -0.13, 
    -0.13, -0.11, -0.09, -0.1, -0.08, -0.09, -0.06, -0.06, 0, -0.08, -0.11, 
    -0.12, -0.15, -0.14, -0.09, 0.11, 0.12, 0.12, 0.11, 0.08, 0.05, 0.19, _,
  -0.2, -0.29, -0.24, -0.17, -0.1, -0.15, -0.17, -0.21, -0.25, -0.3, -0.29, 
    -0.28, -0.32, -0.25, -0.14, -0.12, -0.08, -0.12, -0.07, 0.02, -0.02, 
    -0.02, -0.03, 0.06, -0.02, -0.12, -0.09, _, 0, -0.08, -0.24, -0.26, 
    -0.13, -0.25, -0.18, -0.09, _, _, _, _, _, _, _, _, -0.04, -0.01, -0.02, 
    0, -0.09, -0.22, -0.33, -0.48, 0.12, _, -0.12, 0.07, 0.1, 0.09, 0.05, 
    -0.13, -0.13, 0.01, _, _, _, _, _, _, _, _, _, _,
  _, _, -0.01, -0.1, 0.05, 0.06, 0.05, 0.1, -0.09, -0.06, -0.24, -0.38, 
    -0.55, -0.51, -0.23, 0.03, -0.08, -0.11, 0.01, 0.08, 0.17, 0.2, 0.12, 
    0.2, 0.21, 0.39, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  0.09, -0.02, -0.02, -0.02, -0.01, -0.03, -0.03, 0, -0.03, -0.06, -0.03, 
    -0.01, -0.02, -0.02, 0, 0.04, 0.11, 0.14, 0.13, 0.13, 0.16, 0.19, 0.22, 
    0.23, 0.22, 0.23, 0.25, 0.17, 0.06, 0.02, -0.01, -0.02, -0.02, -0.05, 
    -0.11, -0.17, _, _, _, _, _, _, _, _, -0.22, -0.22, -0.2, -0.18, -0.18, 
    -0.18, -0.15, -0.14, -0.11, -0.13, -0.2, -0.16, -0.12, -0.08, -0.07, 
    -0.07, -0.09, -0.06, -0.03, -0.02, -0.02, 0, 0.02, 0.01, 0, -0.03, 0.02, 
    0.06,
  0.05, 0.04, 0.02, -0.01, 0.06, 0.09, 0.1, 0.11, 0.09, 0.14, 0.19, 0.17, 
    0.12, 0.12, 0.04, 0.03, 0.05, 0.05, 0.07, 0.07, 0.02, 0.05, 0.04, 0.04, 
    0.01, 0.08, 0.07, 0.11, 0.06, 0.08, 0.07, 0.01, 0, 0, -0.01, -0.02, _, _, 
    _, _, _, _, _, _, -0.03, -0.03, 0, 0.03, 0.04, _, _, _, _, 0.17, 0.25, 
    0.15, 0.12, 0.08, 0.1, 0.02, 0.05, -0.1, -0.02, -0.05, 0, -0.01, 0.01, 
    0.16, 0.31, _, 0.05, _,
  0.49, -0.01, -0.02, -0.01, 0.04, -0.01, -0.04, -0.06, -0.04, -0.11, -0.2, 
    -0.23, -0.21, -0.19, -0.14, -0.02, -0.07, -0.04, 0.02, 0.06, -0.08, 0, 
    -0.06, 0.01, -0.03, 0.11, 0.09, 0.12, -0.16, -0.2, -0.11, -0.18, -0.1, 
    -0.11, -0.09, 0.03, _, _, _, _, _, _, _, _, 0.05, 0.01, 0.06, 0.03, 0.02, 
    0.16, 0.41, -0.03, -0.01, _, _, _, 0.24, 0.32, _, 0.26, 0.03, 0, -0.02, 
    0, -0.07, -0.16, -0.21, _, _, _, _, _,
  -0.04, 0.05, -0.02, -0.03, -0.06, -0.02, 0.01, 0.03, 0.03, 0.04, 0.1, 0.16, 
    0.19, 0.34, 0, 0.02, -0.04, 0.04, -0.04, -0.15, -0.16, -0.15, -0.12, 
    -0.13, -0.13, -0.14, -0.11, 0.25, -0.05, 0.01, 0.1, 0.16, 0.2, 0.19, 
    0.23, 0.3, _, _, _, _, _, _, _, _, 0.32, 0.15, 0.15, 0.31, 0.22, 0.16, 
    0.09, 0.08, 0.11, 0.06, 0.03, 0, 0.01, -0.02, -0.04, -0.06, -0.08, -0.09, 
    -0.03, -0.04, -0.08, -0.03, 0.03, 0.11, 0.15, 0.09, _, _,
  0.13, 0.1, 0.09, 0.12, -0.02, -0.05, -0.06, -0.13, -0.13, -0.17, -0.17, 
    -0.2, -0.19, -0.2, -0.18, -0.15, -0.11, -0.06, 0.04, 0.05, 0.06, 0.14, 
    0.09, 0.16, 0, 0.17, 0.15, 0.32, 0.19, 0.19, 0.15, 0.12, 0.12, 0.12, 
    0.11, 0.09, _, _, _, _, _, _, _, _, 0.07, 0.07, 0.07, 0.07, 0.12, 0.13, 
    0.12, 0.06, 0.12, 0.04, 0, -0.06, -0.07, -0.06, _, 0.18, 0.12, 0.06, 
    0.09, -0.02, -0.04, -0.04, 0.02, -0.21, -0.24, _, 0.02, _,
  0.21, 0.2, 0.54, 0.34, 0.21, 0.2, 0.3, 0.08, 0.13, 0.19, 0.14, 0.02, 0.21, 
    0.26, 0.12, 0.57, 0.54, 0.31, 0.72, 1.73, 1.58, 0.68, 0.06, 0.22, 0.22, 
    0.18, 0.09, -0.16, -0.35, -0.48, -0.56, -0.59, -0.57, -0.5, -0.43, -0.37, 
    _, _, _, _, _, _, _, _, -0.34, -0.32, -0.25, -0.18, -0.15, -0.25, -0.02, 
    0.32, -0.01, _, _, _, _, -0.67, 0.03, 0.29, -0.18, 0.3, 0.15, 0.04, 
    -0.09, _, _, -0.12, -0.03, 0.18, _, _,
  0.03, -0.08, -0.13, -0.1, -0.11, -0.08, -0.04, 0.02, 0.06, 0.13, 0.26, 
    0.39, 0.48, 0.58, 0.68, 0.63, 0.79, 0.7, 0.72, 0.81, 0.8, 0.78, 0.5, _, 
    _, _, _, _, 0.6, _, 1.67, _, _, _, 0.41, 0.39, _, _, _, _, _, _, _, _, 
    0.31, 0.01, 0.02, 0.02, 0.03, 0.04, 0.02, -0.04, -0.06, -0.19, -0.29, _, 
    _, -0.01, 0.36, 0.29, 0.23, 0.23, 0.14, 0.25, _, 0.09, -0.21, _, _, _, _, 
    0.05,
  0.12, 0.14, 0.19, 0.14, 0.12, 0.11, -0.04, -0.06, -0.02, -0.01, 0.01, 
    -0.01, -0.08, -0.04, -0.06, -0.1, -0.13, -0.09, -0.09, -0.09, -0.09, 
    -0.08, -0.05, -0.03, 0.05, 0.07, 0.09, 0.1, 0.09, 0.09, 0.07, 0.05, 0.07, 
    0.07, 0.06, 0.04, _, _, _, _, _, _, _, _, 0.05, 0.05, 0.07, 0.09, 0.1, 
    0.1, 0.09, 0.07, 0.06, 0.07, _, 0.18, 0.12, 0.11, 0.13, 0.08, 0.09, 0.08, 
    0.1, 0.1, 0.1, 0.1, 0.02, -0.02, -0.02, -0.02, 0.02, 0.03,
  0.01, 0.02, 0, -0.01, 0.02, 0.15, 0.07, -0.01, -0.01, -0.01, 0.01, 0.01, 0, 
    0.01, 0.12, 0.16, 0.19, 0.22, 0.13, 0.02, -0.03, -0.01, -0.13, -0.21, 
    -0.18, -0.17, -0.26, -0.13, -0.18, -0.18, -0.18, -0.17, -0.17, -0.19, 
    -0.3, -0.38, _, _, _, _, _, _, _, _, -0.44, -0.42, -0.39, -0.33, -0.28, 
    -0.24, -0.17, -0.16, -0.13, -0.32, _, -0.42, -0.22, -0.15, -0.12, -0.04, 
    0.02, 0.03, 0.04, 0.4, 0.15, 0.39, -0.26, -0.31, -0.17, -0.14, -0.03, 0.03,
  0.09, 0.06, 0.08, 0.09, 0.07, 0.06, 0.03, 0.15, 0.41, 0.42, -0.02, -0.14, 
    -0.16, -0.19, -0.09, -0.01, -0.04, -0.04, -0.03, -0.02, -0.14, _, -0.04, 
    -0.06, -0.07, -0.04, -0.01, 0.02, 0.05, 0.03, 0.03, 0.03, 0.06, 0.05, 
    0.05, 0.04, _, _, _, _, _, _, _, _, 0.02, 0.03, -0.01, -0.11, -0.32, 
    -0.24, -0.05, 0, -0.13, _, _, _, 0, _, _, _, _, -0.26, _, _, 0.03, 0.08, 
    -0.07, 0.04, 0.01, _, -0.03, _,
  0.03, -0.05, -0.03, -0.01, -0.04, 0.04, 0.05, 0.16, 0.12, 0.2, 0.31, 0.18, 
    0.19, 0.54, 0.12, 0.18, 0.04, 0.06, -0.08, 0.03, 0.01, _, _, _, _, _, _, 
    _, -0.23, -0.46, -0.02, _, -0.18, _, _, -0.57, _, _, _, _, _, _, _, _, 
    -1.15, -0.39, -0.79, -0.62, -0.54, _, _, -0.19, 0.06, _, _, _, _, _, 
    -0.33, -0.04, -0.07, 0.1, -0.08, _, _, _, -0.58, _, _, _, _, _,
  0.14, 0.1, 0.04, 0.07, 0.11, 0.14, 0.14, 0.26, 0.41, 0.32, 0.15, 0.14, 
    0.15, 0.21, 0.23, 0.2, 0.23, 0.3, 0.11, 0.15, -0.02, 0.01, _, -0.1, 
    -0.04, 0, _, _, -0.12, -0.12, -0.13, -0.11, -0.02, 0.04, -0.1, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, -0.08, 0.15, 0.21, 0.19, _, _, _, _, _, _, 
    0.04, _, _, _, _, _, -0.19, _, _, _, _, _, _, _,
  -0.06, -0.08, -0.09, -0.07, -0.08, -0.08, -0.05, -0.05, -0.04, -0.03, 
    -0.04, -0.05, -0.04, -0.09, -0.04, -0.05, -0.09, -0.1, -0.07, -0.1, 
    -0.12, -0.08, -0.08, -0.07, -0.06, -0.07, -0.07, -0.03, -0.03, -0.01, 
    -0.01, -0.01, -0.03, -0.05, -0.06, -0.05, _, _, _, _, _, _, _, _, -0.05, 
    -0.07, -0.1, -0.13, -0.12, -0.12, -0.16, -0.13, -0.14, -0.11, -0.18, 
    -0.04, -0.19, -0.07, -0.19, -0.14, -0.19, -0.19, -0.12, -0.06, 0, 0.1, 
    0.12, 0.07, 0.05, -0.11, -0.14, -0.11,
  -0.05, -0.02, 0.16, 0.03, 0.14, 0.14, 0.05, -0.09, -0.13, -0.08, -0.12, 
    -0.19, -0.26, -0.32, -0.44, -0.48, -0.51, -0.55, -0.78, -1.04, -1.05, 
    -1.1, -1.13, -1.16, -1.17, -1.09, -1.16, _, -1.03, -1.02, -1, -0.98, 
    -0.91, -0.85, -0.81, -0.77, _, _, _, _, _, _, _, _, -0.74, -0.66, -0.61, 
    -0.56, -0.54, -0.39, -0.24, -0.06, _, 0.1, 0.11, _, _, _, 0.18, 0.25, 
    0.37, 0.38, 0.36, 0.38, 0.37, 0.46, _, _, _, 0.25, 0.05, 0.02,
  _, _, 0.1, 0, -0.19, -0.19, -0.19, -0.29, 0, -0.1, -0.29, _, _, _, _, _, 0, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, 0, -0.01, 0.01, _, 0.41, 0.35, 0.28, 0.38, 0.16, 0.17, 0.16, 0.12, 0.16, 
    0.1, -0.14, -0.33, -0.55, -0.64, -0.54, -0.45, -0.49, -0.65, -0.64, 
    -1.63, -1.87, -1.27, -0.67, -1.07, -1.1, -0.96, -0.92, -0.67, -0.65, 
    -1.08, -0.73, _, _, _, _, _, _, _, _, -0.85, -0.74, -0.56, -0.44, -0.28, 
    -0.19, -0.11, -0.07, _, _, -0.04, 0.06, 0.2, 0.31, 0.31, 0.3, 0.28, 0.24, 
    0.22, 0.12, 0.06, 0.13, 0.13, 0.1, 0.16, _, _, _,
  0.08, 0.08, 0.11, 0.07, 0.07, 0.07, -0.21, -0.05, -0.12, -0.2, -1.14, 0.02, 
    0.06, -2.74, -1.6, -0.42, -0.66, -0.49, -0.29, -0.14, -0.16, -0.17, 
    -0.05, -0.22, -0.12, -0.1, -0.09, -0.59, -0.1, -0.08, 0, 0.03, -0.03, 
    0.11, -0.22, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.01, -0.02, -0.05, -0.04, -0.05, -0.07, -0.13, -0.11, -0.34, -0.03, -0.01, 
    0.01, 0.04, 0.01, -0.03, -0.04, 0.04, 0, 0.02, 0.08, _, _, _, _, _, _, _, 
    _, _, _, _, _, 0.34, 0.17, 0.22, 0.15, _, _, _, _, _, _, _, _, 0.1, 0.16, 
    0.06, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _,
  -0.06, 0.02, 0.05, 0.07, 0.08, 0.17, 0.1, 0.09, 0.12, 0, 0.02, 0.08, -0.06, 
    -0.1, -0.06, -0.09, -0.08, -0.07, -0.16, -0.15, -0.24, -0.14, -0.17, 
    -0.13, -0.2, -0.14, -0.07, _, -0.1, -0.1, -0.04, -0.03, 0.02, 0.03, 0.09, 
    0.11, _, _, _, _, _, _, _, _, 0.13, 0.17, 0.13, -0.01, -0.09, _, _, _, _, 
    _, _, _, _, _, _, _, _, -0.32, -0.58, -0.46, -0.31, -0.34, _, _, _, _, 
    0.04, 0.02 ;

 uvQualityCode =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, 0, _,
  0, 4, _, 0, 0, _, _, 0, 0, 2, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, _, 
    _, _, 0, 0, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, _, 0, _, _, _, _, _, _, 
    0, _, _, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, _, _, 
    0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, 8, _, _, _, _, _, _, _, _,
  4, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _,
  4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, _, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, _, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _,
  _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  4, 4, 0, 0, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, _,
  0, 0, 0, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, _, _, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, 
    _, _, _, 0, _, 2, _, _, _, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, _, _, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, _, 8,
  0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  4, 4, 4, 4, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 0, 4, 4, 0, 2, 2, 0, 0, 2, 8, 2, _, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 2, 
    8, 8, 8, 8, 8, 8, _, 8, _, _, _, 8, 8, _, _, 8, 8, 8, 8, 8, _, 8, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 0, 0, 0, 0, 0, 0, 0, 2, 2, _, _, _, _, 
    _, _, _, 2, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    _, 0, 0, 0, 0, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, 0, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 
    0, _, _, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, 0, 
    0, 0, 0, _, _, _, _, _, 2, 0, 0, _, _, _, _, 2, _, _, _, _, _, _, _,
  4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, _, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, 0, 0, 0,
  _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, 8, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 2, 4, 4, _, 0, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    0, 0, 0, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, 8, _, _, _, _, _, _, _, _, 8,
  4, 4, 4, 0, 0, 0, 0, 4, 4, 2, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, 
    _, _, _, _, _, 2, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, _, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 0, _, _, _, _, 8, 8 ;

 wQualityCode =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, 0, _,
  0, 0, _, 0, 0, _, _, 0, 0, 0, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, _, 
    _, _, 0, 0, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, _, _, _, _, _, _, 
    0, _, _, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, _, _, 
    0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, 0, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, _, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, _, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _,
  _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, _, _, _, 0, 0, _, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, _, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, _, _, 0, 0, 0, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, 
    _, _, _, 0, _, 0, _, _, _, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, _, _, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, _, _, _, _, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, _, _, _, 0, _, _, _, _, 0, _, _, 0, 0, 0, 0, 0, _, 0, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, 
    _, _, _, 0, 0, 0, _, 0, _, _, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    _, _, 0, 0, _, _, _, _, _, 0, 0, 0, 0, 0, _, _, _, 0, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, 0, 0, 
    0, _, _, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, 0, 
    0, 0, 0, _, _, _, _, _, _, 0, _, _, _, _, _, 0, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, _, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    0, 0, 0, _, 0, 0, _, _, _, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, 0, 0, 0,
  _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, 0, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0, 0, 0, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    0, 0, 0, _, _, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, 
    _, _, _, _, _, _, _, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, _, 0, 0, 0, 0, 0, 0, 0, 0, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, 
    _, _, _, _, _, _, _, _, _, _, _, _, 0, 0, 0, 0, 0, _, _, _, _, 0, 0 ;

 HorizSpStdDev =
  7.29, 4.84, 2.56, 2.56, 1.96, 1.44, 1.69, 2.25, 2.89, 2.25, 1.96, 1.69, 
    1.96, 1.96, 1.44, 1.69, 1.69, 1.69, 1.44, 1.44, 1.44, 1.96, 1.96, 2.25, 
    2.25, 1.69, 1.44, 0.81, 4, 4, 4, 3.61, 3.61, 3.61, 3.61, 4, _, _, _, _, 
    _, _, _, _, 4.41, 4.41, 4, 3.61, 3.61, 2.89, 2.89, 3.24, 2.89, 2.56, 4, 
    4.41, 4, 3.24, 4, 4, 4.84, 5.29, 6.25, 5.29, 4.41, 4, 4, 3.61, _, _, 
    3.24, _,
  28.09, 4, _, 5.29, 6.25, _, _, 4.41, 4.41, 4.84, _, _, 3.24, 4, 4, 4.41, 
    4.84, 2.56, 2.89, 7.29, 4, 3.61, 3.24, 2.56, 2.56, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  1.96, 2.25, 2.89, 2.56, 1.44, 1.69, 2.25, 2.25, 2.25, 2.56, 1.21, 1.69, 
    2.25, 1.96, 1.96, 1.69, 0.64, 1.44, 2.56, 2.25, 2.25, 1.96, 1.96, 1.69, 
    2.56, 2.25, 2.25, 1.96, 2.56, 2.56, 2.25, 2.56, 3.24, 2.89, 3.24, 2.89, 
    _, _, _, _, _, _, _, _, 2.56, 3.24, 3.24, 4, _, _, _, 2.89, 3.24, _, _, 
    _, _, _, _, _, 4, 4, 3.61, 3.24, 3.24, _, _, _, _, _, _, _,
  6.25, 4.41, 4, 2.25, 3.24, 4.41, 3.24, 3.24, 2.89, 2.56, 2.89, 4, 4.41, 
    2.89, 2.89, 2.56, 2.25, _, 2.56, _, _, _, _, _, _, 2.56, _, _, 2.56, 4, 
    2.56, 2.56, 2.56, 3.24, 3.24, 2.89, _, _, _, _, _, _, _, _, 3.24, 4, 
    6.25, _, _, 3.24, 3.61, 3.61, 3.61, 3.24, 3.61, 3.24, _, _, _, _, _, _, 
    _, 6.25, _, _, _, _, _, _, _, _,
  14.44, 6.76, 9, 6.76, 5.29, 3.24, 2.25, 1.69, 1.44, 0.25, 0.81, 1.21, 1.44, 
    0.36, 1.96, 1.96, 2.25, 0.49, 2.56, 1.44, 1.44, 1.44, 1.21, 1.21, 1.44, 
    2.25, 2.25, 1.96, 3.61, 3.24, 2.89, 2.89, 2.89, 2.89, 2.89, 2.89, _, _, 
    _, _, _, _, _, _, 2.89, 2.89, 2.56, 3.24, 4, 4, 4.41, 4.41, 4.41, 3.24, 
    3.24, 4, 4.84, 4.84, 5.29, 6.25, 6.25, 6.76, 6.25, 5.29, 4, 4.84, 5.29, 
    4.41, 4.41, 4.41, 4.84, _,
  9, 7.29, 3.24, 1.69, 2.25, 4.41, 2.25, 1.96, 1.44, 1.21, 0.64, 1, 0.49, 
    0.81, 1, 1.44, 1.21, 1, 1.21, 1.44, 0.81, 1.21, 1, 0.81, 0.81, 1, 1.69, 
    _, 4.84, 5.76, 2.89, 4.41, 3.61, 3.61, 3.61, 3.61, _, _, _, _, _, _, _, 
    _, 3.24, 2.89, 2.89, 3.24, 3.24, 3.24, 4, 1, 2.25, _, 4, 4, 3.61, 3.61, 
    3.24, 4.41, 5.76, 5.76, _, _, _, _, _, _, _, _, _, _,
  _, _, 1.69, 2.56, 2.56, 1.44, 1.21, 2.56, 1.96, 2.25, 0.81, 1.96, 1, 1.69, 
    0.64, 1, 0.81, 1, 0.49, 1.96, 2.25, 1.21, 1.21, 1, 0.64, 1, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  12.96, 15.21, 6.25, 4.84, 9, 7.84, 2.25, 2.25, 3.24, 1.69, 1.69, 1.21, 
    0.81, 2.56, 1, 1, 1, 1.21, 1, 1.44, 1, 1, 1.96, 1.44, 0.36, 0.49, 0.64, 
    1.21, 3.24, 3.24, 2.89, 2.89, 2.89, 2.56, 1.96, 2.25, _, _, _, _, _, _, 
    _, _, 2.25, 2.25, 1.96, 1.96, 2.25, 2.56, 3.61, 3.61, 2.89, 3.61, 4, 
    3.61, 3.24, 4.41, 4.84, 5.76, 6.76, 6.25, 4.41, 3.61, 4.41, 4.41, 4.84, 
    4.84, 4.41, 4.41, 4.41, 4,
  4.41, 4, 4.41, 6.76, 10.89, 3.61, 2.89, 2.56, 2.56, 2.25, 1.96, 1.69, 1.96, 
    2.56, 3.61, 1.69, 0.81, 1.69, 1, 0.81, 1.69, 2.25, 1, 1.44, 0.81, 1, 
    0.25, 1.96, 2.56, 3.24, 2.89, 2.56, 2.56, 3.61, 4, 4, _, _, _, _, _, _, 
    _, _, 4, 4, 4.84, 5.29, 2.89, _, _, _, _, 4, 2.89, 3.61, 3.24, 3.24, 
    3.61, 2.89, 3.24, 4.41, 4.84, 4, 4, 3.61, 4, 3.61, 4, _, 3.24, _,
  6.25, 3.24, 6.76, 7.84, 4.84, 4.41, 2.25, 1.96, 2.89, 3.24, 1.21, 0.81, 
    1.96, 4, 3.24, 3.61, 2.56, 0.81, 0.81, 0.09, 2.25, 1.21, 0.49, 1.96, 
    1.44, 1.44, 0.81, 1, 3.24, 0.25, 3.24, 2.25, 1.96, 1.96, 1.21, 2.56, _, 
    _, _, _, _, _, _, _, 2.89, 2.89, 2.89, 3.24, 2.89, 2.89, 3.24, 4, 4, _, 
    _, _, 4.41, 5.76, _, 5.29, 4, 4.41, 5.29, 4, 4, 4.41, 3.61, _, _, _, _, _,
  0.36, 1.96, 1.96, 1.96, 1.96, 1.96, 1.96, 1.96, 1.96, 2.56, 3.24, 1.96, 1, 
    2.25, 1, 1, 0.81, 1.21, 1, 2.25, 1.44, 1.21, 1.44, 1, 1, 1.44, 1.96, 
    1.44, 2.56, 2.56, 2.89, 2.89, 2.56, 3.24, 3.61, 3.24, _, _, _, _, _, _, 
    _, _, 3.61, 2.56, 2.89, 3.61, 3.61, 2.89, 1.96, 2.25, 2.56, 3.24, 4, 
    3.61, 3.24, 3.61, 3.61, 4, 4.41, 5.76, 5.29, 6.25, 6.76, 6.76, 5.29, 
    4.41, 4.84, 3.61, _, _,
  3.61, 2.89, 2.56, 3.61, 1.21, 1.44, 1.21, 0.64, 1.96, 0.81, 1, 1.21, 2.25, 
    1.21, 0.81, 0.81, 1, 1, 0.49, 0.36, 0.36, 1.21, 0.49, 1.44, 1.44, 1.69, 
    2.56, 2.25, 4, 4, 3.24, 1.96, 2.25, 3.61, 2.25, 2.25, _, _, _, _, _, _, 
    _, _, 1.96, 2.25, 2.89, 1.96, 2.89, 3.61, 3.24, 2.89, 2.25, 2.56, 1.44, 
    2.56, 1.96, 3.24, _, 6.25, 5.76, 4.84, 5.29, 5.29, 5.76, 4, 4, 3.61, 4, 
    _, 2.89, _,
  1.44, 1.21, 5.29, 4.41, 2.89, 1.44, 1.21, 1.44, 1.21, 1.44, 1.21, 2.25, 
    3.24, 1.96, 0.64, 3.61, 2.25, 3.24, 5.29, 3.24, 1.44, 1.44, 0.64, 1, 1, 
    1, 0.81, 2.25, 1.69, 1, 1.44, 1.69, 2.56, 2.25, 1.44, 1.21, _, _, _, _, 
    _, _, _, _, 0.49, 0.81, 1.44, 1.96, 1.96, 0.81, 1.44, 2.25, 3.24, _, _, 
    _, _, 6.25, 4.84, 5.76, 6.76, 7.29, 5.76, 4, 4.41, _, _, 4.84, 5.76, 
    5.29, _, _,
  2.89, 4, 3.24, 3.24, 3.61, 4.41, 2.25, 1.69, 4.84, 1.21, 1.96, 1.69, 1.96, 
    1.44, 1.21, 0.64, 1.44, 1, 1, 2.56, 0.81, 1.96, 1, _, _, _, _, _, 2.89, 
    _, 1.21, _, _, _, 2.89, 2.89, _, _, _, _, _, _, _, _, 2.56, 3.24, 4.41, 
    5.76, 6.25, 6.76, 6.25, 5.76, 4.84, 5.29, 4.84, _, _, 4, 4.41, 4, 4.84, 
    4, 3.24, 2.56, _, 8.41, 8.41, _, _, _, _, 9,
  3.61, 6.25, 1.69, 4.41, 4.41, 7.29, 2.56, 4, 3.24, 2.56, 2.89, 2.89, 2.25, 
    2.25, 1.69, 1.69, 1.69, 1.44, 1.69, 1.96, 1.96, 1.69, 1.69, 1.44, 0.81, 
    0.81, 0.64, 1.21, 2.25, 2.89, 3.61, 4.84, 5.76, 4.84, 3.61, 2.56, _, _, 
    _, _, _, _, _, _, 2.25, 1.96, 2.25, 2.89, 2.56, 2.89, 3.24, 4, 4.84, 
    2.56, _, 3.61, 2.56, 2.56, 3.24, 4, 4.41, 4, 4.84, 4.84, 4.84, 5.76, 
    5.76, 4.41, 5.29, 5.76, 5.76, 4.41,
  16, 14.44, 7.29, 8.41, 7.84, 7.29, 5.29, 3.61, 4, 3.24, 2.56, 2.25, 2.56, 
    1.96, 4, 2.89, 1.96, 3.24, 2.25, 1.96, 1.44, 0.81, 1, 0.25, 1.44, 1.44, 
    1.44, 1.69, 5.76, 5.29, 4.41, 4, 4.41, 5.76, 4.84, 4.84, _, _, _, _, _, 
    _, _, _, 5.29, 3.61, 3.61, 4.84, 4.84, 4.84, 4.41, 4.41, 4.41, 4.41, _, 
    7.84, 7.84, 8.41, 7.84, 7.29, 7.29, 6.76, 6.76, 4.84, 5.29, 3.61, 4, 
    6.25, 5.29, 7.29, 7.84, 7.29,
  2.25, 1.69, 2.89, 5.29, 5.76, 7.29, 7.29, 7.29, 6.76, 7.84, 8.41, 8.41, 
    9.61, 3.61, 2.89, 2.56, 4, 5.76, 5.29, 2.89, 1.96, _, 1.69, 1.44, 1.96, 
    1.44, 2.25, 1.44, 2.56, 2.89, 2.89, 2.89, 3.24, 2.89, 2.89, 2.89, _, _, 
    _, _, _, _, _, _, 3.24, 3.24, 3.24, 2.89, 2.56, 2.56, 1.96, 3.24, 4, _, 
    _, _, 4.41, _, _, _, _, 2.89, _, _, 2.89, 2.89, 2.89, 3.61, 3.24, _, 
    3.61, _,
  9, 5.76, 2.56, 6.76, 5.29, 4.84, 4.84, 3.61, 1.69, 4.41, 3.24, 1.69, 1.69, 
    6.25, 1.69, 1.69, 1.44, 0.64, 3.61, 1.21, 2.89, _, _, _, _, _, _, _, 
    3.61, 4, 3.61, _, 4, _, _, 3.61, _, _, _, _, _, _, _, _, 4, 4.84, 4.41, 
    4.41, 3.61, _, _, 4.41, 4, _, _, _, _, _, 5.76, 5.29, 5.29, 4.84, 3.24, 
    _, _, _, 3.61, _, _, _, _, _,
  3.24, 2.56, 3.24, 2.56, 0.81, 3.61, 1.21, 4, 2.89, 2.25, 2.89, 1, 0.64, 
    2.89, 5.29, 1.96, 1.69, 2.89, 1.44, 2.25, 0.49, 1, _, 1.21, 0.49, 1.69, 
    _, _, 3.24, 2.89, 3.61, 4.41, 4.84, 4.41, 5.29, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, 3.24, 3.61, 2.89, 2.25, _, _, _, _, _, _, 3.61, _, _, _, 
    _, _, 3.61, _, _, _, _, _, _, _,
  26.01, 2.25, 2.56, 2.56, 3.24, 3.24, 2.56, 3.24, 1.44, 1.69, 0.36, 0.25, 
    1.21, 2.89, 0.64, 0.64, 1, 0.81, 1.44, 1.69, 1.69, 1.44, 1, 1, 0.64, 
    0.64, 1, 0.64, 2.25, 2.25, 1.96, 1.96, 2.25, 2.25, 2.56, 2.56, _, _, _, 
    _, _, _, _, _, 2.25, 2.25, 2.89, 2.89, 3.24, 2.89, 3.24, 4, 4.41, 4.41, 
    4.41, 4.41, 4, 3.61, 4.84, 7.84, 6.25, 5.29, 4.84, 3.61, 3.61, 4.84, 
    5.29, 5.29, 5.29, 4.84, 5.29, 5.76,
  7.84, 5.29, 5.76, 5.76, 4.41, 4, 3.61, 2.25, 2.25, 1.96, 1.96, 1.96, 1.96, 
    2.25, 2.25, 1.69, 2.56, 2.89, 2.25, 1.44, 1.21, 1.44, 1.69, 1.69, 2.25, 
    2.89, 2.56, _, 6.25, 5.29, 4.41, 4.84, 2.89, 2.56, 2.56, 2.89, _, _, _, 
    _, _, _, _, _, 2.56, 2.56, 3.24, 4, 2.89, 4, 4.41, 4.41, _, 3.61, 3.61, 
    _, _, _, 4, 4.41, 5.76, 5.76, 5.76, 6.76, 5.76, 4.41, _, _, _, 3.61, 
    5.76, 5.29,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 30.25, 11.56, 16.81, _, 4.84, 8.41, 7.29, 4.41, 4, 3.61, 3.24, 5.29, 
    4.84, 4.41, 4.84, 5.76, 4.84, 5.29, 6.76, 7.29, 6.76, 6.25, 6.25, 1, 
    1.69, 7.84, 5.76, 13.69, 17.64, 16.81, 18.49, 12.96, 12.96, 14.44, 19.36, 
    _, _, _, _, _, _, _, _, 17.64, 18.49, 18.49, 13.69, 14.44, 16, 9.61, 9, 
    _, _, 15.21, 7.84, 8.41, 7.84, 7.84, 8.41, 11.56, 10.24, 8.41, 5.29, 
    5.29, 5.29, 5.29, 4.84, 4.41, _, _, _,
  2.25, 1.96, 2.56, 1.69, 5.29, 5.76, 1.69, 3.61, 2.56, 2.89, 6.76, 4.41, 
    4.84, 1.69, 3.61, 0.81, 1.21, 2.25, 1, 1.96, 1.96, 1.96, 3.61, 1.96, 
    1.44, 1.96, 1.21, 1.21, 3.61, 4, 5.29, 4.41, 3.24, 2.25, 1.96, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _,
  10.89, 9, 7.29, 4.41, 4, 4, 5.29, 6.76, 7.84, 4, 7.84, 5.76, 4.84, 4, 2.56, 
    2.25, 1.96, 1.44, 2.56, 2.56, _, _, _, _, _, _, _, _, _, _, _, _, 4, 
    4.41, 4.41, 6.76, _, _, _, _, _, _, _, _, 7.29, 7.84, 3.24, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  3.24, 1.96, 1.69, 2.56, 2.56, 2.89, 1.69, 3.24, 2.56, 2.56, 1.69, 2.25, 
    0.64, 0.64, 1.69, 1.69, 1, 0.49, 1, 1.21, 1.21, 1.69, 1, 1.69, 1.21, 
    1.21, 2.25, _, 5.29, 5.29, 4.41, 4.41, 4.41, 2.56, 2.56, 1.96, _, _, _, 
    _, _, _, _, _, 2.89, 3.61, 3.24, 4, 3.61, _, _, _, _, _, _, _, _, _, _, 
    _, _, 4.84, 5.29, 6.25, 7.29, 6.76, _, _, _, _, 4.84, 0.81 ;

 VertSpStdDev =
  0.2, 0.3, 0.3, 0.3, 0.3, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.3, 0.3, 
    0.3, 0.3, 0.3, 0.3, 0.3, 0.3, 0.3, 0.3, 0.3, 0.3, 0.4, 0.4, 0.4, 0.4, 
    0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, _, _, _, _, _, _, _, _, 0.4, 0.4, 0.5, 
    0.5, 0.6, 0.6, 0.6, 0.6, 0.6, 0.7, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 
    0.5, 0.5, 0.5, 0.4, 0.4, 0.4, 0.4, _, _, 0.5, _,
  6.3, 1.5, _, 0.8, 0.7, _, _, 0.5, 0.5, 0.4, _, _, 0.5, 0.3, 0.4, 0.4, 0.4, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.6, 0.4, 0.3, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.5, 0.4, 0.7, 0.4, 0.4, 0.3, 0.3, 0.3, 
    0.3, 0.4, 0.3, 0.3, 0.3, 0.3, 0.3, 0.3, 0.3, 0.3, 0.3, 0.3, 0.4, 0.3, 
    0.3, 0.3, 0.3, 0.3, 0.4, 0.4, 0.4, _, _, _, _, _, _, _, _, 0.4, 0.4, 0.4, 
    0.3, _, _, _, 0.4, 0.4, _, _, _, _, _, _, _, 0.5, 0.5, 0.5, 0.4, 0.5, _, 
    _, _, _, _, _, _,
  0.6, 0.5, 0.6, 0.5, 0.4, 0.4, 0.3, 0.3, 0.3, 0.3, 0.3, 0.3, 0.3, 0.2, 0.3, 
    0.3, 0.3, _, 0.3, _, _, _, _, _, _, 0.3, _, _, 0.3, 0.3, 0.4, 0.4, 0.4, 
    0.3, 0.4, 0.3, _, _, _, _, _, _, _, _, 0.3, 0.3, 0.4, _, _, 0.4, 0.4, 
    0.4, 0.4, 0.4, 0.5, 0.3, _, _, _, _, _, _, _, 0.5, _, _, _, _, _, _, _, _,
  0.7, 0.7, 0.6, 0.4, 0.4, 0.4, 0.4, 0.4, 0.5, 0.6, 0.7, 0.7, 0.8, 0.8, 0.8, 
    0.9, 0.8, 0.9, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.7, 0.7, 0.6, 0.7, 
    0.7, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, _, _, _, _, _, _, _, _, 0.6, 0.6, 0.6, 
    0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.7, 0.7, 0.8, 0.8, 0.8, 0.8, 0.7, 0.7, 
    0.6, 0.6, 0.6, 0.6, 0.5, 0.5, 0.5, 0.4, 0.4, 0.5, _,
  0.8, 0.7, 1, 1.1, 1.2, 0.9, 0.6, 0.4, 0.4, 0.4, 0.4, 0.5, 0.5, 0.4, 0.5, 
    0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.5, 0.5, 0.5, 0.5, _, 0.6, 0.6, 
    0.7, 0.7, 0.8, 0.8, 0.9, 0.9, _, _, _, _, _, _, _, _, 0.9, 0.9, 0.9, 0.8, 
    0.8, 0.8, 0.7, 0.8, 0.6, _, 0.4, 0.6, 0.6, 0.6, 0.6, 0.5, 0.4, 0.4, _, _, 
    _, _, _, _, _, _, _, _,
  _, _, 0.7, 0.7, 0.7, 0.6, 0.5, 0.7, 0.4, 0.4, 0.6, 0.7, 0.7, 0.3, 0.5, 0.6, 
    0.6, 0.5, 0.7, 0.6, 0.6, 0.5, 0.4, 0.4, 0.5, 0.6, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.9, 0.7, 0.6, 0.5, 0.5, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 
    0.4, 0.4, 0.4, 0.4, 0.3, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, _, _, _, _, _, _, _, _, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.6, 0.6, 0.6, 0.8, 1.1, 1.1, 1.1, 1.1, 1.1, 1, 0.8, 
    0.7, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.4,
  0.4, 0.4, 0.4, 0.4, 0.5, 0.5, 0.6, 0.6, 0.5, 0.6, 0.7, 0.5, 0.4, 0.4, 0.4, 
    0.3, 0.3, 0.3, 0.3, 0.3, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.5, 0.3, 0.4, 
    0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.3, _, _, _, _, _, _, _, _, 0.3, 0.3, 0.4, 
    0.4, 0.4, _, _, _, _, 0.5, 0.5, 0.5, 0.4, 0.5, 0.5, 0.4, 0.4, 0.4, 0.5, 
    0.4, 0.3, 0.4, 0.4, 0.5, 0.5, _, 0.4, _,
  0.5, 0.5, 0.6, 1.4, 1.3, 0.9, 0.9, 0.9, 0.8, 0.7, 0.9, 1, 0.9, 0.5, 0.8, 
    1.1, 0.7, 0.6, 0.5, 0.6, 0.6, 0.5, 0.5, 0.5, 0.5, 0.6, 0.5, 0.5, 1, 1, 
    0.8, 0.8, 0.6, 0.7, 0.7, 0.5, _, _, _, _, _, _, _, _, 0.4, 0.4, 0.5, 0.6, 
    0.7, 0.6, 0.6, 0.6, 0.5, _, _, _, 0.5, 0.5, _, 0.7, 0.6, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.4, _, _, _, _, _,
  0.5, 0.6, 0.3, 0.3, 0.4, 0.4, 0.4, 0.4, 0.4, 0.5, 0.7, 0.6, 0.6, 0.7, 0.4, 
    0.4, 0.4, 0.4, 0.4, 0.4, 0.3, 0.3, 0.4, 0.4, 0.4, 0.4, 0.3, 0.5, 0.4, 
    0.5, 0.5, 0.5, 0.6, 0.6, 0.5, 0.5, _, _, _, _, _, _, _, _, 0.5, 0.6, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.4, 0.4, 0.4, 0.5, 0.5, 0.4, 0.5, 0.5, 
    0.5, 0.6, 0.6, 0.6, 0.6, 0.5, 0.5, 0.6, 0.4, _, _,
  0.9, 0.9, 0.7, 1.1, 0.5, 0.5, 0.5, 0.4, 0.4, 0.3, 0.4, 0.4, 0.4, 0.3, 0.3, 
    0.4, 0.3, 0.3, 0.4, 0.4, 0.4, 0.4, 0.5, 0.5, 0.6, 0.4, 0.5, 0.5, 0.4, 
    0.4, 0.5, 0.5, 0.5, 0.5, 0.4, 0.4, _, _, _, _, _, _, _, _, 0.4, 0.4, 0.4, 
    0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.5, 0.6, 0.5, 0.4, _, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.4, 0.4, _, 0.5, _,
  1.2, 1.1, 1.4, 1.2, 1, 0.8, 0.7, 0.5, 0.4, 0.5, 0.7, 0.5, 0.8, 0.7, 0.4, 
    0.9, 0.9, 0.9, 1.2, 0.8, 0.5, 0.5, 0.4, 0.4, 0.4, 0.4, 0.6, 0.8, 0.7, 
    0.6, 0.6, 0.5, 0.5, 0.6, 0.6, 0.7, _, _, _, _, _, _, _, _, 0.7, 0.7, 0.8, 
    0.7, 0.8, 0.9, 0.9, 0.8, 0.7, _, _, _, _, 0.4, 0.7, 0.7, 0.6, 0.6, 0.6, 
    0.7, 0.7, _, _, 0.4, 0.5, 0.6, _, _,
  0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.6, 0.6, 0.7, 0.7, 0.7, 0.7, 0.7, 0.7, 
    0.7, 0.8, 0.8, 0.7, 0.8, 0.8, 0.9, 0.7, _, _, _, _, _, 0.9, _, 0.4, _, _, 
    _, 0.8, 0.8, _, _, _, _, _, _, _, _, 0.9, 1, 1.1, 1.1, 1.1, 1.1, 1, 1, 1, 
    0.9, 0.8, _, _, 0.7, 0.6, 0.8, 0.8, 0.8, 0.8, 0.8, _, 0.7, 0.5, _, _, _, 
    _, 0.4,
  0.7, 0.9, 0.7, 0.5, 0.6, 0.5, 0.6, 0.6, 0.6, 0.5, 0.5, 0.5, 0.4, 0.4, 0.4, 
    0.4, 0.4, 0.3, 0.3, 0.3, 0.3, 0.3, 0.3, 0.3, 0.4, 0.4, 0.3, 0.3, 0.3, 
    0.3, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, _, _, _, _, _, _, _, _, 0.4, 0.4, 0.4, 
    0.4, 0.4, 0.4, 0.4, 0.5, 0.4, 0.5, _, 0.6, 0.5, 0.7, 0.6, 0.5, 0.6, 0.6, 
    0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.5, 0.6,
  1, 0.5, 0.5, 0.4, 0.4, 0.7, 0.5, 0.7, 0.6, 0.4, 0.5, 0.5, 0.3, 0.4, 0.6, 
    0.8, 0.9, 0.9, 0.8, 0.5, 0.4, 0.5, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 0.6, 
    0.6, 0.6, 0.6, 0.6, 0.6, 0.7, 0.7, _, _, _, _, _, _, _, _, 0.7, 0.7, 0.7, 
    0.8, 0.8, 0.8, 0.8, 0.8, 0.8, 0.7, _, 0.6, 0.7, 0.7, 0.8, 0.8, 0.7, 0.7, 
    0.7, 0.6, 0.4, 0.5, 0.6, 0.5, 0.5, 0.5, 0.6, 0.6,
  0.5, 0.5, 0.4, 0.3, 0.2, 0.3, 0.8, 0.8, 0.8, 0.8, 0.7, 0.7, 0.6, 0.5, 0.3, 
    0.3, 0.3, 0.3, 0.3, 0.3, 0.5, _, 0.3, 0.3, 0.3, 0.4, 0.3, 0.3, 0.4, 0.3, 
    0.3, 0.4, 0.5, 0.4, 0.4, 0.4, _, _, _, _, _, _, _, _, 0.4, 0.5, 0.5, 0.4, 
    0.5, 0.6, 0.5, 0.5, 0.5, _, _, _, 0.4, _, _, _, _, 0.4, _, _, 0.3, 0.3, 
    0.4, 0.4, 0.4, _, 0.3, _,
  0.7, 1.6, 1.2, 1, 1, 1, 0.8, 1, 1.2, 1.4, 1.5, 1.4, 1.5, 1.8, 1.2, 0.8, 
    0.5, 0.6, 0.6, 0.7, 0.5, _, _, _, _, _, _, _, 0.5, 0.3, 0.5, _, 0.3, _, 
    _, 0.7, _, _, _, _, _, _, _, _, 0.7, 0.6, 0.5, 0.5, 0.4, _, _, 0.5, 0.7, 
    _, _, _, _, _, 0.5, 0.8, 0.8, 0.8, 0.9, _, _, _, 0.3, _, _, _, _, _,
  1.1, 0.8, 0.9, 0.9, 1, 1.2, 1, 0.8, 0.9, 0.8, 0.4, 0.4, 0.5, 0.6, 0.6, 0.6, 
    0.7, 0.8, 0.5, 0.7, 0.5, 0.5, _, 0.4, 0.5, 0.4, _, _, 0.5, 0.4, 0.4, 0.4, 
    0.4, 0.5, 0.4, _, _, _, _, _, _, _, _, _, _, _, _, _, 0.3, 0.4, 0.4, 0.5, 
    _, _, _, _, _, _, 0.6, _, _, _, _, _, 0.4, _, _, _, _, _, _, _,
  5.6, 0.8, 0.6, 0.6, 0.6, 0.5, 0.5, 0.5, 0.5, 0.6, 0.5, 0.5, 0.6, 0.8, 0.4, 
    0.4, 0.4, 0.4, 0.4, 0.4, 0.3, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 
    0.4, 0.4, 0.4, 0.4, 0.4, 0.4, 0.4, _, _, _, _, _, _, _, _, 0.5, 0.5, 0.5, 
    0.5, 0.5, 0.5, 0.6, 0.6, 0.6, 0.6, 0.5, 0.6, 0.7, 0.7, 0.8, 0.6, 0.6, 
    0.6, 0.6, 0.5, 0.4, 0.5, 0.4, 0.5, 0.5, 0.5, 0.3, 0.3,
  0.5, 0.9, 0.6, 0.4, 0.5, 0.6, 0.5, 0.4, 0.4, 0.4, 0.4, 0.3, 0.3, 0.3, 0.3, 
    0.3, 0.5, 0.7, 0.7, 0.6, 0.5, 0.4, 0.4, 0.4, 0.5, 0.5, 0.5, _, 0.6, 0.6, 
    0.6, 0.6, 0.7, 0.7, 0.7, 0.7, _, _, _, _, _, _, _, _, 0.7, 0.8, 0.8, 0.8, 
    0.8, 0.7, 0.6, 0.5, _, 0.5, 0.6, _, _, _, 0.8, 0.8, 0.8, 0.8, 0.7, 0.7, 
    0.6, 0.7, _, _, _, 0.6, 0.5, 0.4,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 0.5, 1, 0.7, _, 0.8, 0.7, 1, 0.9, 0.9, 0.8, 0.8, 0.7, 0.7, 0.7, 0.8, 
    0.7, 1.1, 1.1, 1, 1.1, 1.2, 1.1, 1.2, 1.7, 1.7, 2.1, 0.8, 1.9, 2, 1.8, 
    1.9, 1.7, 2.1, 2, 1, _, _, _, _, _, _, _, _, 1.6, 1.6, 1.1, 0.9, 0.8, 
    0.8, 0.9, 0.9, _, _, 0.8, 0.8, 0.9, 0.9, 0.8, 0.8, 0.8, 0.7, 0.7, 0.5, 
    0.6, 0.5, 0.5, 0.5, 0.5, _, _, _,
  0.4, 0.5, 0.5, 0.7, 0.5, 0.3, 1, 0.6, 0.7, 1, 1.9, 0.3, 0.3, 1.4, 1.2, 0.8, 
    0.9, 0.8, 0.6, 0.5, 0.6, 0.7, 0.7, 0.8, 0.7, 0.6, 0.5, 0.4, 0.7, 0.6, 
    0.5, 0.6, 0.6, 0.6, 0.5, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.4, 1.2, 1, 0.9, 1, 0.9, 1, 1.6, 1.3, 0.4, 0.4, 0.3, 0.4, 0.4, 0.6, 0.4, 
    0.3, 0.3, 0.3, 0.3, _, _, _, _, _, _, _, _, _, _, _, _, 0.4, 0.4, 0.4, 
    0.5, _, _, _, _, _, _, _, _, 0.4, 0.5, 0.5, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  0.5, 0.5, 0.7, 1, 1, 0.9, 0.7, 0.9, 0.8, 0.8, 0.7, 0.9, 0.5, 0.4, 0.5, 0.6, 
    0.5, 0.6, 0.5, 0.4, 0.4, 0.4, 0.5, 0.5, 0.5, 0.5, 0.4, _, 0.6, 0.7, 0.6, 
    0.6, 0.7, 0.7, 0.7, 0.8, _, _, _, _, _, _, _, _, 0.8, 0.7, 0.8, 0.5, 0.5, 
    _, _, _, _, _, _, _, _, _, _, _, _, 0.8, 0.9, 0.9, 0.8, 0.8, _, _, _, _, 
    0.6, 0.6 ;

 beamNames =
  "North   ",
  "East    ",
  "Vertical" ;

 azimBeam =
  343, 73, 343,
  10, 100, 10,
  344, 74, 344,
  346, 76, 346,
  350, 80, 350,
  355, 85, 355,
  52, 142, 52,
  352, 82, 352,
  344, 74, 344,
  350, 80, 350,
  15, 105, 15,
  348, 78, 348,
  347, 77, 347,
  1, 91, 1,
  0, 90, 0,
  352, 82, 352,
  338, 68, 338,
  0, 90, 0,
  347, 77, 347,
  349, 79, 349,
  354, 84, 354,
  130, 220, 130,
  351, 81, 351,
  341, 71, 341,
  340, 70, 340,
  355, 85, 355 ;

 elevBeam =
  73.7, 73.7, 90,
  73.7, 73.7, 90,
  73.7, 73.7, 90,
  73.7, 73.7, 90,
  73.7, 73.7, 90,
  73.7, 73.7, 90,
  73.7, 73.7, 90,
  73.7, 73.7, 90,
  73.7, 73.7, 90,
  73.7, 73.7, 90,
  73.7, 73.7, 90,
  73.7, 73.7, 90,
  73.7, 73.7, 90,
  73.7, 73.7, 90,
  73.7, 73.7, 90,
  73.7, 73.7, 90,
  73.7, 73.7, 90,
  73.7, 73.7, 90,
  73.7, 73.7, 90,
  73.7, 73.7, 90,
  73.7, 73.7, 90,
  73.7, 73.7, 90,
  73.7, 73.7, 90,
  73.7, 73.7, 90,
  73.7, 73.7, 90,
  73.7, 73.7, 90 ;

 momentsQualityCode =
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  0, 0, 0,
  _, _, _,
  0, 0, 0,
  4, 4, 4,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  8, 8, 8,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  8, 8, 8,
  0, 0, 0,
  _, _, _,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  2, 2, 2,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  4, 4, 4,
  4, 4, 4,
  4, 4, 4,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  4, 4, 4,
  4, 4, 4,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  4, 4, 4,
  4, 4, 4,
  0, 0, 0,
  0, 0, 0,
  4, 4, 4,
  4, 4, 4,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  4, 4, 4,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  0, 0, 0,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  4, 4, 4,
  4, 4, 4,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  8, 8, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  0, 0, 0,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, _,
  _, _, _,
  _, _, _,
  0, 0, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, _,
  0, 0, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  _, _, _,
  8, 8, 8,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  2, 2, 2,
  0, 0, 0,
  4, 4, 4,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  4, 4, 4,
  4, 4, 4,
  4, 4, 4,
  4, 4, 4,
  0, 0, 0,
  4, 4, 4,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  4, 4, 4,
  4, 4, 4,
  4, 4, 4,
  4, 4, 4,
  0, 0, 0,
  4, 4, 4,
  4, 4, 4,
  0, 0, 0,
  8, 8, 8,
  8, 8, 8,
  0, 0, 0,
  0, 0, 0,
  8, 8, 8,
  2, 2, 2,
  8, 8, 8,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  8, 8, 8,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  8, 8, 8,
  2, 2, 2,
  2, 2, 2,
  2, 2, 2,
  2, 2, 2,
  2, 2, _,
  2, 2, _,
  _, _, _,
  2, 2, 2,
  _, _, _,
  _, _, _,
  _, _, _,
  2, 2, _,
  2, 2, 2,
  _, _, _,
  _, _, _,
  2, 2, 2,
  2, 2, 2,
  2, 2, 2,
  2, 2, 2,
  2, 2, 2,
  _, _, _,
  2, 2, 2,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  4, 4, 4,
  4, 4, 4,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  8, 8, 8,
  8, 8, 8,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  8, 8, 8,
  0, 0, 0,
  0, 0, 0,
  0, 0, _,
  0, 0, 0,
  0, 0, _,
  0, 0, _,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  0, 0, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, _,
  0, 0, _,
  0, 0, _,
  0, 0, 0,
  0, 0, _,
  _, _, _,
  _, _, _,
  0, 0, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  8, 8, _,
  0, 0, 0,
  0, 0, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  8, 8, 8,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  4, 4, 4,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  4, 4, 4,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, _,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  8, 8, 8,
  4, 4, 4,
  4, 4, 4,
  _, _, _,
  0, 0, 0,
  4, 4, 4,
  4, 4, 4,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  8, 8, 8,
  8, 8, 8,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  2, 2, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  2, 2, _,
  4, 4, 4,
  4, 4, 4,
  4, 4, 4,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  4, 4, 4,
  4, 4, 4,
  8, 8, 8,
  8, 8, 8,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  8, 8, _,
  0, 0, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0, 0, _,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  0, 0, 0,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  2, 2, 2,
  2, 2, 2 ;

 consensusNum =
  910, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 
    1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 
    1010, 1010, 1010, 1010, 909, 909, 909, 910, 910, 710, 710, 810, _, _, _, 
    _, _, _, _, _, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1009, 
    1010, 1010, 910, 910, 809, 909, 910, 1010, 910, 1010, 910, 1010, 910, 
    910, 709, _, _, 506, _,
  404, 505, _, 409, 809, _, _, 705, 709, 408, _, _, 409, 709, 609, 709, 709, 
    509, 809, 409, 808, 809, 807, 808, 707, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  809, 809, 809, 809, 809, 809, 809, 809, 809, 809, 809, 809, 709, 809, 809, 
    809, 809, 809, 809, 709, 609, 709, 709, 808, 604, 504, 605, 807, 810, 
    810, 810, 810, 810, 505, 808, 404, _, _, _, _, _, _, _, _, 810, 810, 810, 
    409, _, _, _, 406, 404, _, _, _, _, _, _, _, 405, 404, 506, 605, 405, _, 
    _, _, _, _, _, _,
  1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 
    910, 1010, 1010, 610, 810, _, 810, _, _, _, _, _, _, 609, _, _, 710, 410, 
    510, 610, 510, 510, 710, 810, _, _, _, _, _, _, _, _, 810, 610, 510, _, 
    _, 510, 810, 910, 810, 910, 710, 506, _, _, _, _, _, _, _, 410, _, _, _, 
    _, _, _, _, _,
  909, 909, 709, 909, 1009, 909, 1009, 1009, 1009, 909, 809, 709, 809, 808, 
    907, 807, 807, 907, 807, 908, 1008, 1009, 1008, 809, 909, 909, 809, 909, 
    1009, 1009, 1009, 1009, 909, 1009, 1009, 1009, _, _, _, _, _, _, _, _, 
    1009, 1009, 909, 909, 909, 909, 909, 909, 909, 909, 1009, 909, 909, 1008, 
    1009, 1009, 1009, 1009, 1009, 1009, 909, 1009, 1009, 1009, 1009, 1008, 
    604, _,
  710, 610, 810, 910, 810, 1010, 910, 710, 910, 1010, 1010, 1010, 909, 1010, 
    1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 907, 1010, 
    910, _, 1010, 910, 810, 910, 404, 405, 607, 405, _, _, _, _, _, _, _, _, 
    809, 809, 809, 808, 808, 909, 709, 506, 504, _, 504, 608, 708, 809, 507, 
    506, 406, 404, _, _, _, _, _, _, _, _, _, _,
  _, _, 710, 909, 908, 1010, 1010, 910, 1010, 1010, 1009, 907, 907, 1008, 
    908, 908, 1010, 1010, 1010, 909, 1010, 1009, 1009, 909, 607, 604, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  910, 709, 1009, 1010, 910, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 
    1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 
    1010, 1010, 1010, 1010, 1010, 910, 910, 1010, 1010, 810, 708, _, _, _, _, 
    _, _, _, _, 1010, 1010, 1010, 1010, 1010, 1010, 1009, 1009, 909, 1009, 
    1009, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 
    1010, 1010, 1010, 1010, 809, 606,
  910, 810, 810, 610, 710, 1010, 1010, 1010, 1010, 1010, 1009, 1010, 1010, 
    1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 
    908, 809, 605, 907, 605, 1010, 908, 1010, 808, 908, 504, _, _, _, _, _, 
    _, _, _, 1010, 1010, 1010, 1010, 809, _, _, _, _, 406, 607, 808, 1009, 
    809, 808, 909, 908, 910, 1008, 908, 909, 1009, 608, 407, 605, _, 506, _,
  1005, 1010, 1010, 810, 910, 710, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 
    1010, 810, 1010, 1010, 909, 1010, 1010, 910, 1008, 1010, 909, 910, 1010, 
    1010, 1010, 1010, 910, 1010, 1010, 1010, 806, 708, 505, _, _, _, _, _, _, 
    _, _, 1010, 1010, 809, 808, 807, 1006, 906, 806, 405, _, _, _, 504, 406, 
    _, 806, 909, 1009, 810, 709, 508, 407, 404, _, _, _, _, _,
  1009, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 
    1010, 1010, 1009, 1010, 1010, 1010, 1008, 907, 608, 1009, 1010, 1010, 
    1010, 1010, 907, 804, 704, 506, 406, 1010, 910, 910, 810, 810, _, _, _, 
    _, _, _, _, _, 609, 807, 908, 810, 1009, 1009, 1009, 1009, 807, 905, 807, 
    908, 1008, 1009, 909, 909, 909, 910, 910, 910, 1010, 910, 1009, 907, 907, 
    707, _, _,
  910, 1009, 1009, 1010, 910, 1010, 1010, 1010, 910, 1010, 1010, 1010, 910, 
    1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 808, 
    1010, 910, 910, 1010, 910, 910, 910, 406, 910, 910, 909, _, _, _, _, _, 
    _, _, _, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 909, 506, 
    507, 405, 405, _, 806, 1008, 1008, 908, 909, 909, 910, 809, 606, 506, _, 
    508, _,
  910, 910, 1008, 1008, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 
    1010, 1010, 1010, 1010, 1010, 1009, 1007, 1010, 1006, 1009, 1010, 1010, 
    1010, 1010, 1009, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1008, _, _, 
    _, _, _, _, _, _, 1010, 1010, 1010, 1010, 1010, 909, 909, 808, 605, _, _, 
    _, _, 804, 1005, 1006, 1008, 1008, 1008, 806, 504, _, _, 904, 805, 604, 
    _, _,
  710, 910, 910, 1010, 1009, 909, 909, 910, 1010, 1010, 1010, 1010, 1010, 
    1010, 1010, 610, 910, 710, 809, 910, 910, 710, 408, _, _, _, _, _, 609, 
    _, 405, _, _, _, 608, 708, _, _, _, _, _, _, _, _, 807, 1010, 1010, 1010, 
    1010, 1010, 1010, 910, 710, 710, 410, _, _, 406, 408, 509, 809, 910, 809, 
    708, _, 406, 407, _, _, _, _, 407,
  910, 810, 910, 910, 910, 910, 810, 910, 910, 910, 910, 910, 910, 910, 910, 
    910, 910, 910, 910, 910, 910, 910, 910, 910, 910, 910, 910, 910, 910, 
    609, 508, 506, 910, 606, 809, 910, _, _, _, _, _, _, _, _, 910, 910, 910, 
    910, 910, 910, 910, 910, 810, 709, _, 508, 708, 810, 810, 910, 910, 910, 
    910, 910, 810, 810, 910, 810, 910, 910, 810, 810,
  710, 610, 910, 1010, 910, 808, 909, 1010, 1010, 1010, 1010, 910, 1010, 910, 
    1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 910, 
    910, 910, 1010, 1010, 1009, 909, 706, 704, 910, 909, _, _, _, _, _, _, _, 
    _, 909, 909, 909, 1009, 1009, 1009, 809, 809, 609, 408, _, 407, 609, 909, 
    1009, 909, 909, 709, 508, 506, 406, 405, 404, 506, 507, 608, 808, 1010,
  1010, 1010, 1009, 1010, 1010, 910, 1010, 1010, 1010, 910, 1010, 810, 410, 
    1010, 1010, 810, 910, 1010, 810, 710, 609, _, 909, 1010, 1010, 610, 409, 
    710, 709, 710, 410, 910, 1010, 910, 810, 910, _, _, _, _, _, _, _, _, 
    710, 710, 509, 408, 505, 606, 707, 707, 704, _, _, _, 406, _, _, _, _, 
    406, _, _, 405, 706, 910, 609, 510, _, 607, _,
  610, 408, 409, 809, 810, 808, 806, 907, 1009, 1010, 1010, 910, 909, 907, 
    909, 710, 410, 810, 809, 509, 509, _, _, _, _, _, _, _, 508, 504, 505, _, 
    505, _, _, 506, _, _, _, _, _, _, _, _, 706, 808, 807, 704, 404, _, _, 
    604, 504, _, _, _, _, _, 607, 806, 909, 807, 504, _, _, _, 504, _, _, _, 
    _, _,
  708, 809, 909, 909, 909, 909, 909, 809, 909, 708, 809, 809, 808, 809, 809, 
    909, 809, 909, 909, 909, 708, 608, _, 809, 809, 808, _, _, 604, 807, 909, 
    504, 809, 508, 406, _, _, _, _, _, _, _, _, _, _, _, _, _, 404, 505, 407, 
    404, _, _, _, _, _, _, 504, _, _, _, _, _, 404, _, _, _, _, _, _, _,
  1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 
    1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 
    1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 910, 1010, 1008, 1009, _, 
    _, _, _, _, _, _, _, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 
    1010, 910, 810, 809, 1010, 1010, 1010, 710, 1010, 1010, 1010, 909, 907, 
    806, 808, 908, 808, 806, 806, 704,
  710, 810, 810, 510, 810, 910, 910, 1010, 1010, 1010, 1010, 1010, 1010, 
    1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 910, 
    910, 810, _, 910, 610, 506, 505, 405, 707, 808, 607, _, _, _, _, _, _, _, 
    _, 1010, 1010, 1010, 1010, 910, 909, 909, 707, _, 606, 506, _, _, _, 506, 
    807, 909, 910, 1010, 910, 710, 409, _, _, _, 506, 506, 505,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  _, 910, 810, 508, _, 407, 508, 609, 608, 708, 708, 608, 708, 608, 708, 709, 
    809, 809, 509, 607, 506, 605, 706, 606, 505, 705, 707, 607, 608, 707, 
    606, 408, 608, 604, 407, 406, _, _, _, _, _, _, _, _, 406, 507, 508, 409, 
    510, 709, 608, 507, _, _, 406, 407, 608, 610, 610, 610, 709, 508, 608, 
    408, 508, 608, 608, 608, 407, _, _, _,
  910, 910, 1010, 1010, 709, 707, 1010, 1010, 1010, 1010, 907, 806, 705, 806, 
    908, 1008, 1009, 1010, 1010, 1010, 1010, 1010, 1009, 1010, 1010, 1010, 
    809, 604, 910, 705, 706, 1010, 1009, 906, 604, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  1010, 1010, 1010, 1010, 1010, 1010, 1010, 910, 810, 610, 610, 710, 1010, 
    1010, 1010, 810, 810, 910, 410, 410, _, _, _, _, _, _, _, _, _, _, 410, 
    410, 504, 706, 704, 606, _, _, _, _, _, _, _, _, 608, 608, 405, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _,
  909, 1010, 1010, 1010, 1010, 1010, 1010, 1010, 910, 910, 1010, 1010, 1010, 
    1010, 1010, 1010, 810, 910, 1010, 910, 1009, 1010, 1010, 1009, 806, 910, 
    710, _, 1010, 1010, 1010, 910, 1010, 1010, 1010, 709, _, _, _, _, _, _, 
    _, _, 1010, 1010, 807, 505, 404, _, _, _, _, _, _, _, _, _, _, _, _, 606, 
    707, 707, 608, 607, _, _, _, _, 504, 405 ;

 consensusNumBeam =
  10, 9, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 9, 9,
  9, 9, 9,
  10, 9, 9,
  9, 10, 10,
  9, 10, 10,
  7, 8, 10,
  9, 7, 10,
  9, 8, 10,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 9,
  10, 10, 10,
  10, 10, 10,
  10, 9, 10,
  9, 9, 10,
  8, 9, 9,
  9, 9, 9,
  9, 9, 10,
  10, 10, 10,
  9, 10, 10,
  10, 10, 10,
  9, 10, 10,
  10, 10, 10,
  10, 9, 10,
  9, 9, 10,
  7, 7, 9,
  _, 5, 4,
  _, 6, 4,
  5, 6, 6,
  _, 5, 6,
  4, 6, 4,
  9, 5, 5,
  5, _, 8,
  9, 4, 9,
  8, 8, 9,
  8, 6, _,
  6, 5, _,
  8, 7, 5,
  7, 7, 9,
  4, 4, 8,
  _, _, 9,
  _, 5, 9,
  4, 8, 9,
  7, 8, 9,
  6, 6, 9,
  9, 7, 9,
  9, 7, 9,
  8, 5, 9,
  9, 8, 9,
  9, 4, 9,
  8, 8, 8,
  9, 8, 9,
  9, 8, 7,
  8, 9, 8,
  9, 7, 7,
  _, _, _,
  _, _, _,
  _, _, _,
  _, 8, 9,
  _, 8, 9,
  _, 9, 9,
  _, 8, 9,
  _, 4, 9,
  _, 4, 9,
  _, _, 8,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, 6,
  _, _, 8,
  _, _, 8,
  _, _, 8,
  _, _, 6,
  _, _, _,
  _, _, 4,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, 4,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, 5,
  _, _, 8,
  _, 4, 9,
  _, _, 9,
  _, _, 9,
  _, _, 9,
  9, 8, 9,
  9, 8, 9,
  9, 8, 9,
  9, 8, 9,
  9, 8, 9,
  9, 8, 9,
  9, 8, 9,
  9, 8, 9,
  9, 8, 9,
  8, 8, 9,
  9, 8, 9,
  9, 8, 9,
  7, 8, 9,
  9, 8, 9,
  9, 8, 9,
  9, 8, 9,
  9, 8, 9,
  9, 8, 9,
  9, 8, 9,
  9, 7, 9,
  9, 6, 9,
  9, 7, 9,
  8, 7, 9,
  8, 8, 8,
  6, 8, 4,
  5, 6, 4,
  6, 7, 5,
  9, 8, 7,
  9, 8, 10,
  9, 8, 10,
  9, 8, 10,
  9, 8, 10,
  9, 8, 10,
  5, 7, 5,
  8, 8, 8,
  6, 4, 4,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  9, 8, 10,
  9, 8, 10,
  8, 8, 10,
  4, 8, 9,
  _, 4, 6,
  _, 5, 6,
  _, 6, 6,
  5, 4, 6,
  4, 4, 4,
  _, _, 4,
  _, _, 4,
  4, _, _,
  _, _, 5,
  _, 5, 5,
  _, 5, _,
  _, 5, 5,
  5, 4, 5,
  6, 4, 4,
  7, 5, 6,
  7, 6, 5,
  4, 6, 5,
  _, 4, 5,
  _, _, 6,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, 4,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 9, 10,
  10, 10, 10,
  10, 10, 10,
  10, 6, 10,
  10, 8, 10,
  10, _, 10,
  10, 8, 10,
  8, _, 9,
  6, _, 5,
  _, _, _,
  _, _, _,
  _, _, _,
  7, _, 8,
  10, 6, 9,
  10, _, 9,
  10, _, 9,
  10, 7, 10,
  10, 4, 10,
  10, 5, 10,
  10, 6, 10,
  10, 5, 10,
  10, 5, 10,
  10, 7, 10,
  9, 8, 10,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  10, 8, 10,
  10, 6, 10,
  10, 5, 10,
  10, _, 10,
  9, _, 10,
  9, 5, 10,
  9, 8, 10,
  9, 9, 10,
  9, 8, 10,
  9, 9, 10,
  9, 7, 10,
  9, 5, 6,
  6, _, _,
  6, _, 4,
  6, _, 6,
  6, _, 6,
  4, _, 7,
  5, _, 6,
  6, _, 9,
  7, 4, 10,
  8, _, 10,
  7, _, 10,
  8, _, 10,
  7, _, 9,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  9, 10, 9,
  10, 9, 9,
  7, 10, 9,
  10, 9, 9,
  10, 10, 9,
  9, 10, 9,
  10, 10, 9,
  10, 10, 9,
  10, 10, 9,
  9, 10, 9,
  8, 10, 9,
  7, 10, 9,
  8, 10, 9,
  8, 10, 8,
  9, 10, 7,
  8, 10, 7,
  9, 8, 7,
  9, 9, 7,
  10, 8, 7,
  10, 9, 8,
  10, 10, 8,
  10, 10, 9,
  10, 10, 8,
  8, 10, 9,
  9, 9, 9,
  9, 9, 9,
  8, 9, 9,
  9, 10, 9,
  10, 10, 9,
  10, 10, 9,
  10, 10, 9,
  10, 10, 9,
  9, 10, 9,
  10, 10, 9,
  10, 10, 9,
  10, 10, 9,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  10, 10, 9,
  10, 10, 9,
  10, 9, 9,
  10, 9, 9,
  10, 9, 9,
  10, 9, 9,
  10, 9, 9,
  10, 9, 9,
  10, 9, 9,
  10, 9, 9,
  10, 10, 9,
  10, 9, 9,
  10, 9, 9,
  10, 10, 8,
  10, 10, 9,
  10, 10, 9,
  10, 10, 9,
  10, 10, 9,
  10, 10, 9,
  10, 10, 9,
  10, 9, 9,
  10, 10, 9,
  10, 10, 9,
  10, 10, 9,
  10, 10, 9,
  10, 10, 8,
  6, 7, 4,
  _, 7, 6,
  7, 9, 10,
  7, 6, 10,
  8, 9, 10,
  9, 10, 10,
  8, 10, 10,
  10, 10, 10,
  9, 10, 10,
  7, 10, 10,
  9, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  9, 10, 9,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  9, 9, 7,
  10, 10, 10,
  9, 10, 10,
  4, 5, _,
  10, 10, 10,
  10, 9, 10,
  8, 9, 10,
  9, 10, 10,
  4, 8, 4,
  4, 9, 5,
  6, 9, 7,
  4, 8, 5,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  8, 10, 9,
  8, 10, 9,
  8, 10, 9,
  8, 10, 8,
  8, 10, 8,
  9, 9, 9,
  7, 9, 9,
  5, 8, 6,
  5, 8, 4,
  _, 6, _,
  6, 5, 4,
  8, 6, 8,
  7, 8, 8,
  8, 9, 9,
  5, 9, 7,
  5, 7, 6,
  4, 8, 6,
  4, 8, 4,
  _, 6, _,
  _, 6, _,
  _, _, 4,
  _, _, 4,
  _, _, _,
  _, _, _,
  _, _, _,
  4, _, _,
  6, _, _,
  _, 4, 4,
  _, _, 10,
  _, 4, _,
  8, 7, 10,
  9, 10, 9,
  9, 10, 8,
  10, 10, 10,
  10, 10, 10,
  9, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 9,
  10, 9, 7,
  10, 9, 7,
  10, 10, 8,
  9, 10, 8,
  10, 9, 8,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 9, 9,
  10, 10, 10,
  10, 10, 9,
  10, 10, 9,
  10, 9, 9,
  6, 6, 7,
  7, 6, 4,
  4, _, _,
  _, _, _,
  4, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  9, 10, 10,
  7, 9, 9,
  10, 10, 9,
  10, 10, 10,
  10, 9, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 9, 10,
  10, 9, 10,
  10, 10, 10,
  10, 10, 10,
  9, 8, 10,
  8, 7, 8,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 9,
  10, 10, 9,
  10, 9, 9,
  10, 10, 9,
  10, 10, 9,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 8, 9,
  6, 9, 6,
  9, 10, 10,
  8, 10, 10,
  8, 9, 10,
  6, 9, 10,
  7, 9, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 9,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 9, 8,
  8, 10, 9,
  6, 8, 5,
  9, 9, 7,
  7, 6, 5,
  10, 10, 10,
  9, 10, 8,
  10, 10, 10,
  9, 8, 8,
  10, 9, 8,
  5, 7, 4,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  8, 10, 9,
  _, 10, 7,
  _, 8, 4,
  _, 7, 5,
  _, 7, 5,
  4, 9, 6,
  6, 10, 7,
  8, 10, 8,
  10, 10, 9,
  8, 10, 9,
  8, 10, 8,
  10, 9, 9,
  10, 9, 8,
  9, 10, 10,
  10, 10, 8,
  9, 10, 8,
  9, 10, 9,
  10, 10, 9,
  6, 8, 8,
  4, 7, 7,
  6, 7, 5,
  _, _, 7,
  5, 9, 6,
  _, 8, 5,
  10, 10, 5,
  10, 10, 10,
  10, 10, 10,
  10, 8, 10,
  10, 9, 10,
  10, 7, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 8, 10,
  10, 10, 10,
  10, 10, 10,
  10, 9, 9,
  10, 10, 10,
  10, 10, 10,
  10, 9, 10,
  10, 10, 8,
  10, 10, 10,
  10, 9, 9,
  10, 9, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 9, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 8, 6,
  8, 7, 8,
  7, 5, 5,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  10, 10, 10,
  10, 10, 10,
  10, 8, 9,
  10, 8, 8,
  10, 8, 7,
  10, 10, 6,
  10, 9, 6,
  9, 8, 6,
  6, 4, 5,
  _, _, _,
  5, _, _,
  6, 4, _,
  7, 5, 4,
  8, 4, 6,
  8, 6, _,
  10, 8, 6,
  10, 9, 9,
  10, 10, 9,
  10, 8, 10,
  8, 7, 9,
  10, 5, 8,
  9, 4, 7,
  6, 4, 4,
  4, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  10, 10, 9,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 9,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 8,
  9, 10, 7,
  6, 10, 8,
  10, 10, 9,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 9, 7,
  8, 8, 4,
  8, 7, 4,
  6, 5, 6,
  4, 6, 6,
  10, 10, 10,
  10, 9, 10,
  10, 9, 10,
  8, 8, 10,
  8, 8, 10,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  6, 10, 9,
  8, 10, 7,
  9, 10, 8,
  8, 10, 10,
  10, 10, 9,
  10, 10, 9,
  10, 10, 9,
  10, 10, 9,
  9, 8, 7,
  9, 9, 5,
  8, 9, 7,
  9, 10, 8,
  10, 10, 8,
  10, 10, 9,
  10, 9, 9,
  10, 9, 9,
  10, 9, 9,
  10, 9, 10,
  10, 9, 10,
  10, 9, 10,
  10, 10, 10,
  10, 9, 10,
  10, 10, 9,
  9, 9, 7,
  9, 9, 7,
  7, 9, 7,
  4, _, 5,
  _, _, 4,
  10, 9, 10,
  10, 10, 9,
  10, 10, 9,
  10, 10, 10,
  9, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 9, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 9, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 8, 8,
  10, 10, 10,
  10, 9, 10,
  9, 10, 10,
  10, 10, 10,
  10, 9, 10,
  9, 9, 10,
  9, 9, 10,
  7, 4, 6,
  9, 9, 10,
  9, 9, 10,
  10, 9, 9,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  9, 9, 9,
  5, 7, 6,
  5, 6, 7,
  5, 4, 5,
  5, 4, 5,
  4, 6, _,
  8, 10, 6,
  10, 10, 8,
  10, 10, 8,
  9, 10, 8,
  9, 10, 9,
  9, 10, 9,
  9, 10, 10,
  8, 9, 9,
  8, 6, 6,
  6, 5, 6,
  6, _, 7,
  5, 5, 8,
  _, 5, 6,
  9, 10, 10,
  9, 10, 10,
  10, 10, 8,
  10, 10, 8,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 9,
  10, 10, 7,
  10, 10, 10,
  10, 10, 6,
  10, 10, 9,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 9,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 8,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  9, 10, 9,
  9, 10, 9,
  8, 10, 8,
  6, 10, 5,
  4, 7, _,
  _, 5, 4,
  _, 5, _,
  6, 7, _,
  8, 9, 4,
  10, 10, 5,
  10, 10, 6,
  10, 10, 8,
  10, 10, 8,
  10, 10, 8,
  8, 10, 6,
  5, 10, 4,
  4, 7, _,
  7, 9, _,
  9, 10, 4,
  8, 9, 5,
  8, 6, 4,
  5, 8, _,
  _, 10, _,
  10, 7, 10,
  10, 9, 10,
  9, 9, 10,
  10, 10, 10,
  10, 10, 9,
  9, 10, 9,
  10, 9, 9,
  10, 9, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 6, 10,
  10, 9, 10,
  10, 7, 10,
  10, 8, 9,
  10, 9, 10,
  10, 9, 10,
  10, 7, 10,
  9, 4, 8,
  8, _, 7,
  7, _, 5,
  5, _, 5,
  _, _, 4,
  _, _, _,
  9, 6, 9,
  9, _, 8,
  4, 4, 5,
  9, _, 9,
  4, _, 4,
  10, _, 9,
  10, 6, 8,
  10, 7, 8,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  10, 8, 7,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 9, 10,
  10, 7, 10,
  10, 7, 10,
  10, 4, 10,
  9, _, 9,
  8, _, 6,
  8, 4, 6,
  10, 4, 8,
  10, 5, 9,
  10, 8, 9,
  10, 9, 10,
  10, 8, 9,
  10, 7, 8,
  5, _, 7,
  9, 4, 6,
  6, 4, 7,
  4, _, 7,
  4, _, 5,
  _, _, 5,
  _, _, 6,
  4, 4, 7,
  9, 9, 10,
  9, 8, 10,
  9, 9, 10,
  9, 9, 10,
  9, 9, 10,
  9, 9, 10,
  9, 8, 10,
  9, 9, 10,
  9, 9, 10,
  9, 9, 10,
  9, 9, 10,
  9, 9, 10,
  9, 9, 10,
  9, 9, 10,
  9, 9, 10,
  9, 9, 10,
  9, 9, 10,
  9, 9, 10,
  9, 9, 10,
  9, 9, 10,
  9, 9, 10,
  9, 9, 10,
  9, 9, 10,
  9, 9, 10,
  9, 9, 10,
  9, 9, 10,
  9, 9, 10,
  9, 9, 10,
  9, 9, 10,
  8, 6, 9,
  7, 5, 8,
  5, 5, 6,
  9, 9, 10,
  6, 8, 6,
  9, 8, 9,
  9, 9, 10,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  9, 9, 10,
  9, 9, 10,
  9, 9, 10,
  9, 9, 10,
  9, 9, 10,
  9, 9, 10,
  9, 9, 10,
  9, 9, 10,
  9, 8, 10,
  9, 7, 9,
  7, _, 8,
  7, 5, 8,
  7, 7, 8,
  8, 8, 10,
  8, 9, 10,
  9, 9, 10,
  9, 9, 10,
  9, 9, 10,
  9, 9, 10,
  9, 9, 10,
  9, 8, 10,
  9, 8, 10,
  9, 9, 10,
  9, 8, 10,
  9, 9, 10,
  9, 9, 10,
  9, 8, 10,
  9, 8, 10,
  7, 10, 10,
  6, 8, 10,
  9, 9, 10,
  10, 10, 10,
  10, 9, 10,
  9, 8, 8,
  9, 10, 9,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 9, 10,
  10, 10, 10,
  9, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  9, 10, 10,
  9, 10, 10,
  9, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 9,
  9, 10, 9,
  7, 10, 6,
  7, 10, 4,
  9, 10, 10,
  9, 10, 9,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  9, 10, 9,
  9, 10, 9,
  9, 10, 9,
  10, 10, 9,
  10, 10, 9,
  10, 10, 9,
  8, 10, 9,
  8, 10, 9,
  6, 10, 9,
  6, 4, 8,
  5, _, 7,
  5, 4, 7,
  6, 8, 9,
  9, 10, 9,
  10, 10, 9,
  9, 10, 9,
  9, 10, 9,
  7, 10, 9,
  5, 10, 8,
  5, 8, 6,
  4, 9, 6,
  4, 9, 5,
  4, 9, 4,
  5, 10, 6,
  5, 10, 7,
  6, 10, 8,
  8, 10, 8,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 9,
  10, 10, 10,
  10, 10, 10,
  9, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 9, 10,
  10, 10, 10,
  10, 8, 10,
  10, 4, 10,
  10, 10, 10,
  10, 10, 10,
  10, 8, 10,
  10, 9, 10,
  10, 10, 10,
  10, 8, 10,
  10, 7, 10,
  10, 6, 9,
  10, _, 4,
  10, 9, 9,
  10, 10, 10,
  10, 10, 10,
  10, 6, 10,
  10, 4, 9,
  10, 7, 10,
  10, 7, 9,
  10, 7, 10,
  10, 4, 10,
  10, 9, 10,
  10, 10, 10,
  10, 9, 10,
  10, 8, 10,
  10, 9, 10,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  10, 7, 10,
  10, 7, 10,
  9, 5, 9,
  8, 4, 8,
  9, 5, 5,
  9, 6, 6,
  10, 7, 7,
  9, 7, 7,
  8, 7, 4,
  4, 6, _,
  4, 10, _,
  _, 8, _,
  4, 6, 6,
  _, 9, 6,
  _, 8, 4,
  _, 8, 4,
  4, 10, _,
  4, 8, 6,
  _, 7, 6,
  _, 8, 5,
  4, 8, 5,
  7, 10, 6,
  9, 9, 10,
  10, 6, 9,
  9, 5, 10,
  6, _, 8,
  8, 6, 7,
  7, _, 8,
  6, 8, 10,
  4, 7, 8,
  4, 6, 9,
  9, 8, 9,
  9, 8, 10,
  8, 8, 8,
  9, 8, 6,
  10, 9, 7,
  10, 10, 9,
  10, 10, 10,
  10, 10, 10,
  9, 9, 10,
  10, 9, 9,
  9, 9, 7,
  9, 9, 9,
  7, 9, 10,
  4, 9, 10,
  8, 9, 10,
  8, 10, 9,
  5, 9, 9,
  5, 9, 9,
  _, 9, 8,
  _, 7, _,
  _, _, _,
  4, _, _,
  4, _, _,
  _, 5, _,
  _, _, _,
  5, 7, 8,
  5, 7, 4,
  5, 7, 5,
  5, 6, _,
  5, 5, 5,
  4, 6, _,
  5, 7, _,
  5, 8, 6,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  7, 9, 6,
  8, 9, 8,
  8, 9, 7,
  7, 8, 4,
  4, 6, 4,
  _, 4, _,
  4, 5, _,
  6, 7, 4,
  5, 8, 4,
  5, 8, _,
  _, 8, _,
  _, 7, _,
  _, 6, _,
  _, 7, _,
  6, 6, 7,
  8, 8, 6,
  9, 9, 9,
  8, 9, 7,
  5, 7, 4,
  5, 5, _,
  5, 4, _,
  6, 5, _,
  5, 7, 4,
  4, 4, _,
  _, 5, _,
  _, _, _,
  4, 5, _,
  _, 5, _,
  7, 7, 8,
  8, 8, 9,
  9, 9, 9,
  9, 9, 9,
  9, 9, 9,
  9, 9, 9,
  9, 9, 9,
  8, 9, 9,
  9, 9, 9,
  9, 7, 8,
  8, 8, 9,
  9, 8, 9,
  9, 8, 8,
  9, 8, 9,
  8, 9, 9,
  9, 9, 9,
  8, 9, 9,
  9, 9, 9,
  9, 9, 9,
  9, 9, 9,
  7, 9, 8,
  7, 6, 8,
  6, _, 6,
  9, 8, 9,
  9, 8, 9,
  8, 8, 8,
  4, _, 5,
  _, _, _,
  6, 8, 4,
  9, 8, 7,
  9, 9, 9,
  5, 5, 4,
  8, 9, 9,
  5, 9, 8,
  4, 7, 6,
  4, 8, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, 7, 4,
  _, _, _,
  _, 4, _,
  _, 4, _,
  4, 6, 4,
  5, 5, 5,
  6, 4, 7,
  4, 5, 4,
  _, _, 4,
  _, _, _,
  _, _, _,
  4, _, _,
  4, _, _,
  4, 5, _,
  5, 7, 4,
  5, 6, _,
  _, 8, 4,
  _, 7, _,
  _, 4, 4,
  _, 4, 6,
  4, 4, 4,
  _, _, 6,
  _, 4, _,
  _, _, _,
  4, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  9, 10, 10,
  10, 10, 10,
  10, 10, 8,
  10, 10, 9,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  9, 9, 10,
  9, 8, 10,
  10, 8, 9,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 7, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 9, 9,
  10, 9, 7,
  10, 8, 6,
  9, 8, 8,
  9, 10, 8,
  8, 10, 8,
  8, 10, 6,
  8, 10, 6,
  7, 8, 4,
  9, 7, 10,
  8, 9, 10,
  9, 8, 10,
  5, 9, 10,
  8, 10, 10,
  9, 10, 10,
  9, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  9, 10, 10,
  9, 10, 10,
  8, 9, 10,
  _, _, _,
  9, 10, 10,
  6, 10, 10,
  5, 6, 6,
  5, 5, 5,
  4, 5, 5,
  8, 7, 7,
  9, 8, 8,
  8, 6, 7,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 9, 10,
  9, 9, 9,
  9, 10, 9,
  7, 8, 7,
  6, 7, _,
  6, 6, 6,
  6, 5, 6,
  6, _, 5,
  6, _, 5,
  6, _, 5,
  6, 5, 6,
  9, 8, 7,
  9, 9, 9,
  9, 9, 10,
  10, 10, 10,
  10, 9, 10,
  10, 7, 10,
  10, 4, 9,
  6, 5, _,
  5, _, _,
  7, _, 6,
  5, 6, 6,
  6, 5, 6,
  5, 5, 5,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  10, _, 10,
  10, 9, 10,
  9, 8, 10,
  6, 5, 8,
  4, _, 7,
  4, 4, 7,
  5, 5, 8,
  6, 6, 9,
  6, 6, 8,
  7, 7, 8,
  7, 7, 8,
  6, 8, 8,
  7, 7, 8,
  8, 6, 8,
  8, 7, 8,
  8, 7, 9,
  8, 8, 9,
  8, 8, 9,
  8, 5, 9,
  8, 6, 7,
  5, 5, 6,
  6, 9, 5,
  7, 8, 6,
  6, 9, 6,
  5, 10, 5,
  7, 9, 5,
  7, 7, 7,
  6, 8, 7,
  6, 8, 8,
  7, 7, 7,
  6, 6, 6,
  4, 7, 8,
  6, 7, 8,
  6, 6, 4,
  4, 4, 7,
  4, 5, 6,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  4, 5, 6,
  5, 5, 7,
  6, 5, 8,
  8, 4, 9,
  9, 5, 10,
  8, 7, 9,
  7, 6, 8,
  7, 5, 7,
  6, _, 6,
  6, _, 6,
  5, 4, 6,
  8, 4, 7,
  8, 6, 8,
  8, 6, 10,
  7, 6, 10,
  7, 6, 10,
  7, 7, 9,
  7, 5, 8,
  6, 6, 8,
  6, 4, 8,
  6, 5, 8,
  7, 6, 8,
  8, 6, 8,
  7, 6, 8,
  6, 4, 7,
  _, 4, 7,
  5, _, 6,
  4, _, _,
  9, 10, 10,
  9, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 7, 9,
  8, 7, 7,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 9, 7,
  8, 8, 6,
  7, 8, 5,
  8, 8, 6,
  10, 9, 8,
  10, 10, 8,
  10, 10, 9,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 9,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  8, 9, 9,
  7, 6, 4,
  9, 10, 10,
  7, 8, 5,
  7, 9, 6,
  10, 10, 10,
  10, 10, 9,
  9, 9, 6,
  6, 7, 4,
  4, 5, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, 4,
  _, 4, 4,
  _, _, 4,
  _, 4, 4,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, 4, _,
  _, _, _,
  _, _, _,
  _, _, 4,
  _, _, _,
  _, _, _,
  _, 4, _,
  _, 6, _,
  5, 5, _,
  7, _, _,
  4, _, _,
  5, _, _,
  _, _, _,
  _, _, _,
  5, _, _,
  4, _, _,
  4, _, _,
  4, 4, _,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  9, 10, 10,
  8, 10, 10,
  6, 6, 10,
  6, 6, 10,
  7, 8, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 8, 10,
  10, 8, 10,
  9, 9, 10,
  4, 4, 10,
  4, 6, 10,
  4, _, 10,
  _, _, 10,
  _, _, 10,
  _, 4, 10,
  _, _, 10,
  _, _, 10,
  _, _, 9,
  _, _, 9,
  _, _, 10,
  _, _, 10,
  4, 4, 10,
  9, 4, 10,
  8, 5, 4,
  9, 7, 6,
  10, 7, 4,
  10, 6, 6,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  10, 6, 8,
  9, 6, 8,
  4, 5, 5,
  _, _, 4,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, 4,
  _, _, _,
  _, _, 4,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  9, 10, 9,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  9, 10, 10,
  9, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  8, 10, 10,
  9, 10, 10,
  10, 10, 10,
  9, 9, 10,
  10, 10, 9,
  10, 10, 10,
  10, 10, 10,
  10, 10, 9,
  8, 8, 6,
  9, 9, 10,
  8, 7, 10,
  7, _, _,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  10, 9, 10,
  10, 10, 10,
  10, 10, 10,
  10, 10, 10,
  7, 9, 9,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  10, 10, 10,
  10, 10, 10,
  9, 8, 7,
  8, 5, 5,
  9, 4, 4,
  9, _, _,
  4, _, 8,
  _, 5, 6,
  _, 4, 4,
  _, _, 5,
  _, _, _,
  _, _, 5,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  4, 5, _,
  9, 6, 6,
  9, 7, 7,
  9, 7, 7,
  10, 6, 8,
  9, 6, 7,
  5, _, 6,
  _, _, 4,
  _, _, 6,
  4, _, 4,
  5, 5, 4,
  7, 4, 5 ;

 peakPower =
  59, 56, 51, 42, 42, 49, 67, 69, 63, 62, 62, 60, 53, 49, 54, 57, 52, 50, 47, 
    47, 47, 46, 43, 43, 43, 43, 44, 39, 36, 35, 36, 37, 33, 29, 29, 30, _, _, 
    _, _, _, _, _, _, 44, 44, 44, 44, 44, 43, 42, 41, 40, 39, 39, 39, 38, 38, 
    38, 37, 38, 39, 39, 38, 36, 34, 33, 32, 33, 33, 32, 32,
  55, 55, 58, 55, 59, _, _, 44, 44, 42, 43, 45, 51, 52, 55, 55, 51, 46, 44, 
    46, 45, 44, 42, 41, 42, _, _, _, 46, 41, 40, 40, 39, 38, 35, _, _, _, _, 
    _, _, _, _, _, _, _, 37, 36, 37, 36, 36, _, 33, _, _, _, _, _, _, _, 33, 
    _, _, _, _, _, 36, 37, 38, 39, 39, 39,
  56, 61, 58, 66, 67, 65, 52, 40, 40, 42, 41, 41, 39, 38, 40, 35, 33, 38, 42, 
    44, 38, 39, 37, 38, 32, 31, 35, 31, 46, 45, 43, 42, 42, 33, 31, 31, _, _, 
    _, _, _, _, _, _, 42, 39, 36, 32, 32, 33, 33, 33, 33, 33, 33, _, 31, 31, 
    _, 31, 33, 34, 33, 32, 32, 33, 33, _, _, _, _, 35,
  64, 68, 61, 65, 67, 59, 68, 67, 64, 63, 59, 54, 51, 54, 46, 35, 37, 33, 34, 
    30, 27, _, _, _, 33, 33, 31, 30, 41, 39, 38, 39, 40, 41, 41, 42, _, _, _, 
    _, _, _, _, _, 41, 40, 38, 36, 37, 38, 39, 39, 39, 37, 35, 33, _, 32, 33, 
    34, 33, 33, 34, 37, 39, 39, 37, 33, _, _, _, _,
  76, 77, 67, 68, 72, 73, 74, 73, 72, 73, 73, 74, 70, 67, 64, 62, 60, 61, 63, 
    64, 65, 67, 66, 63, 61, 60, 57, 55, 54, 51, 48, 47, 45, 43, 42, 42, _, _, 
    _, _, _, _, _, _, 54, 52, 50, 49, 47, 45, 43, 41, 41, 43, 44, 45, 44, 43, 
    42, 43, 43, 43, 42, 40, 38, 38, 38, 38, 37, 35, 35, 36,
  47, 47, 53, 62, 67, 64, 51, 40, 41, 44, 42, 40, 41, 43, 41, 39, 41, 41, 40, 
    38, 41, 45, 44, 39, 32, 35, 35, _, 43, 40, 39, 40, 29, 33, 32, 32, _, _, 
    _, _, _, _, _, _, 45, 44, 44, 43, 43, 41, 39, 37, 34, _, 32, 33, 35, 35, 
    35, 34, 33, 33, _, _, 32, 31, _, _, _, _, _, 31,
  65, _, 41, 50, 61, 59, 54, 56, 62, 64, 59, 59, 63, 69, 56, 54, 60, 64, 63, 
    50, 46, 44, 44, 42, 38, 40, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  63, 58, 48, 67, 70, 71, 72, 66, 59, 60, 63, 58, 59, 54, 55, 54, 58, 58, 57, 
    60, 61, 66, 61, 56, 55, 55, 51, 50, 52, 51, 50, 49, 48, 44, 42, 44, _, _, 
    _, _, _, _, _, _, 54, 54, 53, 52, 50, 49, 48, 48, 47, 45, 47, 51, 54, 56, 
    56, 55, 53, 50, 48, 46, 44, 44, 46, 47, 46, 44, 40, 37,
  64, 63, 58, 65, 73, 80, 75, 66, 58, 48, 47, 48, 62, 59, 48, 55, 57, 55, 63, 
    59, 48, 38, 43, 40, 40, 34, 33, 33, 33, 34, 45, 34, 35, 33, 33, 31, _, _, 
    _, _, _, _, _, _, 43, 42, 41, 39, 38, 37, 36, 31, 35, 36, 36, 37, 36, 36, 
    36, 36, 36, 36, 37, 38, 38, 38, 36, 34, 34, 35, 36, 38,
  19, 32, 42, 57, 62, 68, 64, 59, 55, 58, 59, 56, 56, 57, 60, 57, 53, 54, 52, 
    51, 49, 43, 38, 37, 45, 44, 42, 39, 38, 39, 37, 38, 36, 36, 33, 32, _, _, 
    _, _, _, _, _, _, 43, 41, 41, 40, 40, 39, 37, 37, 35, _, _, _, 36, 36, _, 
    38, 38, 38, 37, 36, 35, 35, 33, _, _, _, _, _,
  58, 63, 64, 62, 65, 69, 63, 58, 52, 51, 47, 48, 49, 43, 48, 49, 46, 40, 35, 
    33, 35, 46, 50, 53, 51, 43, 35, 35, 31, 30, 30, 42, 41, 39, 38, 37, _, _, 
    _, _, _, _, _, _, 37, 38, 39, 38, 38, 38, 38, 37, 36, 35, 36, 38, 40, 41, 
    40, 39, 40, 42, 44, 44, 43, 40, 37, 36, 35, 34, 33, 33,
  67, 67, 59, 58, 54, 51, 47, 60, 66, 73, 75, 66, 57, 65, 64, 62, 55, 47, 48, 
    51, 48, 43, 41, 42, 41, 39, 38, 38, 44, 43, 41, 39, 34, 40, 43, 37, _, _, 
    _, _, _, _, _, _, 48, 48, 46, 42, 39, 37, 36, 37, 36, 36, 36, 34, 32, 31, 
    _, 34, 37, 40, 42, 41, 39, 36, 33, 33, 33, 33, 33, 32,
  54, 57, 57, 66, 65, 64, 60, 58, 61, 56, 47, 46, 43, 44, 52, 54, 50, 55, 53, 
    46, 39, 34, 41, 42, 41, 46, 46, 45, 44, 43, 42, 41, 39, 38, 37, 35, _, _, 
    _, _, _, _, _, _, 48, 47, 45, 43, 42, 40, 38, 36, 35, _, 31, _, _, 30, 
    35, 36, 36, 37, 36, 35, 35, _, _, 32, 33, 33, _, _,
  42, 48, 50, 44, 42, 44, 42, 42, 51, 53, 46, 48, 50, 48, 45, 36, 36, 37, 37, 
    39, 38, 37, 34, 37, 35, 33, 32, _, 41, 40, 30, 40, 31, 39, 40, 40, _, _, 
    _, _, _, _, _, _, 41, 42, 45, 47, 49, 49, 49, 47, 46, 43, 41, 38, 35, 37, 
    38, 40, 42, 43, 42, 41, 38, 36, 34, 34, 34, 34, 34, 35,
  64, 62, 59, 75, 79, 68, 73, 73, 66, 60, 61, 60, 58, 64, 66, 64, 58, 62, 60, 
    50, 48, 58, 59, 56, 58, 57, 55, 49, 41, 33, 33, 31, 50, 34, 40, 44, _, _, 
    _, _, _, _, _, _, 57, 56, 56, 55, 53, 50, 46, 43, 41, 40, 38, 36, 36, 37, 
    38, 38, 40, 43, 45, 45, 44, 42, 40, 40, 41, 41, 40, 39,
  68, 74, 63, 68, 68, 56, 63, 63, 58, 57, 60, 57, 56, 56, 59, 61, 61, 56, 53, 
    51, 50, 48, 44, 42, 43, 41, 40, 40, 41, 42, 42, 39, 38, 33, 48, 47, _, _, 
    _, _, _, _, _, _, 48, 48, 48, 48, 47, 46, 44, 43, 41, 40, 39, 37, 39, 43, 
    46, 47, 46, 44, 41, 37, 34, 35, 37, 36, 36, 36, 38, 39,
  50, 51, 47, 69, 76, 76, 63, 57, 54, 52, 54, 53, 49, 40, 41, 50, 47, 60, 63, 
    51, 37, 31, 38, 41, 45, 37, 35, 41, 41, 44, 35, 51, 48, 45, 46, 45, _, _, 
    _, _, _, _, _, _, 43, 40, 36, 33, 34, 35, 36, 35, 34, _, _, _, 33, 33, 
    33, 33, _, 33, 33, 33, 32, 33, 34, 35, 34, 34, 34, 33,
  58, 58, 50, 59, 61, 65, 57, 56, 59, 60, 56, 57, 58, 58, 54, 44, 37, 39, 41, 
    38, 45, 41, _, _, _, _, _, _, 33, 32, 32, _, 30, _, _, 34, _, _, _, _, _, 
    _, _, _, 35, 35, 34, 33, 31, _, _, 33, 33, _, _, _, _, _, 33, 37, 37, 36, 
    35, _, _, _, 31, _, _, _, _, _,
  54, 60, 65, 70, 72, 70, 67, 65, 60, 51, 40, 38, 47, 50, 56, 57, 57, 51, 52, 
    46, 41, 45, 43, 38, 40, 33, 32, _, 33, 33, 43, 32, 40, 38, 37, _, _, _, 
    _, _, _, _, _, _, 44, _, _, _, 37, 36, 35, 35, 34, _, _, _, _, _, 34, _, 
    34, _, 32, 32, 32, 32, _, _, _, _, _, _,
  69, 64, 55, 65, 69, 69, 67, 63, 65, 62, 64, 70, 65, 55, 50, 56, 57, 57, 54, 
    51, 50, 48, 49, 50, 50, 48, 50, 50, 42, 41, 43, 43, 42, 39, 36, 35, _, _, 
    _, _, _, _, _, _, 49, 48, 47, 45, 44, 43, 42, 41, 40, 38, 37, 37, 38, 39, 
    39, 39, 40, 41, 40, 38, 36, 36, 37, 38, 38, 37, 34, 33,
  70, 67, 62, 67, 72, 73, 66, 66, 64, 61, 60, 57, 52, 51, 51, 55, 52, 52, 51, 
    51, 49, 51, 51, 47, 40, 35, 35, _, 46, 47, 38, 42, 41, 37, 35, 32, _, _, 
    _, _, _, _, _, _, 46, 45, 44, 42, 41, 39, 37, 35, _, 34, 36, 36, 35, 35, 
    37, 39, 41, 43, 43, 42, 40, 37, _, _, 35, 35, 34, 34,
  42, 50, 51, 53, 56, 53, 53, 61, 57, 43, 17, 104, _, _, _, 110, 0, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _,
  70, 70, 71, 71, 66, 72, 73, 73, 69, 69, 68, 66, 73, 73, 71, 71, 73, 73, 72, 
    71, 67, 66, 66, 65, 65, 60, 55, 51, 48, 45, 52, 68, 65, 36, 58, 49, _, _, 
    _, _, _, _, _, _, 54, 52, 49, 48, 48, 48, 48, 47, 45, 42, 41, 41, 45, 48, 
    50, 51, 49, 46, 42, 38, 39, 40, 40, 40, 38, 37, 34, _,
  64, 68, 67, 60, 53, 53, 62, 72, 72, 70, 64, 56, 56, 64, 64, 62, 61, 57, 53, 
    56, 57, 56, 54, 55, 60, 54, 44, 41, 55, 42, 42, 49, 47, 45, 44, _, _, _, 
    _, _, _, _, _, _, 44, 46, 45, 44, _, _, _, _, _, _, _, _, _, 41, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _,
  44, 56, 59, 61, 67, 70, 69, 61, 52, 54, 52, 49, 51, 53, 46, 44, 48, 43, 40, 
    39, 38, 38, 38, 38, 38, 37, 38, 38, 38, 38, 38, 38, 36, 35, 36, 37, _, _, 
    _, _, _, _, _, _, 37, 37, 36, 33, _, _, _, _, _, _, _, 34, _, 32, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _,
  50, 67, 74, 76, 73, 73, 73, 69, 67, 64, 59, 57, 54, 53, 50, 45, 46, 50, 52, 
    53, 51, 46, 43, 39, 34, 35, 36, _, 46, 45, 44, 43, 44, 46, 36, 34, _, _, 
    _, _, _, _, _, _, 45, 42, 38, 36, 36, _, 35, 35, 35, 34, _, 34, _, _, _, 
    _, _, 40, 42, 43, 42, 39, 37, 34, 34, 36, 37, 36 ;

 peakPowerBeam =
  40, 44, 59,
  43, 45, 56,
  42, 41, 51,
  37, 35, 42,
  39, 38, 42,
  59, 61, 49,
  70, 71, 67,
  71, 71, 69,
  67, 65, 63,
  67, 64, 62,
  63, 63, 62,
  56, 60, 60,
  48, 53, 53,
  44, 51, 49,
  48, 58, 54,
  47, 59, 57,
  43, 56, 52,
  41, 56, 50,
  42, 51, 47,
  49, 51, 47,
  50, 49, 47,
  48, 48, 46,
  48, 46, 43,
  48, 45, 43,
  46, 43, 43,
  44, 43, 43,
  44, 43, 44,
  39, 39, 39,
  35, 35, 36,
  34, 36, 35,
  36, 37, 36,
  38, 37, 37,
  33, 32, 33,
  30, 29, 29,
  30, 29, 29,
  31, 31, 30,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  45, 44, 44,
  44, 43, 44,
  44, 43, 44,
  44, 43, 44,
  43, 43, 44,
  43, 42, 43,
  42, 41, 42,
  40, 40, 41,
  39, 39, 40,
  38, 38, 39,
  39, 38, 39,
  38, 38, 39,
  38, 38, 38,
  38, 37, 38,
  38, 37, 38,
  37, 37, 37,
  36, 38, 38,
  37, 38, 39,
  37, 39, 39,
  37, 38, 38,
  36, 38, 36,
  35, 37, 34,
  34, 36, 33,
  33, 34, 32,
  _, 32, 33,
  _, 33, 33,
  31, 33, 32,
  _, 32, 32,
  41, 36, 55,
  51, 54, 55,
  61, _, 58,
  58, 61, 55,
  55, 63, 59,
  52, 54, _,
  44, 44, _,
  40, 45, 44,
  40, 42, 44,
  37, 36, 42,
  _, _, 43,
  _, 41, 45,
  40, 54, 51,
  47, 57, 52,
  53, 59, 55,
  55, 56, 55,
  52, 49, 51,
  48, 43, 46,
  46, 43, 44,
  47, 49, 46,
  44, 43, 45,
  46, 43, 44,
  45, 40, 42,
  43, 40, 41,
  43, 40, 42,
  _, _, _,
  _, _, _,
  _, _, _,
  _, 42, 46,
  _, 38, 41,
  _, 38, 40,
  _, 38, 40,
  _, 36, 39,
  _, 36, 38,
  _, _, 35,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, 37,
  _, _, 36,
  _, _, 37,
  _, _, 36,
  _, _, 36,
  _, _, _,
  _, _, 33,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, 33,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, 36,
  _, _, 37,
  _, 37, 38,
  _, _, 39,
  _, _, 39,
  _, _, 39,
  57, 57, 56,
  63, 62, 61,
  63, 61, 58,
  68, 67, 66,
  68, 67, 67,
  64, 62, 65,
  53, 51, 52,
  42, 41, 40,
  38, 43, 40,
  35, 44, 42,
  45, 43, 41,
  42, 43, 41,
  40, 44, 39,
  42, 43, 38,
  46, 45, 40,
  43, 40, 35,
  42, 42, 33,
  46, 47, 38,
  51, 45, 42,
  49, 47, 44,
  39, 44, 38,
  37, 42, 39,
  38, 43, 37,
  37, 44, 38,
  32, 36, 32,
  37, 36, 31,
  35, 38, 35,
  34, 36, 31,
  47, 50, 46,
  44, 49, 45,
  41, 46, 43,
  40, 45, 42,
  40, 44, 42,
  33, 31, 33,
  32, 31, 31,
  31, 29, 31,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  42, 42, 42,
  39, 39, 39,
  36, 37, 36,
  35, 34, 32,
  _, 34, 32,
  _, 34, 33,
  _, 33, 33,
  33, 34, 33,
  34, 32, 33,
  _, _, 33,
  _, _, 33,
  30, _, _,
  _, _, 31,
  _, 32, 31,
  _, 32, _,
  _, 32, 31,
  35, 34, 33,
  37, 34, 34,
  38, 34, 33,
  39, 33, 32,
  40, 33, 32,
  _, 34, 33,
  _, _, 33,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, 35,
  66, 66, 64,
  69, 65, 68,
  62, 60, 61,
  64, 61, 65,
  61, 59, 67,
  61, 57, 59,
  71, 66, 68,
  68, 63, 67,
  64, 60, 64,
  63, 58, 63,
  59, 54, 59,
  54, 51, 54,
  52, 49, 51,
  59, 51, 54,
  49, 41, 46,
  37, 33, 35,
  39, 34, 37,
  33, _, 33,
  36, 35, 34,
  32, _, 30,
  28, _, 27,
  _, _, _,
  _, _, _,
  _, _, _,
  33, _, 33,
  33, 32, 33,
  32, _, 31,
  31, _, 30,
  45, 40, 41,
  43, 40, 39,
  41, 37, 38,
  42, 37, 39,
  44, 39, 40,
  46, 40, 41,
  48, 39, 41,
  45, 38, 42,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  48, 37, 41,
  49, 36, 40,
  52, 35, 38,
  60, _, 36,
  39, _, 37,
  41, 34, 38,
  42, 36, 39,
  42, 36, 39,
  41, 36, 39,
  39, 35, 37,
  37, 34, 35,
  34, 34, 33,
  33, _, _,
  33, _, 32,
  32, _, 33,
  33, _, 34,
  34, _, 33,
  63, _, 33,
  61, _, 34,
  57, 35, 37,
  45, _, 39,
  50, _, 39,
  51, _, 37,
  46, _, 33,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  76, 73, 76,
  77, 74, 77,
  65, 64, 67,
  66, 66, 68,
  71, 71, 72,
  73, 74, 73,
  75, 75, 74,
  76, 74, 73,
  72, 75, 72,
  72, 74, 73,
  74, 72, 73,
  71, 73, 74,
  66, 70, 70,
  63, 67, 67,
  63, 65, 64,
  63, 65, 62,
  62, 64, 60,
  61, 62, 61,
  64, 64, 63,
  66, 67, 64,
  68, 68, 65,
  68, 69, 67,
  68, 68, 66,
  66, 66, 63,
  64, 63, 61,
  62, 61, 60,
  59, 57, 57,
  56, 55, 55,
  54, 53, 54,
  52, 50, 51,
  49, 48, 48,
  47, 47, 47,
  47, 46, 45,
  44, 44, 43,
  43, 43, 42,
  42, 40, 42,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  55, 54, 54,
  54, 52, 52,
  52, 51, 50,
  51, 50, 49,
  49, 49, 47,
  47, 46, 45,
  44, 44, 43,
  43, 42, 41,
  43, 42, 41,
  44, 42, 43,
  45, 43, 44,
  44, 43, 45,
  42, 42, 44,
  41, 40, 43,
  43, 41, 42,
  45, 42, 43,
  46, 43, 43,
  45, 43, 43,
  43, 42, 42,
  41, 40, 40,
  39, 38, 38,
  40, 38, 38,
  40, 39, 38,
  40, 39, 38,
  39, 37, 37,
  37, 35, 35,
  36, 35, 35,
  _, 36, 36,
  49, 51, 47,
  50, 49, 47,
  56, 56, 53,
  64, 66, 62,
  65, 70, 67,
  57, 61, 64,
  49, 52, 51,
  40, 43, 40,
  44, 44, 41,
  45, 48, 44,
  42, 46, 42,
  40, 42, 40,
  41, 42, 41,
  43, 44, 43,
  41, 45, 41,
  39, 44, 39,
  43, 43, 41,
  42, 42, 41,
  38, 41, 40,
  39, 40, 38,
  42, 43, 41,
  44, 45, 45,
  43, 46, 44,
  39, 41, 39,
  32, 33, 32,
  36, 38, 35,
  34, 37, 35,
  31, 34, _,
  43, 45, 43,
  44, 43, 40,
  40, 42, 39,
  42, 44, 40,
  32, 32, 29,
  34, 34, 33,
  33, 34, 32,
  32, 33, 32,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  43, 45, 45,
  41, 44, 44,
  40, 43, 44,
  40, 42, 43,
  39, 42, 43,
  38, 41, 41,
  37, 40, 39,
  35, 37, 37,
  32, 35, 34,
  _, 35, _,
  33, 35, 32,
  34, 35, 33,
  35, 36, 35,
  35, 36, 35,
  35, 36, 35,
  36, 35, 34,
  35, 34, 33,
  34, 35, 33,
  _, 36, _,
  _, 33, _,
  _, _, 32,
  _, _, 31,
  _, _, _,
  _, _, _,
  _, _, _,
  36, _, _,
  35, _, _,
  _, 32, 31,
  _, _, 65,
  _, 48, _,
  39, 40, 41,
  37, 38, 50,
  54, 55, 61,
  58, 59, 59,
  57, 57, 54,
  59, 58, 56,
  64, 65, 62,
  65, 66, 64,
  64, 61, 59,
  63, 55, 59,
  62, 60, 63,
  64, 65, 69,
  67, 62, 56,
  63, 59, 54,
  61, 60, 60,
  63, 64, 64,
  61, 62, 63,
  48, 50, 50,
  47, 50, 46,
  43, 46, 44,
  45, 47, 44,
  43, 44, 42,
  37, 35, 38,
  37, 36, 40,
  34, _, _,
  _, _, _,
  34, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  62, 61, 63,
  54, 52, 58,
  47, 47, 48,
  69, 68, 67,
  72, 69, 70,
  73, 71, 71,
  74, 75, 72,
  67, 69, 66,
  59, 59, 59,
  60, 60, 60,
  63, 63, 63,
  58, 59, 58,
  60, 62, 59,
  56, 56, 54,
  56, 56, 55,
  55, 56, 54,
  58, 59, 58,
  59, 61, 58,
  57, 56, 57,
  57, 54, 60,
  62, 62, 61,
  67, 67, 66,
  62, 61, 61,
  55, 56, 56,
  55, 57, 55,
  55, 56, 55,
  50, 53, 51,
  50, 53, 50,
  53, 51, 52,
  53, 51, 51,
  52, 49, 50,
  50, 48, 49,
  49, 47, 48,
  47, 43, 44,
  44, 42, 42,
  42, 42, 44,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  54, 53, 54,
  53, 52, 54,
  53, 52, 53,
  51, 51, 52,
  50, 49, 50,
  48, 48, 49,
  47, 47, 48,
  45, 45, 48,
  44, 44, 47,
  44, 44, 45,
  47, 46, 47,
  50, 50, 51,
  53, 53, 54,
  55, 55, 56,
  55, 55, 56,
  53, 54, 55,
  51, 51, 53,
  49, 49, 50,
  47, 47, 48,
  45, 45, 46,
  44, 44, 44,
  45, 45, 44,
  48, 46, 46,
  49, 47, 47,
  48, 47, 46,
  46, 45, 44,
  42, 42, 40,
  40, 39, 37,
  60, 62, 64,
  60, 62, 63,
  52, 54, 58,
  67, 64, 65,
  71, 75, 73,
  78, 82, 80,
  76, 77, 75,
  66, 67, 66,
  57, 59, 58,
  49, 50, 48,
  47, 48, 47,
  51, 52, 48,
  63, 64, 62,
  59, 60, 59,
  50, 51, 48,
  57, 60, 55,
  58, 60, 57,
  60, 61, 55,
  66, 69, 63,
  60, 64, 59,
  48, 51, 48,
  39, 41, 38,
  44, 46, 43,
  40, 43, 40,
  42, 41, 40,
  36, 36, 34,
  34, 35, 33,
  33, 33, 33,
  34, 35, 33,
  32, 35, 34,
  47, 49, 45,
  34, 36, 34,
  37, 39, 35,
  35, 35, 33,
  33, 34, 33,
  32, 33, 31,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  45, 45, 43,
  43, 43, 42,
  42, 42, 41,
  40, 41, 39,
  36, 39, 38,
  _, 38, 37,
  _, 36, 36,
  _, 36, 31,
  _, 37, 35,
  37, 37, 36,
  36, 38, 36,
  37, 38, 37,
  37, 37, 36,
  36, 38, 36,
  36, 38, 36,
  36, 38, 36,
  36, 39, 36,
  37, 39, 36,
  38, 40, 37,
  39, 40, 38,
  39, 41, 38,
  38, 40, 38,
  37, 39, 36,
  37, 37, 34,
  36, 37, 34,
  _, _, 35,
  35, 36, 36,
  _, 38, 38,
  37, 32, 19,
  42, 39, 32,
  53, 50, 42,
  63, 60, 57,
  68, 63, 62,
  69, 67, 68,
  66, 63, 64,
  63, 59, 59,
  60, 57, 55,
  61, 59, 58,
  61, 58, 59,
  59, 58, 56,
  59, 58, 56,
  61, 57, 57,
  62, 58, 60,
  60, 55, 57,
  57, 55, 53,
  57, 55, 54,
  55, 52, 52,
  52, 51, 51,
  50, 50, 49,
  45, 43, 43,
  43, 41, 38,
  42, 40, 37,
  49, 46, 45,
  46, 45, 44,
  44, 44, 42,
  43, 41, 39,
  43, 38, 38,
  43, 39, 39,
  42, 38, 37,
  41, 38, 38,
  39, 37, 36,
  37, 36, 36,
  35, 34, 33,
  33, 33, 32,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  46, 45, 43,
  45, 43, 41,
  44, 43, 41,
  44, 43, 40,
  43, 42, 40,
  41, 40, 39,
  40, 39, 37,
  38, 37, 37,
  36, 35, 35,
  _, _, _,
  33, _, _,
  35, 33, _,
  37, 37, 36,
  38, 40, 36,
  39, 39, _,
  40, 38, 38,
  41, 38, 38,
  41, 37, 38,
  40, 37, 37,
  40, 36, 36,
  38, 36, 35,
  36, 36, 35,
  34, 34, 33,
  33, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  67, 67, 58,
  72, 73, 63,
  70, 70, 64,
  66, 66, 62,
  67, 68, 65,
  68, 71, 69,
  62, 65, 63,
  57, 60, 58,
  56, 57, 52,
  53, 54, 51,
  50, 50, 47,
  50, 49, 48,
  51, 49, 49,
  47, 46, 43,
  51, 55, 48,
  53, 55, 49,
  50, 50, 46,
  43, 44, 40,
  36, 39, 35,
  33, 37, 33,
  39, 40, 35,
  46, 48, 46,
  51, 52, 50,
  54, 56, 53,
  50, 53, 51,
  41, 46, 43,
  35, 37, 35,
  34, 34, 35,
  31, 32, 31,
  31, 31, 30,
  29, 30, 30,
  42, 43, 42,
  40, 41, 41,
  39, 39, 39,
  38, 36, 38,
  37, 36, 37,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  37, 38, 37,
  37, 39, 38,
  38, 40, 39,
  39, 40, 38,
  39, 40, 38,
  39, 40, 38,
  39, 40, 38,
  38, 39, 37,
  38, 38, 36,
  37, 36, 35,
  39, 39, 36,
  40, 41, 38,
  42, 43, 40,
  42, 43, 41,
  41, 42, 40,
  40, 41, 39,
  40, 41, 40,
  42, 44, 42,
  44, 46, 44,
  44, 46, 44,
  44, 45, 43,
  42, 42, 40,
  39, 39, 37,
  37, 38, 36,
  37, 37, 35,
  36, 35, 34,
  35, _, 33,
  _, _, 33,
  63, 64, 67,
  62, 61, 67,
  59, 58, 59,
  60, 58, 58,
  55, 54, 54,
  52, 53, 51,
  53, 52, 47,
  65, 66, 60,
  68, 67, 66,
  75, 76, 73,
  75, 75, 75,
  66, 66, 66,
  58, 57, 57,
  65, 67, 65,
  65, 67, 64,
  62, 62, 62,
  56, 55, 55,
  50, 49, 47,
  49, 49, 48,
  50, 50, 51,
  48, 48, 48,
  43, 43, 43,
  43, 41, 41,
  45, 42, 42,
  42, 41, 41,
  41, 41, 39,
  39, 39, 38,
  39, 38, 38,
  46, 49, 44,
  44, 49, 43,
  41, 47, 41,
  39, 43, 39,
  33, 32, 34,
  43, 43, 40,
  46, 46, 43,
  43, 40, 37,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  50, 49, 48,
  48, 48, 48,
  45, 46, 46,
  41, 43, 42,
  38, 40, 39,
  37, 39, 37,
  37, 38, 36,
  37, 38, 37,
  37, 37, 36,
  36, 36, 36,
  37, 35, 36,
  36, 33, 34,
  35, 33, 32,
  35, 33, 31,
  35, 33, _,
  38, 35, 34,
  42, 39, 37,
  44, 41, 40,
  45, 42, 42,
  43, 41, 41,
  41, 39, 39,
  37, 36, 36,
  34, 33, 33,
  33, 32, 33,
  34, 34, 33,
  33, _, 33,
  32, 34, 33,
  _, 33, 32,
  53, 57, 54,
  55, 58, 57,
  63, 66, 57,
  70, 71, 66,
  65, 66, 65,
  69, 69, 64,
  75, 66, 60,
  71, 64, 58,
  64, 67, 61,
  59, 58, 56,
  46, 46, 47,
  44, 49, 46,
  45, 50, 43,
  48, 50, 44,
  58, 60, 52,
  57, 60, 54,
  54, 60, 50,
  58, 62, 55,
  55, 59, 53,
  48, 51, 46,
  40, 45, 39,
  41, 45, 34,
  49, 49, 41,
  48, 50, 42,
  46, 49, 41,
  50, 52, 46,
  48, 50, 46,
  46, 49, 45,
  47, 50, 44,
  46, 49, 43,
  45, 48, 42,
  43, 47, 41,
  41, 46, 39,
  40, 45, 38,
  39, 43, 37,
  37, 42, 35,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  47, 55, 48,
  46, 53, 47,
  46, 52, 45,
  45, 50, 43,
  44, 48, 42,
  42, 46, 40,
  40, 44, 38,
  38, 41, 36,
  37, 39, 35,
  36, 38, _,
  _, 37, 31,
  _, 35, _,
  34, 34, _,
  37, 37, 30,
  40, 39, 35,
  41, 42, 36,
  41, 42, 36,
  40, 42, 37,
  37, 40, 36,
  35, 38, 35,
  34, 37, 35,
  35, 36, _,
  35, 37, _,
  35, 38, 32,
  35, 38, 33,
  34, 38, 33,
  33, 36, _,
  _, 36, _,
  47, 41, 42,
  51, 45, 48,
  52, 46, 50,
  44, 39, 44,
  44, 38, 42,
  45, 39, 44,
  45, 38, 42,
  45, 40, 42,
  52, 47, 51,
  52, 46, 53,
  45, 40, 46,
  47, 41, 48,
  49, 42, 50,
  47, 42, 48,
  44, 39, 45,
  35, 30, 36,
  37, 31, 36,
  37, 30, 37,
  37, 31, 37,
  39, 34, 39,
  37, 33, 38,
  35, 31, 37,
  33, 28, 34,
  36, _, 37,
  32, _, 35,
  31, _, 33,
  _, _, 32,
  _, _, _,
  40, 36, 41,
  40, _, 40,
  29, 27, 30,
  40, _, 40,
  27, _, 31,
  39, _, 39,
  39, 36, 40,
  40, 37, 40,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  41, 37, 41,
  42, 38, 42,
  45, 41, 45,
  47, 42, 47,
  48, 43, 49,
  48, 43, 49,
  47, 42, 49,
  46, 41, 47,
  45, 38, 46,
  43, 37, 43,
  41, 35, 41,
  39, _, 38,
  38, _, 35,
  38, 33, 37,
  38, 33, 38,
  40, 34, 40,
  42, 36, 42,
  43, 36, 43,
  42, 37, 42,
  40, 35, 41,
  41, _, 38,
  45, 34, 36,
  49, 34, 34,
  52, _, 34,
  52, _, 34,
  _, _, 34,
  _, _, 34,
  48, 34, 35,
  64, 63, 64,
  62, 53, 62,
  60, 58, 59,
  76, 75, 75,
  78, 77, 79,
  68, 66, 68,
  75, 72, 73,
  73, 71, 73,
  64, 62, 66,
  61, 59, 60,
  62, 59, 61,
  59, 58, 60,
  60, 58, 58,
  66, 64, 64,
  66, 63, 66,
  63, 61, 64,
  57, 58, 58,
  64, 63, 62,
  61, 61, 60,
  50, 52, 50,
  49, 50, 48,
  58, 57, 58,
  59, 57, 59,
  59, 57, 56,
  59, 59, 58,
  57, 56, 57,
  56, 51, 55,
  50, 46, 49,
  41, 36, 41,
  33, 31, 33,
  33, 33, 33,
  32, 32, 31,
  51, 50, 50,
  38, 35, 34,
  43, 41, 40,
  44, 44, 44,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  56, 57, 57,
  56, 56, 56,
  55, 54, 56,
  55, 52, 55,
  53, 49, 53,
  50, 46, 50,
  47, 43, 46,
  44, 41, 43,
  41, 40, 41,
  39, 38, 40,
  38, _, 38,
  35, 34, 36,
  36, 35, 36,
  39, 36, 37,
  40, 36, 38,
  40, 38, 38,
  43, 40, 40,
  46, 43, 43,
  48, 45, 45,
  48, 45, 45,
  46, 42, 44,
  43, 40, 42,
  41, 39, 40,
  41, 40, 40,
  43, 40, 41,
  47, 40, 41,
  50, 39, 40,
  51, 39, 39,
  67, 73, 68,
  59, 64, 74,
  57, 62, 63,
  59, 64, 68,
  60, 62, 68,
  56, 65, 56,
  60, 65, 63,
  60, 64, 63,
  58, 61, 58,
  55, 59, 57,
  58, 63, 60,
  51, 57, 57,
  50, 56, 56,
  54, 62, 56,
  59, 67, 59,
  60, 69, 61,
  61, 66, 61,
  56, 61, 56,
  51, 57, 53,
  50, 56, 51,
  53, 58, 50,
  51, 54, 48,
  44, 51, 44,
  41, 49, 42,
  40, 48, 43,
  40, 46, 41,
  40, 46, 40,
  42, 46, 40,
  43, 48, 41,
  44, 49, 42,
  40, 46, 42,
  38, 43, 39,
  36, 40, 38,
  34, 39, 33,
  49, 56, 48,
  49, 55, 47,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  49, 55, 48,
  49, 55, 48,
  49, 55, 48,
  48, 55, 48,
  47, 54, 47,
  46, 52, 46,
  44, 50, 44,
  42, 48, 43,
  42, 45, 41,
  41, 43, 40,
  40, _, 39,
  40, 46, 37,
  41, 49, 39,
  43, 52, 43,
  44, 54, 46,
  45, 54, 47,
  44, 53, 46,
  43, 49, 44,
  42, 44, 41,
  40, 40, 37,
  40, 39, 34,
  39, 39, 35,
  39, 39, 37,
  40, 40, 36,
  40, 40, 36,
  42, 42, 36,
  43, 44, 38,
  42, 44, 39,
  55, 44, 50,
  57, 49, 51,
  51, 45, 47,
  74, 66, 69,
  75, 70, 76,
  71, 68, 76,
  57, 59, 63,
  55, 56, 57,
  52, 51, 54,
  53, 47, 52,
  54, 48, 54,
  53, 47, 53,
  49, 45, 49,
  40, 41, 40,
  44, 41, 41,
  59, 41, 50,
  54, 44, 47,
  63, 55, 60,
  63, 55, 63,
  51, 46, 51,
  37, 37, 37,
  32, _, 31,
  48, 37, 38,
  49, 39, 41,
  48, 37, 45,
  40, 32, 37,
  40, 34, 35,
  41, 31, 41,
  44, 32, 41,
  45, 34, 44,
  36, 31, 35,
  54, 41, 51,
  50, 40, 48,
  48, 39, 45,
  48, 39, 46,
  48, 38, 45,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  46, 37, 43,
  42, 37, 40,
  38, 36, 36,
  36, 32, 33,
  35, 33, 34,
  36, 35, 35,
  35, 35, 36,
  35, 35, 35,
  35, 36, 34,
  35, 36, _,
  34, 36, _,
  _, 36, _,
  36, 37, 33,
  _, 37, 33,
  _, 37, 33,
  _, 37, 33,
  34, 37, _,
  33, 37, 33,
  _, 37, 33,
  _, 36, 33,
  34, 36, 32,
  34, 36, 33,
  35, 35, 34,
  36, 36, 35,
  35, 35, 34,
  37, _, 34,
  36, 34, 34,
  36, _, 33,
  51, 58, 58,
  48, 47, 58,
  44, 40, 50,
  62, 52, 59,
  61, 57, 61,
  60, 55, 65,
  60, 58, 57,
  56, 59, 56,
  56, 61, 59,
  58, 61, 60,
  58, 60, 56,
  58, 61, 57,
  60, 64, 58,
  58, 64, 58,
  51, 57, 54,
  43, 45, 44,
  38, 43, 37,
  41, 44, 39,
  44, 49, 41,
  42, 43, 38,
  39, 37, 45,
  _, 33, 41,
  _, 33, _,
  _, _, _,
  31, _, _,
  29, _, _,
  _, 29, _,
  _, _, _,
  35, 37, 33,
  34, 38, 32,
  34, 38, 32,
  33, 37, _,
  32, 35, 30,
  32, 34, _,
  33, 36, _,
  35, 39, 34,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  35, 41, 35,
  36, 41, 35,
  35, 40, 34,
  33, 38, 33,
  32, 36, 31,
  _, 38, _,
  32, 35, _,
  33, 36, 33,
  34, 36, 33,
  32, 35, _,
  _, 34, _,
  _, 35, _,
  _, 35, _,
  _, 37, _,
  34, 38, 33,
  37, 40, 37,
  37, 41, 37,
  37, 40, 36,
  36, 37, 35,
  33, 33, _,
  33, 34, _,
  32, 34, _,
  33, 33, 31,
  32, 33, _,
  _, 32, _,
  _, _, _,
  31, 33, _,
  _, 34, _,
  56, 57, 54,
  62, 64, 60,
  66, 69, 65,
  71, 73, 70,
  74, 76, 72,
  72, 74, 70,
  70, 69, 67,
  68, 67, 65,
  61, 60, 60,
  52, 49, 51,
  42, 43, 40,
  42, 45, 38,
  51, 51, 47,
  52, 54, 50,
  59, 58, 56,
  61, 60, 57,
  60, 59, 57,
  54, 53, 51,
  53, 53, 52,
  48, 47, 46,
  46, 46, 41,
  49, 52, 45,
  47, _, 43,
  41, 39, 38,
  41, 42, 40,
  35, 35, 33,
  33, _, 32,
  _, _, _,
  35, 35, 33,
  34, 35, 33,
  45, 48, 43,
  32, 32, 32,
  42, 45, 40,
  40, 43, 38,
  41, 41, 37,
  48, 48, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, 54, 44,
  _, _, _,
  _, 61, _,
  _, 59, _,
  50, 54, 37,
  44, 50, 36,
  39, 44, 35,
  37, 37, 35,
  _, _, 34,
  _, _, _,
  _, _, _,
  33, _, _,
  33, _, _,
  33, 38, _,
  35, 38, 34,
  35, 39, _,
  _, 36, 34,
  _, 35, _,
  _, 34, 32,
  _, 34, 32,
  32, 33, 32,
  _, _, 32,
  _, 34, _,
  _, _, _,
  33, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  65, 67, 69,
  63, 64, 64,
  57, 58, 55,
  69, 70, 65,
  72, 73, 69,
  72, 72, 69,
  69, 67, 67,
  65, 65, 63,
  67, 67, 65,
  63, 63, 62,
  67, 66, 64,
  72, 72, 70,
  64, 66, 65,
  56, 58, 55,
  54, 54, 50,
  60, 60, 56,
  61, 62, 57,
  58, 60, 57,
  57, 57, 54,
  55, 54, 51,
  54, 52, 50,
  54, 52, 48,
  52, 51, 49,
  50, 54, 50,
  49, 54, 50,
  48, 51, 48,
  51, 53, 50,
  50, 53, 50,
  43, 44, 42,
  44, 45, 41,
  45, 45, 43,
  43, 45, 43,
  41, 44, 42,
  41, 41, 39,
  39, 37, 36,
  39, 37, 35,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  50, 52, 49,
  49, 51, 48,
  48, 50, 47,
  47, 48, 45,
  45, 46, 44,
  44, 45, 43,
  43, 44, 42,
  42, 43, 41,
  40, 41, 40,
  39, 39, 38,
  38, 38, 37,
  39, 38, 37,
  40, 40, 38,
  42, 41, 39,
  42, 42, 39,
  41, 44, 39,
  41, 43, 40,
  41, 43, 41,
  41, 42, 40,
  38, 39, 38,
  37, 37, 36,
  37, 38, 36,
  38, 40, 37,
  39, 41, 38,
  39, 41, 38,
  38, 39, 37,
  37, 38, 34,
  36, 38, 33,
  68, 65, 70,
  69, 64, 67,
  61, 58, 62,
  66, 60, 67,
  73, 70, 72,
  73, 69, 73,
  68, 63, 66,
  67, 64, 66,
  64, 63, 64,
  62, 61, 61,
  59, 58, 60,
  55, 54, 57,
  54, 50, 52,
  52, 48, 51,
  55, 53, 51,
  54, 51, 55,
  52, 49, 52,
  51, 47, 52,
  52, 47, 51,
  51, 47, 51,
  49, 46, 49,
  52, 50, 51,
  50, 48, 51,
  45, 43, 47,
  37, 35, 40,
  36, 34, 35,
  35, 31, 35,
  _, _, _,
  45, 43, 46,
  42, 44, 47,
  39, 35, 38,
  41, 37, 42,
  38, 38, 41,
  34, 35, 37,
  34, 32, 35,
  33, 30, 32,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  45, 42, 46,
  45, 42, 45,
  44, 41, 44,
  43, 39, 42,
  41, 37, 41,
  40, 36, 39,
  37, 34, 37,
  36, 33, 35,
  36, 32, _,
  36, 32, 34,
  38, 32, 36,
  39, _, 36,
  38, _, 35,
  37, _, 35,
  38, 33, 37,
  40, 37, 39,
  43, 40, 41,
  45, 41, 43,
  45, 41, 43,
  44, 39, 42,
  42, 36, 40,
  39, 34, 37,
  37, 32, _,
  37, _, _,
  37, _, 35,
  38, 32, 35,
  38, 34, 34,
  38, 35, 34,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  77, _, 70,
  82, 63, 70,
  80, 75, 71,
  71, 65, 71,
  68, _, 66,
  72, 71, 72,
  72, 71, 73,
  75, 73, 73,
  70, 70, 69,
  66, 64, 69,
  66, 74, 68,
  65, 71, 66,
  62, 63, 73,
  69, 68, 73,
  73, 69, 71,
  72, 70, 71,
  75, 75, 73,
  75, 75, 73,
  73, 73, 72,
  71, 73, 71,
  70, 70, 67,
  67, 71, 66,
  65, 70, 66,
  62, 68, 65,
  58, 67, 65,
  51, 64, 60,
  48, 61, 55,
  64, 64, 51,
  56, 65, 48,
  46, 45, 45,
  42, 44, 52,
  63, 74, 68,
  58, 73, 65,
  35, 62, 36,
  54, 50, 58,
  55, 47, 49,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  55, 46, 54,
  55, 65, 52,
  55, 65, 49,
  54, 47, 48,
  53, 48, 48,
  53, 50, 48,
  47, 49, 48,
  44, 47, 47,
  43, _, 45,
  41, _, 42,
  41, 58, 41,
  44, 43, 41,
  48, 46, 45,
  51, 49, 48,
  53, 51, 50,
  52, 51, 51,
  50, 52, 49,
  47, 46, 46,
  43, 41, 42,
  40, 39, 38,
  41, 39, 39,
  41, 40, 40,
  40, 39, 40,
  38, 38, 40,
  36, 36, 38,
  _, 35, 37,
  36, _, 34,
  33, _, _,
  67, 65, 64,
  72, 71, 68,
  70, 70, 67,
  62, 62, 60,
  54, 57, 53,
  50, 55, 53,
  63, 70, 62,
  74, 78, 72,
  75, 75, 72,
  74, 75, 70,
  64, 66, 64,
  60, 63, 56,
  59, 60, 56,
  62, 62, 64,
  62, 62, 64,
  62, 63, 62,
  61, 63, 61,
  58, 60, 57,
  55, 59, 53,
  60, 60, 56,
  58, 59, 57,
  57, 57, 56,
  55, 55, 54,
  57, 57, 55,
  60, 61, 60,
  52, 55, 54,
  44, 44, 44,
  40, 41, 41,
  55, 58, 55,
  42, 43, 42,
  41, 41, 42,
  52, 53, 49,
  49, 50, 47,
  46, 47, 45,
  44, 44, 44,
  43, 45, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, 44,
  _, 45, 46,
  _, _, 45,
  _, 44, 44,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, 41, _,
  _, _, _,
  _, _, _,
  _, _, 41,
  _, _, _,
  _, _, _,
  _, 43, _,
  _, 44, _,
  44, 44, _,
  44, _, _,
  43, _, _,
  44, _, _,
  _, _, _,
  _, _, _,
  42, _, _,
  44, _, _,
  45, _, _,
  44, 42, _,
  52, 53, 44,
  58, 60, 56,
  60, 61, 59,
  64, 63, 61,
  68, 67, 67,
  71, 70, 70,
  69, 67, 69,
  60, 58, 61,
  50, 50, 52,
  46, 46, 54,
  44, 48, 52,
  42, 46, 49,
  52, 51, 51,
  52, 50, 53,
  43, 44, 46,
  46, 44, 44,
  48, 45, 48,
  37, 34, 43,
  34, 33, 40,
  35, 31, 39,
  30, _, 38,
  _, _, 38,
  _, _, 38,
  _, 31, 38,
  _, _, 38,
  _, _, 37,
  _, _, 38,
  _, _, 38,
  _, _, 38,
  _, _, 38,
  39, 35, 38,
  39, 36, 38,
  40, 37, 36,
  40, 36, 35,
  39, 35, 36,
  44, 35, 37,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  49, 36, 37,
  42, 35, 37,
  34, 33, 36,
  _, _, 33,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, 34,
  _, _, _,
  _, _, 32,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  53, 54, 50,
  71, 70, 67,
  77, 77, 74,
  78, 78, 76,
  78, 77, 73,
  75, 76, 73,
  76, 75, 73,
  72, 71, 69,
  70, 69, 67,
  66, 66, 64,
  61, 61, 59,
  57, 57, 57,
  58, 54, 54,
  56, 54, 53,
  52, 49, 50,
  50, 48, 45,
  49, 49, 46,
  50, 51, 50,
  51, 54, 52,
  53, 53, 53,
  51, 49, 51,
  47, 47, 46,
  45, 43, 43,
  40, 38, 39,
  34, 34, 34,
  35, 37, 35,
  37, 34, 36,
  33, _, _,
  47, 47, 46,
  45, 45, 45,
  44, 44, 44,
  44, 43, 43,
  47, 43, 44,
  49, 45, 46,
  37, 34, 36,
  35, 34, 34,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  48, 45, 45,
  44, 42, 42,
  38, 38, 38,
  38, 34, 36,
  37, 35, 36,
  37, _, _,
  37, _, 35,
  _, 36, 35,
  _, 35, 35,
  _, _, 34,
  _, _, _,
  _, _, 34,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  40, 37, _,
  41, 40, 40,
  43, 42, 42,
  44, 43, 43,
  42, 42, 42,
  40, 38, 39,
  38, _, 37,
  _, _, 34,
  _, _, 34,
  37, _, 36,
  38, 34, 37,
  37, 33, 36 ;

 radVelocity =
  -4.48, -2.68, 0,
  -3.81, -4.03, 0.01,
  -2.99, -4.04, 0,
  -2.4, -4.24, -0.01,
  -2.06, -4.23, 0,
  -2.2, -3.6, 0.02,
  -2.31, -3.23, 0.02,
  -2.05, -2.61, 0.03,
  -1.2, -2.43, 0.05,
  -0.59, -3.06, 0.08,
  -0.45, -3.52, 0.06,
  -0.27, -3.67, 0.05,
  -0.26, -3.42, 0.03,
  -0.11, -3.05, -0.02,
  0.05, -2.76, -0.04,
  0.03, -2.63, -0.02,
  -0.04, -2.2, 0.02,
  0.01, -1.84, 0.04,
  0.14, -1.81, 0.05,
  0.24, -1.84, 0.05,
  0.28, -1.87, 0,
  0.26, -2.14, -0.02,
  0.3, -2.35, -0.04,
  0.48, -2.5, -0.03,
  1.04, -2.95, -0.04,
  1.54, -3.32, -0.02,
  1.77, -3.75, 0,
  2.1, -4.03, -0.01,
  1.97, -4.24, -0.02,
  1.26, -3.97, -0.03,
  1.08, -3.74, -0.04,
  0.8, -3.73, -0.02,
  0.82, -3.94, -0.03,
  0.83, -4.34, 0.05,
  0.87, -4.07, 0.05,
  0.89, -4.17, 0.11,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0.9, -4.35, -0.05,
  1.24, -4.56, -0.06,
  2, -4.83, -0.08,
  2.45, -5.24, -0.04,
  2.78, -5.66, -0.04,
  3.08, -5.93, -0.03,
  3.3, -6.24, -0.03,
  3.27, -6.54, 0.01,
  3.23, -6.77, -0.02,
  3.25, -6.98, -0.03,
  3.33, -7.15, -0.1,
  3.46, -7.48, -0.08,
  3.57, -7.78, -0.11,
  3.51, -8.01, -0.22,
  3.84, -7.36, -0.14,
  3.72, -7.39, -0.15,
  3.37, -6.71, -0.06,
  2.95, -5.99, -0.07,
  2.01, -5.47, -0.07,
  1.47, -4.75, -0.08,
  0.98, -4.41, -0.11,
  1.24, -4.36, -0.08,
  1.42, -4.3, -0.07,
  1.26, -4.32, 0.01,
  _, -2, 0.11,
  _, -1.89, 0.14,
  0.47, -1.56, 0.17,
  _, -1.64, 0.19,
  -0.05, 0.45, 1.37,
  -0.17, 0.8, 0.07,
  -0.1, _, -0.22,
  0.17, 0.74, 0.06,
  0.16, 0.81, 0.09,
  0.17, 0.48, _,
  -0.19, 0.18, _,
  -0.99, 0.18, 0.16,
  -0.87, 0.1, -0.03,
  -0.45, -7.52, 0,
  _, _, 0.13,
  _, -0.16, 0.1,
  0.19, -0.32, 0.05,
  0.08, -0.29, -0.03,
  0.24, -0.07, 0.13,
  0.39, 0.05, 0.26,
  0.39, -0.89, 0.37,
  0.59, -2.25, 0.36,
  0.46, -2.5, 0.2,
  0.46, -1.14, 0.13,
  0.57, -2.36, 0.2,
  0.71, -2.35, 0.16,
  0.54, -2.76, 0.04,
  0.43, -2.58, 0.02,
  0.31, -2.57, 0.03,
  _, _, _,
  _, _, _,
  _, _, _,
  _, -2.78, 0.06,
  _, -2.9, 0.02,
  _, -2.9, 0.05,
  _, -2.99, 0.04,
  _, -7.65, 0.06,
  _, -7.57, 0.09,
  _, _, 0.08,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, -0.11,
  _, _, -0.12,
  _, _, -0.1,
  _, _, -0.03,
  _, _, 0,
  _, _, _,
  _, _, 0.02,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, -10.5,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, -0.09,
  _, _, 0.03,
  _, -0.54, 0.03,
  _, _, 0,
  _, _, 0.04,
  _, _, 0,
  -2.27, -3.56, 0.04,
  -1.88, -3.51, 0.04,
  -0.95, -3.88, 0.04,
  -1.12, -3.82, 0.06,
  -1.47, -3.94, 0.07,
  -1.29, -4.19, 0.09,
  -1.03, -4.14, 0.09,
  -0.6, -3.75, -0.03,
  -0.4, -2.99, -0.08,
  -0.41, -2.81, -0.18,
  -0.27, -2.66, -0.1,
  -0.27, -2.43, -0.11,
  -0.25, -1.64, -0.11,
  -0.3, -1.56, -0.13,
  -0.26, -1.49, -0.11,
  -0.47, -1.44, -0.13,
  -1.21, -0.49, 0.07,
  -1.28, -0.26, 0.07,
  -0.86, -0.26, 0.11,
  -0.49, -0.28, 0.11,
  -0.36, -0.21, 0.07,
  -0.24, -0.17, 0.01,
  0.09, -0.24, 0.02,
  0.22, -0.29, -0.02,
  0.18, -0.39, 0.12,
  0.24, -0.42, -0.01,
  0.24, -0.39, -0.09,
  0.07, -0.49, 0.06,
  0.1, -0.63, -0.02,
  0.1, -0.78, -0.03,
  0.06, -0.95, -0.03,
  0.06, -1.2, -0.03,
  0.14, -1.64, -0.02,
  0.03, -1.71, -0.16,
  0.25, -2.44, -0.04,
  0.39, -3.06, -0.14,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0.37, -2.78, 0.02,
  0.28, -2.92, 0.01,
  0.47, -2.95, -0.01,
  0.5, -3.17, -0.04,
  _, -3.24, -0.03,
  _, -3.44, -0.02,
  _, -3.18, -0.03,
  0.03, -3.33, -0.18,
  0.19, -3.92, -0.38,
  _, _, -0.15,
  _, _, 0,
  -11.54, _, _,
  _, _, 0.1,
  _, -4.87, 0.02,
  _, -4.93, _,
  _, -4.61, -0.22,
  1.33, -4.01, -0.05,
  0.76, -3.78, -0.09,
  0.43, -3.65, -0.1,
  0.05, -3.29, -0.05,
  0.19, -3.28, 0.11,
  _, -3.48, 0.1,
  _, _, 0.27,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, 1.19,
  -3.02, -0.83, 0,
  -3.41, -0.64, 0,
  -3.37, -0.38, -0.03,
  -3, -0.56, 0.03,
  -2.56, -0.97, 0.06,
  -1.47, -1.6, 0.06,
  -1.04, -1.87, 0.02,
  -1.35, -1.63, 0.01,
  -1.8, -1.56, 0,
  -1.93, -1.67, 0.01,
  -1.93, -1.51, 0.02,
  -1.8, -0.94, 0.06,
  -1.35, -1.22, 0.08,
  -0.97, -1.56, 0.11,
  -0.89, -1.67, 0.09,
  -0.83, 5.04, 0.04,
  -1.27, 0.37, 0,
  -0.82, _, -0.05,
  -0.58, 0.98, -0.07,
  -1.09, _, -0.08,
  -1.83, _, -0.21,
  _, _, _,
  _, _, _,
  _, _, _,
  -2.34, _, 0.05,
  -2.27, 0.79, 0.05,
  -1.49, _, 0.18,
  -1.35, _, -0.01,
  -1.47, 0.38, 0.03,
  -1.4, 0.7, 0.04,
  -1.28, 0.37, 0.04,
  -1.12, 0.13, 0.01,
  -1.02, -0.02, 0.02,
  -0.95, 0.1, -0.02,
  -0.84, 0.45, -0.04,
  -0.66, 0.54, -0.04,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  -0.68, 0.6, -0.02,
  -1.04, 0.56, -0.01,
  -1.65, 0.72, -0.01,
  -2.31, _, 0.05,
  -3.11, _, 0.05,
  -3.05, -0.46, 0.07,
  -2.79, -0.53, 0.06,
  -2.34, -0.51, 0.05,
  -2, -0.63, 0.04,
  -1.76, -0.62, 0.04,
  -1.59, -0.46, 0.07,
  -1.58, -0.48, 0.03,
  -1.61, _, _,
  -2.06, _, -0.13,
  -1.98, _, -0.01,
  -1.72, _, 0.01,
  -0.6, _, -0.29,
  -1.31, _, -0.17,
  -0.91, _, -0.06,
  -0.79, -0.59, 0.02,
  -0.72, _, 0.04,
  -0.86, _, 0.05,
  -0.62, _, 0,
  -0.68, _, 0.08,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  -6.06, -3.73, -0.14,
  -5.86, -6.02, -0.2,
  -4.89, -6.64, -0.15,
  -2.63, -6.34, -0.1,
  -2.45, -5.86, -0.14,
  -2.9, -4.7, -0.11,
  -2.88, -4.07, -0.13,
  -2.89, -3.68, -0.13,
  -2.83, -3.48, -0.14,
  -2.9, -3.4, -0.21,
  -2.67, -3.07, -0.21,
  -3.05, -3.08, -0.16,
  -2.91, -2.95, -0.12,
  -2.86, -2.99, 0.02,
  -3.04, -2.9, -0.19,
  -2.97, -2.86, -0.24,
  -3.27, -3.11, -0.38,
  -3.34, -2.85, 0.05,
  -3.27, -2.38, 0.25,
  -3.25, -2.31, 0.21,
  -3.43, -2.27, 0.28,
  -3.55, -2.59, 0.52,
  -3.69, -2.98, 0.59,
  -4.02, -3.35, 0.54,
  -4.31, -4.15, 0.57,
  -3.58, -3.7, 0.51,
  -3.21, -4.25, 0.49,
  -2.61, -4.15, 0.49,
  -2, -3.94, 0.45,
  -1.95, -3.66, 0.39,
  -2.34, -3.57, 0.35,
  -2.59, -3.79, 0.38,
  -2.47, -4.17, 0.36,
  -2.38, -4.51, 0.41,
  -2.45, -4.71, 0.25,
  -2.72, -4.91, 0.16,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  -2.73, -4.81, 0.19,
  -2.85, -5, 0.15,
  -2.96, -5, 0.13,
  -3.15, -4.84, 0.13,
  -3.45, -4.55, 0.13,
  -3.81, -4.23, 0.13,
  -4.32, -4.17, 0.11,
  -5, -4.5, 0.09,
  -5.53, -5.19, 0.1,
  -5.64, -5.78, 0.08,
  -5.58, -6.22, 0.09,
  -5.58, -6.58, 0.06,
  -5.54, -7.36, 0.06,
  -4.81, -8.08, 0,
  -4.25, -8.07, 0.08,
  -3.82, -7.67, 0.11,
  -3.5, -7.13, 0.12,
  -3.24, -6.55, 0.15,
  -2.99, -5.96, 0.14,
  -2.74, -5.37, 0.09,
  -2.53, -4.76, -0.11,
  -2.19, -4.43, -0.12,
  -1.84, -4.23, -0.12,
  -1.58, -4.06, -0.11,
  -1.34, -3.98, -0.08,
  -1.06, -4.01, -0.05,
  -0.72, -3.92, -0.19,
  _, -2.93, -0.16,
  -4.69, -2.36, 0.2,
  -4.57, -4.46, 0.29,
  -4.57, -6.32, 0.24,
  -3.85, -5.85, 0.17,
  -3.13, -5.28, 0.1,
  -3.11, -4.66, 0.15,
  -2.14, -3.58, 0.17,
  -1.93, -3.09, 0.21,
  -2.09, -2.62, 0.25,
  -2.17, -2.5, 0.3,
  -2.22, -2.31, 0.29,
  -2.19, -2.02, 0.28,
  -2.14, -1.81, 0.32,
  -2.12, -1.82, 0.25,
  -2.1, -1.9, 0.14,
  -1.83, -2.06, 0.12,
  -1.43, -2.17, 0.08,
  -1.27, -2.22, 0.12,
  -1.4, -2.5, 0.07,
  -1.72, -2.43, -0.02,
  -2.07, -2.55, 0.02,
  -2.25, -2.74, 0.02,
  -2.44, -2.95, 0.03,
  -2.87, -2.86, -0.06,
  -3.43, -3.2, 0.02,
  -3.73, -3.5, 0.12,
  -3.85, -3.94, 0.09,
  -4.42, -5.21, _,
  -4.07, -4.37, 0,
  -5.02, -5.08, 0.08,
  -6.25, -5.36, 0.24,
  -6.68, -5.03, 0.26,
  -6.12, -5.06, 1.07,
  -6.54, -4.99, 0.79,
  -7.53, -4.54, 0.32,
  -8.22, -3.97, 0.3,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  -8.24, -4.18, 0.04,
  -8.43, -4.16, 0.01,
  -8.56, -4.29, 0.02,
  -8.54, -4.6, 0,
  -9, -4.86, 0.09,
  -8.81, -5.19, 0.22,
  -8.65, -5.35, 0.33,
  -8.69, -5.41, 0.48,
  -8.03, -5.86, -0.12,
  _, -6.16, _,
  -6.62, -5.54, 0.12,
  -6.66, -5.1, -0.07,
  -6.86, -5.52, -0.1,
  -6.73, -5.78, -0.09,
  -6.66, -5.74, -0.05,
  -7.07, -5.37, 0.13,
  -7.4, -5.61, 0.13,
  -4.87, -5.67, -0.01,
  _, -6.61, _,
  _, -5.79, _,
  _, _, 0.26,
  _, _, 0.16,
  _, _, _,
  _, _, _,
  _, _, _,
  -4.15, _, _,
  -3.47, _, _,
  _, 7.29, 0.48,
  _, _, 0,
  _, 1.85, _,
  -0.42, 1.82, 0.01,
  -0.69, 1.51, 0.1,
  -0.89, 1.32, -0.05,
  -0.65, 1.47, -0.06,
  -0.35, 1.24, -0.05,
  -0.48, 0.78, -0.1,
  -0.77, 0.61, 0.09,
  -1.24, 0.54, 0.06,
  -1.27, 0.59, 0.24,
  -1.25, 0.62, 0.38,
  -0.71, 0.85, 0.55,
  -0.9, 0.56, 0.51,
  -0.73, 0.84, 0.23,
  -0.52, 1.09, -0.03,
  -0.92, 1.37, 0.08,
  -1.32, 1.41, 0.11,
  -1.47, 1.18, -0.01,
  -1.19, 0.47, -0.08,
  -1.33, 0.34, -0.17,
  -2.07, 0.45, -0.2,
  -2.4, 0.55, -0.12,
  -2.45, 0.67, -0.2,
  -2.88, 0.52, -0.21,
  -3.48, 0.27, -0.39,
  -3.74, _, _,
  _, _, _,
  -4.84, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  -5.24, -4.12, -0.09,
  -4.32, -3.9, 0.02,
  -5.24, -5.19, 0.02,
  -4.47, -4.46, 0.02,
  -3.59, -3.7, 0.01,
  -2.68, -3.37, 0.03,
  -2.72, -2.65, 0.03,
  -2.6, -2.53, 0,
  -2.52, -2.53, 0.03,
  -2.98, -2.79, 0.06,
  -3.13, -3.01, 0.03,
  -3.22, -2.74, 0.01,
  -3.12, -2.46, 0.02,
  -2.99, -2.28, 0.02,
  -3.05, -2.02, 0,
  -3.55, -1.66, -0.04,
  -3.78, -1.18, -0.11,
  -3.64, -0.79, -0.14,
  -3.56, -0.67, -0.13,
  -3.37, -0.61, -0.13,
  -3.21, -0.98, -0.16,
  -3.3, -1.38, -0.19,
  -3.29, -2.01, -0.22,
  -2.97, -3.03, -0.23,
  -2.83, -3.31, -0.22,
  -2.74, -3.48, -0.23,
  -2.6, -3.6, -0.25,
  -2.33, -3.58, -0.17,
  -2.06, -3.79, -0.09,
  -1.91, -4.11, 0.01,
  -2.18, -4.25, 0.05,
  -2.69, -4.26, 0.03,
  -2.86, -4.18, 0.03,
  -2.97, -4.05, 0.06,
  -3.09, -3.72, 0.19,
  -2.68, -3.73, 0.2,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  -2.62, -4.04, 0.22,
  -2.6, -4.13, 0.22,
  -2.73, -4.21, 0.2,
  -2.86, -4.27, 0.18,
  -3.1, -4.3, 0.18,
  -3.52, -4.35, 0.18,
  -3.89, -4.28, 0.15,
  -4.41, -4.31, 0.14,
  -5.19, -4.23, 0.11,
  -5.71, -4.13, 0.13,
  -6.01, -4.55, 0.2,
  -6.25, -5.09, 0.16,
  -6.16, -5.59, 0.12,
  -5.92, -5.86, 0.08,
  -5.52, -6.06, 0.07,
  -4.91, -6.21, 0.07,
  -3.97, -6.24, 0.09,
  -2.77, -5.98, 0.06,
  -2.01, -5.29, 0.03,
  -1.83, -4.73, 0.02,
  -1.93, -4.46, 0.02,
  -1.94, -4.32, 0,
  -1.71, -4.33, -0.02,
  -1.58, -4.22, -0.01,
  -1.44, -4.02, 0,
  -1.31, -3.81, 0.03,
  -1.1, -3.36, -0.02,
  -0.76, -2.64, -0.06,
  -3.49, -2.68, -0.05,
  -3.26, -3.07, -0.04,
  -3.22, -3.45, -0.02,
  -3.22, -3.52, 0.01,
  -1.86, -3.8, -0.06,
  -3.24, -4, -0.09,
  -3.1, -3.93, -0.1,
  -2.67, -3.74, -0.11,
  -2.38, -3.7, -0.09,
  -1.86, -3.65, -0.14,
  -1.71, -3.51, -0.19,
  -1.12, -3.33, -0.17,
  -0.82, -3.12, -0.12,
  -0.83, -2.78, -0.12,
  -1.81, -0.56, -0.04,
  -2.32, 0.73, -0.03,
  -2.43, 1.2, -0.05,
  -1.96, 0.63, -0.05,
  -1.95, 0.38, -0.07,
  -2.07, 0.32, -0.07,
  -2.61, 0.76, -0.02,
  -2.67, 0.67, -0.05,
  -2.87, 0.39, -0.04,
  -3.14, 0.33, -0.04,
  -3.22, -0.01, -0.01,
  -3.3, -0.32, -0.08,
  -3.43, -0.4, -0.07,
  -3.06, -0.4, -0.11,
  -2.68, -0.63, -0.05,
  -2.88, -1, 0,
  -2.85, -1.3, -0.07,
  -2.93, -1.84, -0.03,
  -2.68, -1.61, -0.07,
  -2.19, -1.37, -0.09,
  -1.94, -1.07, 0.03,
  -1.26, -1.11, 0.11,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  -1.01, -1.27, 0.03,
  -0.72, -1.64, 0.03,
  -1.06, -1.93, 0,
  -1.35, -2.22, -0.03,
  -2.83, -2.48, -0.04,
  _, -2.55, -0.01,
  _, -2.6, 0.06,
  _, -2.81, -7,
  _, -2.87, 0,
  -1.23, -3.03, -0.17,
  -0.99, -3.12, -0.25,
  -0.88, -3.15, -0.15,
  -0.86, -3.11, -0.12,
  -1.35, -3.33, -0.08,
  -1.42, -3.41, -0.1,
  -1.3, -3.2, -0.02,
  -1.03, -3.16, -0.05,
  -0.81, -2.85, 0.1,
  -0.47, -2.46, 0.02,
  -0.47, -2.08, 0.05,
  -0.43, -1.84, 0,
  -0.33, -1.68, 0.01,
  0.15, -2.32, -0.01,
  0.41, -2.69, -0.16,
  0.43, -2.76, -0.31,
  _, _, -0.05,
  0.37, -0.86, -0.05,
  _, -0.75, 0.08,
  -5.29, -2.05, -0.49,
  -4.79, -3.27, 0.01,
  -4.64, -4.2, 0.02,
  -4.11, -3.98, 0.01,
  -2.78, -3.83, -0.04,
  -2.08, -3.26, 0.01,
  -1.81, -2.99, 0.04,
  -1.87, -2.68, 0.06,
  -1.9, -2.63, 0.04,
  -2.14, -2.86, 0.11,
  -2.47, -3.02, 0.2,
  -2.75, -3.08, 0.23,
  -3.19, -3.06, 0.21,
  -3.42, -2.92, 0.19,
  -3.56, -2.73, 0.14,
  -3.19, -3.2, 0.02,
  -3.09, -3.18, 0.07,
  -3.23, -3.28, 0.04,
  -3.45, -3.06, -0.02,
  -3.7, -2.93, -0.06,
  -4.08, -2.99, 0.08,
  -4.26, -3.09, 0,
  -4.36, -3.15, 0.06,
  -3.97, -2.93, -0.01,
  -3.65, -2.89, 0.03,
  -3.31, -3.28, -0.11,
  -3.38, -3.65, -0.09,
  -3.52, -3.58, -0.12,
  -3.67, -3.48, -0.08,
  -3.63, -3.71, 0.04,
  -3.36, -3.73, 0.01,
  -3.18, -3.79, 0.07,
  -3.25, -3.81, 0.05,
  -3.03, -3.65, 0.07,
  -2.63, -3.04, -0.32,
  -3.37, -3.38, 0.24,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  -3.43, -3.83, -0.05,
  -3.65, -3.89, -0.01,
  -3.87, -3.96, -0.06,
  -4.23, -3.84, -0.03,
  -4.55, -3.76, -0.02,
  -4.9, -3.67, -0.16,
  -5.21, -3.75, -0.41,
  -5.61, -3.63, 0.03,
  -6.22, -3.83, 0.01,
  _, _, _,
  -6.76, _, _,
  -6.3, -11.29, _,
  -5.81, -6.02, -0.24,
  -5.25, -6.49, -0.32,
  -4.6, -6.78, _,
  -3.34, -5.64, -0.26,
  -2.84, -5.47, -0.03,
  -2.61, -5.33, 0,
  -2.16, -5.03, 0.02,
  -1.48, -4.98, 0,
  -1.32, -4.9, 0.07,
  -1.13, -4.35, 0.16,
  -2.2, -4.03, 0.21,
  -3.39, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  -0.76, 0.59, 0.04,
  -0.85, 0.52, -0.05,
  -0.89, 0.95, 0.02,
  -0.76, 1.59, 0.03,
  -0.33, 2.54, 0.06,
  -0.33, 3.18, 0.02,
  -0.32, 3.74, -0.01,
  -0.35, 4.14, -0.03,
  -1.25, 3.8, -0.03,
  -1.59, 3.76, -0.04,
  -1.68, 3.76, -0.1,
  -1.86, 3.48, -0.16,
  -1.76, 3.12, -0.19,
  -1.31, 2.29, -0.34,
  -0.6, 2.37, 0,
  -0.36, 2.44, -0.02,
  -0.44, 2.43, 0.04,
  -0.23, 2.3, -0.04,
  0.25, 2.35, 0.04,
  -0.13, 2.41, 0.15,
  -0.01, 2.54, 0.16,
  -0.13, 2.58, 0.15,
  0.06, 2.17, 0.12,
  0.12, 2.41, 0.13,
  0.05, 2.88, 0.13,
  -0.03, 3.23, 0.14,
  -0.46, 2.99, 0.11,
  -0.68, 2.98, -0.25,
  -0.83, 2.92, -0.12,
  -1.03, 3.04, -0.02,
  -0.4, 3.29, -0.11,
  -0.71, 2.92, -0.16,
  -0.88, 2.91, -0.2,
  -1.08, 2.85, -0.19,
  -0.98, 2.43, -0.23,
  -0.83, 2.04, -0.3,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  -0.16, 1.88, -0.32,
  0.2, 1.98, -0.15,
  0.26, 2.34, -0.15,
  0.06, 2.7, -0.31,
  -0.12, 3.05, -0.22,
  -0.28, 3.42, -0.16,
  -0.38, 3.69, -0.09,
  -0.36, 3.78, -0.08,
  -0.54, 3.66, -0.11,
  -0.59, 3.35, -0.06,
  -0.16, 2.86, -0.03,
  0.21, 2.5, 0,
  0.53, 2.39, -0.01,
  0.57, 2.55, 0.02,
  0.69, 2.87, 0.04,
  0.76, 3.22, 0.06,
  0.67, 3.41, 0.08,
  0.31, 3.04, 0.09,
  0.17, 2.5, 0.03,
  0.28, 1.52, 0.04,
  0.51, 1.21, 0.08,
  0.82, 0.2, 0.03,
  1.37, -0.72, -0.03,
  1.75, -0.96, -0.11,
  1.8, -0.77, -0.15,
  1.61, -0.7, -0.09,
  1.47, _, -0.14,
  _, _, -0.07,
  -6.03, -4.41, -0.13,
  -5.77, -5.1, -0.1,
  -4.88, -5.06, -0.09,
  -4.26, -4.65, -0.12,
  -3.64, -4.45, 0.02,
  -3.14, -4.31, 0.05,
  -2.56, -3.62, 0.06,
  -2.25, -3.05, 0.13,
  -2.12, -2.82, 0.13,
  -2.04, -1.61, 0.17,
  -2.32, -1.9, 0.17,
  -2.53, -2.4, 0.2,
  -2.51, -1.78, 0.19,
  -2.57, -0.75, 0.2,
  -2.71, -0.42, 0.18,
  -2.81, -0.13, 0.15,
  -2.69, 0.13, 0.11,
  -2.66, 0.18, 0.06,
  -3.13, 0.19, -0.04,
  -3.52, 0.18, -0.05,
  -3.88, 0.14, -0.06,
  -4.13, -0.06, -0.14,
  -4.33, -0.56, -0.09,
  -4.47, -0.84, -0.16,
  -4.5, -1.36, 0,
  -4.23, -1.7, -0.17,
  -4.13, -1.88, -0.15,
  -3.63, -3.19, -0.32,
  -3.44, -3.27, -0.19,
  -3.13, -3.54, -0.19,
  -2.91, -3.86, -0.15,
  -2.72, -4.22, -0.12,
  -2.72, -4.55, 0.02,
  -2.12, -3.98, -0.12,
  -1.98, -3.94, -0.11,
  -1.86, -3.75, -0.03,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  -1.9, -3.9, -0.07,
  -1.91, -3.82, -0.07,
  -1.93, -3.69, -0.07,
  -2.04, -3.74, -0.07,
  -2.32, -3.67, -0.12,
  -2.77, -3.63, -0.13,
  -3.04, -3.56, -0.12,
  -3.51, -3.53, -0.06,
  -3.67, -3.65, -0.12,
  -3.65, -3.97, -0.04,
  -3.74, -4.01, 0,
  -4.09, -4.18, 0.06,
  -4.13, -4.39, 0.07,
  -4.37, -4.48, 0.06,
  -4.95, -4.46, _,
  -3.38, -3.91, -0.18,
  -2.96, -3.72, -0.12,
  -2.91, -3.67, -0.06,
  -2.77, -3.75, -0.09,
  -2.51, -3.7, 0.02,
  -2.18, -3.67, 0.04,
  -1.3, -3.76, 0.04,
  -0.92, -3.66, -0.02,
  -1.4, -4.59, 0.21,
  -1.48, -4.01, 0.24,
  -1.29, _, 0.07,
  -0.98, -2.56, -0.02,
  _, -2.5, -0.04,
  -4.26, -4.02, -0.21,
  -4.39, -5.33, -0.2,
  -2.75, -5.71, -0.54,
  -2.6, -5.38, -0.34,
  -2.16, -4.69, -0.21,
  -1.19, -4.76, -0.2,
  -0.81, -4.87, -0.3,
  -0.22, -4.37, -0.08,
  -0.48, -4.38, -0.13,
  -0.58, -4.64, -0.19,
  -0.97, -4.29, -0.14,
  -1.46, -3.09, -0.02,
  -2.06, -2.68, -0.21,
  -1.8, -2.42, -0.26,
  -1.73, -2.29, -0.12,
  -1.76, -2.19, -0.57,
  -2.04, -0.98, -0.54,
  -2.29, -0.66, -0.31,
  -2.1, -0.47, -0.72,
  -1.72, -0.39, -1.73,
  -1.26, -0.31, -1.58,
  -0.81, -0.55, -0.68,
  -0.69, -0.96, -0.06,
  -0.49, -1.24, -0.22,
  -0.47, -1.56, -0.22,
  -0.71, -2.3, -0.18,
  -0.72, -2.32, -0.09,
  -0.13, -2.29, 0.16,
  0.4, -2.62, 0.56,
  0.53, -2.74, 0.68,
  0.38, -2.74, 0.72,
  0, -2.88, 0.64,
  -0.28, -2.89, 0.6,
  -0.43, -3.04, 0.46,
  -0.46, -3.24, 0.37,
  -0.48, -3.39, 0.41,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  -0.37, -3.49, 0.34,
  -0.48, -3.7, 0.32,
  -0.63, -3.89, 0.25,
  -0.81, -4.02, 0.18,
  -0.98, -4.09, 0.15,
  -1.25, -4.11, 0.25,
  -1.55, -4.16, 0.02,
  -1.89, -4.33, -0.32,
  -1.87, -4.61, 0.01,
  -1.91, -4.67, _,
  _, -5.16, 3.2,
  _, -5.63, _,
  -1.63, -6.28, _,
  -0.67, -6.03, 0.67,
  -0.73, -6.19, -0.03,
  -0.53, -5.8, -0.29,
  -0.31, -5.43, 0.18,
  -0.03, -4.68, -0.3,
  -0.04, -3.43, -0.15,
  0.1, -2.8, -0.04,
  -0.98, -2.73, 0.09,
  -0.28, -3.99, _,
  0.22, -5.04, _,
  0.38, -4.99, 0.12,
  0.5, -4.96, 0.03,
  0.73, -4.46, -0.18,
  0.37, -2.22, _,
  _, -2.23, _,
  0.16, -2.72, -0.03,
  0.74, -2.77, 0.08,
  0.56, -2.98, 0.13,
  -0.07, -2.73, 0.1,
  -1.76, -2.24, 0.11,
  -2.78, -2.97, 0.08,
  -3.34, -3.85, 0.04,
  -4.33, -4.46, -0.02,
  -5.29, -4.77, -0.06,
  -5.84, -5.24, -0.13,
  -6.95, -5.19, -0.26,
  -7.75, -4.95, -0.39,
  -7.76, -5.39, -0.48,
  -7.75, -5.93, -0.58,
  -7.34, -6.18, -0.68,
  -7.26, -6.2, -0.63,
  -7.26, -6.95, -0.79,
  -7.55, -6.96, -0.7,
  -7.85, -7.38, -0.72,
  -8.21, -7.7, -0.81,
  -9.05, -8.01, -0.8,
  -8.99, -6.62, -0.78,
  -9.16, -7.29, -0.5,
  -9.54, _, -0.6,
  -9.28, _, -0.59,
  -9.78, _, 0.06,
  _, _, 0.13,
  _, _, _,
  -9.93, -7.77, -0.6,
  -10.24, _, -0.38,
  -10.86, -1.61, -1.67,
  -11.04, _, -0.31,
  -10.59, _, -0.64,
  -11.03, _, -0.34,
  -11.2, -6.35, -0.41,
  -11.15, -6.36, -0.39,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  -11.33, -6.64, -0.31,
  -11.65, -6.1, -0.01,
  -11.79, -5.89, -0.02,
  -11.68, -6.28, -0.02,
  -11.43, -6.64, -0.03,
  -11.03, -6.89, -0.04,
  -10.59, -6.94, -0.02,
  -10.36, -6.84, 0.04,
  -10.37, -6.77, 0.06,
  -10.4, -5.82, 0.19,
  -10.03, -5.95, 0.29,
  -8.7, _, 0.34,
  -7.88, _, 0.65,
  -7.54, -7.4, 0.01,
  -6.31, -5.73, -0.36,
  -5.71, -5.32, -0.29,
  -5.49, -4.8, -0.23,
  -5.38, -4.15, -0.23,
  -5.38, -3.75, -0.14,
  -5.23, -3.99, -0.25,
  -3.04, _, -0.22,
  -1.27, -1.43, -0.09,
  -0.99, -1.2, 0.21,
  -0.93, _, 0.12,
  -0.88, _, 0.05,
  _, _, 0.03,
  _, _, -0.14,
  -0.93, -1.55, -0.05,
  -5.97, -1.91, -0.12,
  -5.89, -2.98, -0.14,
  -5.32, -3.73, -0.19,
  -4.32, -3.79, -0.14,
  -3.89, -3.88, -0.12,
  -2.56, -3.43, -0.11,
  -1.43, -3.58, 0.04,
  -1.77, -3.67, 0.06,
  -1.99, -4.17, 0.02,
  -2.13, -4.42, 0.01,
  -1.89, -3.56, -0.01,
  -2.09, -2.23, 0.01,
  -1.86, -1.26, 0.08,
  -2.03, -0.64, 0.04,
  -2.48, -0.33, 0.06,
  -2.8, 0.21, 0.1,
  -2.83, 0.39, 0.13,
  -3.04, 0.38, 0.09,
  -3.09, 0.43, 0.09,
  -2.67, 0.51, 0.09,
  -2.38, 0.74, 0.09,
  -2.37, 0.68, 0.08,
  -2.52, 0.5, 0.05,
  -2.95, 0.22, 0.03,
  -3.43, -0.28, -0.05,
  -3.45, -0.28, -0.07,
  -3.38, -0.2, -0.09,
  -3.47, -0.39, -0.1,
  -3.49, -0.72, -0.06,
  -3.23, -1.22, -0.03,
  -3.05, -1.81, -0.11,
  -2.79, -2.49, -0.15,
  -3.04, -1.48, -0.07,
  -2.72, -2.56, -0.11,
  -2.45, -3.11, -0.06,
  -2.08, -3.25, 0.02,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  -2.06, -3.37, -0.05,
  -2.04, -3.5, -0.05,
  -2.01, -3.67, -0.07,
  -1.95, -3.91, -0.09,
  -1.9, -4.25, -0.1,
  -1.85, -4.4, -0.1,
  -1.83, -4.39, -0.09,
  -1.88, -4.29, -0.07,
  -1.89, -4.49, -0.06,
  -2.25, -4.83, -0.07,
  -2.4, _, -0.15,
  -2.66, -4.6, -0.18,
  -2.83, -4.77, -0.12,
  -2.96, -4.78, -0.11,
  -3.1, -4.63, -0.13,
  -3.4, -4.06, -0.08,
  -3.63, -3.47, -0.09,
  -3.71, -3.27, -0.08,
  -3.58, -3.22, -0.1,
  -3.37, -3.21, -0.1,
  -3.06, -3.02, -0.1,
  -2.56, -3.08, -0.1,
  -1.68, -3.7, -0.02,
  -0.97, -3.92, 0.02,
  -0.8, -3.79, 0.02,
  -0.57, -3.47, 0.02,
  -0.25, -2.49, -0.02,
  -0.25, -1.59, -0.03,
  -6.46, -4.69, -0.01,
  -4.5, -3.93, -0.02,
  -3.96, -7.15, 0,
  -3.87, -7.61, 0.01,
  -3.95, -7.73, -0.02,
  -3.47, -7.4, -0.15,
  -2.97, -7.51, -0.07,
  -2.81, -7.25, 0.01,
  -2.66, -6.55, 0.01,
  -2.83, -5.52, 0.01,
  -3.11, -5.1, -0.01,
  -3.68, -4.75, -0.01,
  -4.23, -4.04, 0,
  -4.56, -3.7, -0.01,
  -4.47, -3.48, -0.12,
  -4.61, -3.23, -0.16,
  -4.84, -2.87, -0.19,
  -4.94, -2.67, -0.22,
  -4.75, -2.6, -0.13,
  -4.31, -2.53, -0.02,
  -3.7, -2.53, 0.03,
  -3.55, -2.57, 0.01,
  -3.96, -2.77, 0.13,
  -4.8, -2.94, 0.21,
  -5.41, -3.2, 0.18,
  -5.37, -3.42, 0.17,
  -5.12, -3.71, 0.26,
  -4.63, -4.04, 0.13,
  -4.24, -4.41, 0.19,
  -4.18, -4.88, 0.19,
  -3.95, -5.03, 0.08,
  -3.48, -5.3, 0.15,
  -3.34, -5.82, 0.21,
  -3.63, -5.88, 0.33,
  -3.99, -5.72, 0.3,
  -4.34, -5.82, 0.38,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  -4.65, -5.88, 0.44,
  -4.9, -5.97, 0.42,
  -4.99, -6.15, 0.39,
  -5.26, -6.5, 0.33,
  -5.34, -6.91, 0.28,
  -5.36, -7.24, 0.24,
  -5.46, -7.7, 0.17,
  -5.39, -8.17, 0.16,
  -5.25, -8.48, 0.13,
  -5.35, -8.61, 0.32,
  -5.4, _, 0.52,
  -4.22, -8.37, 0.42,
  -3.89, -8.06, 0.22,
  -2.89, -7.67, 0.15,
  -2.83, -7.27, 0.12,
  -2.78, -6.88, 0.04,
  -2.87, -6.55, -0.02,
  -2.95, -6.14, -0.03,
  -2.9, -5.48, -0.04,
  -3.2, -4.55, -0.4,
  -2.12, -4.33, -0.15,
  -3.59, -4.93, -0.39,
  -2.02, -5.15, 0.26,
  -0.46, -5.19, 0.31,
  -1.21, -5.1, 0.17,
  -1.71, -4.37, 0.14,
  -1.81, -3.64, 0.03,
  -1.8, -3.29, -0.03,
  -0.29, -0.03, -0.09,
  -0.34, -0.15, -0.06,
  -0.32, -0.22, -0.08,
  -0.33, -0.9, -0.09,
  -0.2, -1.07, -0.07,
  -0.15, -0.92, -0.06,
  -0.21, -0.84, -0.03,
  -0.23, -0.71, -0.15,
  -0.36, -1.18, -0.41,
  -0.07, -1.3, -0.42,
  0.58, -0.96, 0.02,
  0.49, -1.36, 0.14,
  0.4, -2.02, 0.16,
  0.02, -5.19, 0.19,
  0.2, -5.36, 0.09,
  0.38, -5.49, 0.01,
  0.5, 0.81, 0.04,
  0.28, 1.65, 0.04,
  0.17, 2.23, 0.03,
  0.09, -3.59, 0.02,
  0.15, -4.25, 0.14,
  0.2, _, 0.16,
  -0.27, 0.1, 0.04,
  -0.23, 0.16, 0.06,
  0.19, 0.17, 0.07,
  0.4, -0.06, 0.04,
  0.78, 6.79, 0.01,
  0.53, 0.11, -0.02,
  0.82, -0.21, -0.03,
  1.09, -0.15, -0.04,
  1.17, 0.33, -0.13,
  0.94, 0.05, -0.03,
  1, 0.05, -0.06,
  1.01, 0.27, -0.05,
  0.95, 0.18, -0.05,
  0.95, 0.04, -0.04,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0.98, 0.02, -0.02,
  1.14, -0.03, -0.03,
  1.39, -0.07, 0.01,
  1.48, 2.34, 0.11,
  1.73, 8.69, 0.32,
  1.69, 8.58, 0.24,
  1.93, 8.69, 0.05,
  1.58, 8.69, 0,
  2.24, 8.3, 0.13,
  1.88, 8.68, _,
  2.02, 8.73, _,
  _, 8.71, _,
  1.1, 8.9, 0,
  _, 8.43, 0.05,
  _, 8.44, 0.23,
  _, 8.47, 0.2,
  2.8, 8.78, _,
  2.78, 8.49, 0.26,
  _, 8.65, 0.24,
  _, 8.81, 0.04,
  2.38, 8.72, -0.03,
  2.29, 8.78, -0.08,
  2.21, 8.81, 0.07,
  2.09, 9.08, -0.04,
  1.93, 9, -0.01,
  0.92, _, -0.01,
  0.52, 8.99, 0.03,
  0.2, _, 0.07,
  2.58, 0.13, -0.03,
  1.13, 1.29, 0.05,
  1.15, 0.93, 0.03,
  0.37, 1.08, 0.01,
  -0.01, 0.81, 0.04,
  -0.53, 0.31, -0.04,
  -1.35, -0.04, -0.05,
  -2.13, -0.45, -0.16,
  -2.86, -1.21, -0.12,
  -3.32, -1.88, -0.2,
  -3.65, -2.68, -0.31,
  -4.08, -3.56, -0.18,
  -4.63, -4.68, -0.19,
  -5.27, -5.47, -0.54,
  -6.19, -5.61, -0.12,
  -6.28, -5.12, -0.18,
  -6.02, -4.75, -0.04,
  -6.28, -5.04, -0.06,
  -6.44, -5.29, 0.08,
  -0.14, -5.33, -0.03,
  0.06, -5.11, -0.01,
  _, -5.06, 0,
  _, -4.89, _,
  _, _, _,
  -15.21, _, _,
  -5.71, _, _,
  _, -5.5, _,
  _, _, _,
  -26.71, -5.81, 0.23,
  -6.73, -6.19, 0.46,
  -6.24, -6.36, 0.02,
  -6.69, -6.23, _,
  -7.16, -6.4, 0.18,
  -7.71, -6.49, _,
  -8.19, -5.44, _,
  -9.17, -5.24, 0.57,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  -9.57, -5.08, 1.15,
  -9.89, -4.94, 0.39,
  -10.6, -4.8, 0.79,
  -10.83, -4.58, 0.62,
  -11.26, -4.8, 0.54,
  _, -13.57, _,
  -12.47, -5.9, _,
  -11.57, -6.38, 0.19,
  -10.73, -6.69, -0.06,
  -10.8, -6.68, _,
  _, -6.6, _,
  _, -6.85, _,
  _, -6.85, _,
  _, -6.84, _,
  -3.8, -5.34, 0.33,
  -3.81, -4.71, 0.04,
  -3.93, -4.43, 0.07,
  -4.13, -4.27, -0.1,
  -4.05, -3.87, 0.08,
  -4.11, -3.08, _,
  -4.54, -1.47, _,
  -4.69, -1.37, _,
  -4.71, -1.44, 0.58,
  -4.36, -1.59, _,
  _, -2.16, _,
  _, _, _,
  -3.25, -1.3, _,
  _, -1.3, _,
  -3.16, -4.2, -0.14,
  -2.89, -3.42, -0.1,
  -3.23, -3.41, -0.04,
  -3.8, -3.54, -0.07,
  -3.9, -3.71, -0.11,
  -3.84, -3.94, -0.14,
  -3.5, -4.19, -0.14,
  -3.64, -4.05, -0.26,
  -3.59, -3.83, -0.41,
  -3.37, -3.55, -0.32,
  -3.28, -3.34, -0.15,
  -3.08, -3.03, -0.14,
  -3.1, -3.27, -0.15,
  -2.96, -3.08, -0.21,
  -2.95, -0.75, -0.23,
  -3.42, 0.75, -0.2,
  -3.54, 1.17, -0.23,
  -3.25, 1.08, -0.3,
  -3.41, 0.53, -0.11,
  -3.75, 0.52, -0.15,
  -3.9, 0.5, 0.02,
  -3.93, 0.38, -0.01,
  -4.03, _, -0.07,
  -4.28, -0.15, 0.1,
  -4.26, -0.29, 0.04,
  -4.1, -0.32, 0,
  -3.96, _, 0.29,
  _, _, _,
  -3.78, -0.86, 0.07,
  -3.81, -0.77, 0.05,
  -3.66, -0.65, 0.13,
  -3.08, -0.81, -0.11,
  -3.3, -0.7, 0.02,
  -3.01, -0.83, -0.04,
  -1.78, -1.13, 0.1,
  -1.83, -1.67, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, -1.24, -0.07,
  _, _, _,
  _, -2.03, _,
  _, -2.28, _,
  -3.31, -2.09, 0.08,
  -3.17, -2.29, -0.15,
  -3.22, -2.15, -0.21,
  -2.65, -1.49, -0.19,
  _, _, -0.01,
  _, _, _,
  _, _, _,
  9.29, _, _,
  9.46, _, _,
  8.62, -1.68, _,
  -3.41, -1.36, -0.04,
  -3.43, -1.83, _,
  _, -2.15, -0.06,
  _, -2.22, _,
  _, -1.79, -0.16,
  _, -1.74, -0.13,
  6.73, -2.38, 0.19,
  _, _, 0.09,
  _, -2.12, _,
  _, _, _,
  15.22, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  -4.7, -3.12, 0.06,
  -4.31, -4.88, 0.08,
  -3.5, -4.57, 0.09,
  -2.71, -4.01, 0.07,
  -2.09, -4.2, 0.08,
  -1.04, -4.5, 0.08,
  -0.7, -4.44, 0.05,
  -0.93, -2.98, 0.05,
  -1.94, -2.56, 0.04,
  -2.46, -2.75, 0.03,
  -2.68, -3.32, 0.04,
  -2.63, -3.45, 0.05,
  -2.47, -3.37, 0.04,
  -2.31, -3.14, 0.09,
  -2.09, -2.4, 0.04,
  -2.19, -2.3, 0.05,
  -2.23, -2.28, 0.09,
  -2.11, -2.28, 0.1,
  -1.53, -2.37, 0.07,
  -0.9, -2.51, 0.1,
  -0.48, -2.82, 0.12,
  -0.41, -3.12, 0.08,
  -0.44, -3.37, 0.08,
  -0.17, -3.54, 0.07,
  -0.19, -3.53, 0.06,
  -0.03, -3.77, 0.07,
  -0.01, -4.03, 0.07,
  -0.15, -4.31, 0.03,
  -0.47, -4.48, 0,
  -0.57, -4.58, 0,
  -0.37, -4.39, -0.02,
  -0.19, -4.44, -0.02,
  -0.29, -4.25, 0.11,
  -0.35, -4.27, 0.07,
  -0.74, -4.59, 0.1,
  -1.1, -4.75, 0.19,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  -0.84, -4.65, 0.05,
  -0.9, -4.68, 0.07,
  -0.71, -4.65, 0.1,
  -0.8, -4.6, 0.13,
  -0.91, -4.61, 0.12,
  -1.27, -4.77, 0.12,
  -1.45, -5.2, 0.16,
  -1.69, -5.61, 0.13,
  -1.75, -6.21, 0.14,
  -1.78, -6.86, 0.11,
  -1.97, -7.12, 0.18,
  -1.9, -8.47, 0.04,
  -2.06, -8.72, 0.19,
  -1.98, -8.88, 0.07,
  -1.65, -8.81, 0.19,
  -1.07, -7.36, 0.14,
  -0.64, -6.01, 0.19,
  -0.62, -5.23, 0.19,
  -0.65, -4.81, 0.12,
  -0.74, -4.35, 0.06,
  -0.89, -4.15, 0,
  -0.77, -4.68, -0.1,
  -0.57, -4.66, -0.12,
  -0.37, -4.28, -0.07,
  -0.18, -3.86, -0.05,
  -0.06, -3.51, 0.11,
  0.2, -2.53, 0.14,
  0.21, -1.45, 0.11,
  -4.19, -3.12, 0.05,
  -4.78, -3.15, 0.02,
  -5.15, -3.28, -0.16,
  -2.86, -4.22, -0.03,
  -3, -4.23, -0.14,
  -1.92, -4.32, -0.14,
  -1.32, -3.98, -0.05,
  -1.2, -3.65, 0.09,
  -0.87, -3.43, 0.13,
  -0.62, -3.25, 0.08,
  -0.41, -2.99, 0.12,
  -0.56, -2.95, 0.19,
  -0.55, -2.27, 0.26,
  -0.64, -1.9, 0.32,
  -1.3, -1.65, 0.44,
  -1.18, -1.02, 0.48,
  -0.98, -0.99, 0.51,
  -1.28, -2.17, 0.55,
  -0.34, -2.64, 0.78,
  -0.32, -3.14, 1.04,
  -0.61, -3.43, 1.05,
  -0.82, -3.57, 1.1,
  -1.35, -3.4, 1.13,
  -1.79, -3.44, 1.16,
  -2.05, -3.9, 1.17,
  -2.92, -4.15, 1.09,
  -3.45, -4.47, 1.16,
  _, _, _,
  -2.7, -3.82, 1.03,
  -1.88, -3.75, 1.02,
  -5.36, -3.74, 1.1,
  -6.38, -4.69, 0.96,
  -5.97, -3.92, 0.91,
  -5.95, -4.01, 0.99,
  -6.52, -3.84, 0.82,
  -6.84, -3.76, 0.98,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  -6.63, -3.65, 0.74,
  -6.79, -3.5, 0.66,
  -6.8, -3.41, 0.61,
  -6.8, -3.35, 0.56,
  -6.9, -3.82, 0.54,
  -7.02, -3.63, 0.39,
  -6.9, -3.98, 0.24,
  -6.75, -4.33, 0.06,
  -6.36, -4.38, _,
  -6.27, -5.16, -0.1,
  -5.99, -5.35, -0.11,
  -5.61, _, -0.16,
  -4.95, _, -0.18,
  -4.06, _, -0.19,
  -4.05, -7.21, -0.18,
  -3.95, -7.06, -0.25,
  -3.62, -6.49, -0.37,
  -3.38, -6.36, -0.38,
  -3.37, -5.96, -0.36,
  -3.33, -5.59, -0.38,
  -3.55, -4.47, -0.37,
  -3.65, -4.05, -0.46,
  -4.24, -3.56, _,
  -4.69, _, _,
  -4.89, _, -0.23,
  -3.6, -4.07, -0.25,
  -3.32, -2.83, -0.05,
  -3, -2.61, -0.02,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  -4.76, _, 0,
  -5.38, 0.41, 0,
  -4.84, -6.35, 0.01,
  -5.38, -7.49, -0.01,
  -1.27, _, -0.64,
  -3.65, -6.99, -0.41,
  -4.39, -7.11, -0.35,
  -4.11, -6.86, -0.28,
  -4.23, -6.29, -0.38,
  -4.11, -5.87, -0.16,
  -3.67, -5.61, -0.17,
  -3.82, -5.62, -0.16,
  -3.46, -5.55, -0.12,
  -3.02, -5.45, -0.16,
  -2.93, -5.11, -0.1,
  -2.73, -4.85, 0.14,
  -2.71, -4.54, 0.33,
  -2.87, -4.36, 0.55,
  -2.75, -5.11, 0.64,
  -2.63, -4.33, 0.54,
  -3.69, -4.7, 0.45,
  -2.72, -4.25, 0.49,
  -3, -4.35, 0.65,
  -3.08, -3.93, 0.64,
  -3.74, -3.83, 1.63,
  -4.09, -3.7, 1.87,
  -3.96, -3.76, 1.27,
  -2.69, -4.22, 0.67,
  -2.48, -4.32, 0.56,
  -2.31, -4.3, 0.42,
  -2.37, -4.27, 0.66,
  -0.17, -4.68, 0.92,
  -2.52, -4.31, 0.67,
  9.83, -4.91, 0.76,
  9.78, -4.72, 1.08,
  -3.03, -4.31, 0.73,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  -3.18, -4.48, 0.85,
  -3.06, -5.04, 0.74,
  -3.16, -5.19, 0.56,
  -3.48, -6.78, 0.44,
  -3.51, -8.35, 0.28,
  -3.79, -10.1, 0.19,
  -3.64, -10.75, 0.11,
  -3.73, -11.2, 0.07,
  -4.03, _, 0.06,
  -4.11, _, 0.01,
  -3.39, -10.36, 0.04,
  -2.03, -10.36, -0.06,
  -1.31, -10.12, -0.2,
  -0.94, -9.19, -0.31,
  -0.68, -8.78, -0.31,
  -0.43, -8.35, -0.3,
  -0.23, -7.64, -0.28,
  -0.09, -7.57, -0.24,
  -0.22, -5.63, -0.22,
  -0.81, -4.68, -0.12,
  -0.99, -4.78, -0.06,
  -0.86, -4.76, -0.13,
  -0.53, -4.43, -0.13,
  -0.3, -3.85, -0.1,
  -0.12, -3.11, -0.16,
  _, -2.64, -0.08,
  -1.23, _, 0.01,
  -2.66, _, _,
  -2.53, -0.42, -0.08,
  -1.72, -0.53, -0.08,
  -1.26, -1.07, -0.11,
  -0.92, -1.91, -0.07,
  -0.46, -2.13, -0.07,
  -0.18, -2.55, -0.07,
  0.55, -2.07, 0.21,
  0.61, -1.85, 0.05,
  0.89, -1.49, 0.12,
  0.91, -1.25, 0.2,
  1.65, -0.95, 1.14,
  1.48, -0.13, -0.02,
  1.62, 0.02, -0.06,
  3.25, 0.04, 2.74,
  2.25, -0.7, 1.6,
  1.71, -0.73, 0.42,
  1.53, -0.53, 0.66,
  1.01, -0.73, 0.49,
  1.69, -0.95, 0.29,
  2.09, -0.83, 0.14,
  2.03, -0.92, 0.16,
  1.71, -1.14, 0.17,
  1.93, -1.09, 0.05,
  2.21, -1.12, 0.22,
  2.37, -1.58, 0.12,
  2.64, -1.7, 0.1,
  2.47, -1.89, 0.09,
  2.75, -1.03, 0.59,
  3.05, -1.33, 0.1,
  3.53, -2.35, -0.16,
  3.9, -2.49, 0.16,
  3.51, -2.5, -0.03,
  3.73, -2.95, 0.03,
  3.77, -3.25, -0.11,
  4.09, -3.46, 0.22,
  3.98, -2.72, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, 0.11,
  _, -3.14, -0.61,
  _, _, -0.01,
  _, -3.51, -0.17,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, -17.06, _,
  _, _, _,
  _, _, _,
  _, _, 1.45,
  _, _, _,
  _, _, _,
  _, -2.81, _,
  _, -2.41, _,
  3.81, -1.85, _,
  3.87, _, _,
  4.24, _, _,
  3.73, _, _,
  _, _, _,
  _, _, _,
  18.67, _, _,
  0.81, _, _,
  0.95, _, _,
  1.4, 12.49, _,
  -0.41, -0.19, -0.01,
  -1.66, -0.19, 0.02,
  -1.87, 0.4, 0.05,
  -2.14, 0.69, 0.04,
  -2, 0.71, 0.05,
  -2.13, 0.73, 0.07,
  -2.27, 0.56, 0.13,
  -2.35, -0.07, 0.11,
  -2.33, 0.66, 0.34,
  -2.25, 3.5, 0.03,
  -7.03, 2.03, 0.01,
  -3.19, 2.22, -0.01,
  -2.81, 0.75, -0.04,
  -2.24, 0.64, -0.01,
  -1.59, 0.82, 0.03,
  -0.96, 0.98, 0.04,
  -0.87, 1.25, -0.04,
  -0.7, 1.4, 0,
  -0.18, 0.88, -0.02,
  -0.11, 1.51, -0.08,
  -0.32, _, -0.07,
  _, _, 0,
  _, _, -0.06,
  _, 2.39, -0.04,
  _, _, -0.05,
  _, _, 0.01,
  _, _, -0.04,
  _, _, 0.01,
  _, _, -0.01,
  _, _, 0.03,
  -2.68, 10.63, 0,
  -2.53, 2.63, 0,
  -2.55, 1.94, -0.34,
  -2.23, 2.38, -0.17,
  -1.73, 2.84, -0.22,
  -1.23, 3.09, -0.15,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  -1.48, 2.61, -0.1,
  -1.68, 2.84, -0.16,
  -2.13, 2.96, -0.06,
  _, _, -0.01,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, -0.15,
  _, _, _,
  _, _, -3.55,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  -2.26, -1.46, 0.06,
  -1.85, -1.98, -0.02,
  -1.87, -2.34, -0.05,
  -2.2, -2.52, -0.07,
  -2.34, -2.42, -0.08,
  -2.36, -2.42, -0.17,
  -2.19, -2.26, -0.1,
  -1.82, -2.19, -0.09,
  -1.49, -2.08, -0.12,
  -1.53, -2.21, 0,
  -1.38, -2.35, -0.02,
  -1.17, -2.56, -0.08,
  -0.79, -2.85, 0.06,
  -0.7, -3.14, 0.1,
  -0.68, -3.22, 0.06,
  -1.12, -3.44, 0.09,
  -1.42, -3.63, 0.08,
  -2, -3.74, 0.07,
  -2.62, -3.66, 0.16,
  -2.57, -3.23, 0.15,
  -2.71, -3.54, 0.24,
  -2.99, -3.49, 0.14,
  -3.2, -3.38, 0.17,
  -3.06, -3.54, 0.13,
  -2.87, -3.84, 0.2,
  -3.77, -4.38, 0.14,
  -4.09, -4.87, 0.07,
  -4.63, _, _,
  -4.33, -4.63, 0.1,
  -4.94, -4.67, 0.1,
  -5.76, -4.76, 0.04,
  -6.41, -4.84, 0.03,
  -6.71, -4.58, -0.02,
  -6.87, -4.45, -0.03,
  -6.84, -4.33, 0.05,
  -6.76, -4.57, -0.1,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  -6.78, -4.62, -0.13,
  -6.7, -4.76, -0.17,
  -6.41, -5.05, -0.13,
  -6.64, -5.4, 0.01,
  -6.24, -5.48, 0.09,
  -6.17, _, _,
  -5.86, _, -0.1,
  _, -6.77, -0.17,
  _, -6.77, -0.01,
  _, _, -0.05,
  _, _, _,
  _, _, 0.08,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  -2.04, -7.54, _,
  -2.08, -7.44, 0.32,
  -2.05, -7.28, 0.58,
  -2.23, -6.92, 0.46,
  -2.15, -6.87, 0.31,
  -1.9, -6.4, 0.34,
  -3.56, _, 0.26,
  _, _, -0.01,
  _, _, -0.09,
  -2.53, _, 0.14,
  -2.44, -3.48, -0.04,
  -2.91, -2.91, -0.02 ;

 specWidth =
  2.2801, 1.96, 0.0361,
  1, 0.8836, 0.1024,
  0.36, 0.3025, 0.1024,
  0.3969, 0.2704, 0.0676,
  0.2304, 0.2025, 0.0729,
  0.16, 0.2601, 0.1296,
  0.1521, 0.36, 0.1521,
  0.3969, 0.2704, 0.1444,
  0.7225, 0.2304, 0.16,
  0.4489, 0.2025, 0.1296,
  0.3364, 0.2116, 0.1296,
  0.2809, 0.2025, 0.1369,
  0.3249, 0.25, 0.1369,
  0.2916, 0.1764, 0.1089,
  0.2209, 0.1089, 0.09,
  0.25, 0.1369, 0.09,
  0.2401, 0.1764, 0.0841,
  0.2916, 0.0729, 0.0784,
  0.2304, 0.0784, 0.0841,
  0.2116, 0.0729, 0.0784,
  0.2304, 0.0961, 0.0784,
  0.3844, 0.0961, 0.1024,
  0.4096, 0.09, 0.1024,
  0.4761, 0.09, 0.1156,
  0.5041, 0.1225, 0.1156,
  0.3969, 0.1444, 0.1681,
  0.2916, 0.1681, 0.1521,
  0.2116, 0.1936, 0.1849,
  0.4624, 0.2116, 0.2116,
  0.4489, 0.4624, 0.2025,
  0.3481, 0.3025, 0.2401,
  0.3969, 0.2025, 0.2025,
  0.4489, 0.2025, 0.2209,
  0.4489, 0.3969, 0.2025,
  0.4096, 0.2704, 0.3025,
  0.5929, 0.2809, 0.2916,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  1.44, 0.4489, 0.1681,
  1.4884, 0.5476, 0.1936,
  0.9604, 0.6084, 0.2209,
  0.7569, 0.7396, 0.2809,
  0.7569, 0.8281, 0.36,
  0.8649, 0.6084, 0.4096,
  0.7396, 0.64, 0.3844,
  1.1236, 0.4761, 0.4096,
  0.7569, 0.5929, 0.4096,
  0.6561, 0.7056, 0.4356,
  1.0201, 0.9409, 0.3969,
  1.0201, 1.1664, 0.3969,
  0.6724, 1.1449, 0.3364,
  0.8464, 0.7921, 0.4096,
  0.9409, 1.1025, 0.4225,
  1, 0.9216, 0.3721,
  1.1449, 1.5129, 0.3481,
  1.0609, 1.7424, 0.2809,
  1.9321, 1.8496, 0.2704,
  1.3689, 1.3924, 0.25,
  0.8649, 1.0609, 0.1764,
  0.6889, 0.9216, 0.16,
  0.64, 0.8464, 0.1521,
  0.7569, 0.6084, 0.1369,
  _, 0.64, 0.1764,
  _, 0.9025, 0.2025,
  0.2916, 1.0201, 0.2304,
  _, 0.5476, 0.2025,
  3.0625, 7.7841, 39.9424,
  0.9604, 4.3264, 2.2201,
  1.7161, _, 1.7424,
  0.7056, 2.6244, 0.6724,
  0.7921, 3.2041, 0.5041,
  0.9801, 3.2041, _,
  0.9801, 1.7161, _,
  1.2321, 0.9604, 0.2916,
  1.4884, 0.5625, 0.25,
  1.5625, 0.4225, 0.16,
  _, _, 0.2401,
  _, 0.81, 0.3249,
  0.5184, 0.8836, 0.2809,
  0.6561, 0.8649, 0.0841,
  0.5625, 0.9409, 0.16,
  0.5625, 1.44, 0.1764,
  0.5929, 1.7161, 0.1681,
  0.6241, 0.3136, 0.2116,
  0.6724, 0.3364, 0.2209,
  0.4761, 4.3681, 0.2116,
  0.7921, 0.8281, 0.2304,
  0.7921, 0.7056, 0.2209,
  0.7225, 0.6241, 0.3136,
  0.6561, 0.1225, 0.1444,
  0.5476, 0.1156, 0.1024,
  _, _, _,
  _, _, _,
  _, _, _,
  _, 0.2916, 0.1936,
  _, 0.3364, 0.1764,
  _, 0.5329, 0.1681,
  _, 0.4624, 0.2116,
  _, 0.3249, 0.1444,
  _, 0.25, 0.1849,
  _, _, 0.25,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, 0.2401,
  _, _, 0.1764,
  _, _, 0.1369,
  _, _, 0.1156,
  _, _, 0.1089,
  _, _, _,
  _, _, 0.0784,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, 0.0841,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, 0.1521,
  _, _, 0.1024,
  _, 1.2996, 0.1089,
  _, _, 0.0784,
  _, _, 0.1369,
  _, _, 0.1089,
  0.2916, 0.2209, 0.1296,
  0.49, 0.2209, 0.1444,
  0.6724, 0.36, 0.1764,
  0.5329, 0.2401, 0.1681,
  0.3025, 0.2116, 0.1849,
  0.3721, 0.1936, 0.1764,
  0.4761, 0.2304, 0.1681,
  0.5329, 0.4096, 0.2809,
  0.5625, 0.2116, 0.1849,
  0.36, 0.1369, 0.5476,
  0.2809, 0.0961, 0.1521,
  0.2304, 0.2704, 0.1369,
  0.4489, 0.1296, 0.0961,
  0.4225, 0.0676, 0.0841,
  0.3844, 0.0625, 0.09,
  0.2916, 0.1089, 0.0841,
  0.16, 0.1521, 0.1521,
  0.1156, 0.2304, 0.0961,
  0.3249, 0.2809, 0.0625,
  0.3136, 0.2304, 0.0625,
  0.2916, 0.3025, 0.0841,
  0.2209, 0.2401, 0.1089,
  0.3025, 0.2401, 0.1156,
  0.25, 0.16, 0.0841,
  0.4761, 0.1849, 0.1024,
  0.2304, 0.2916, 0.0729,
  0.2401, 0.3969, 0.1089,
  0.1444, 0.36, 0.1296,
  0.3249, 0.3136, 0.0676,
  0.3136, 0.3249, 0.0729,
  0.2401, 0.3364, 0.0729,
  0.2209, 0.4225, 0.0841,
  0.2401, 0.6889, 0.09,
  0.16, 0.1764, 0.2916,
  0.2304, 0.2304, 0.1681,
  0.2116, 0.1936, 0.1024,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0.3721, 0.4356, 0.1444,
  0.5625, 0.5184, 0.1296,
  0.3844, 0.64, 0.1369,
  0.8649, 0.6084, 0.1156,
  _, 0.2916, 0.1849,
  _, 0.8649, 0.2025,
  _, 0.2704, 0.2601,
  0.6561, 0.3136, 0.1764,
  0.81, 0.3025, 0.1936,
  _, _, 0.36,
  _, _, 0.5476,
  0.1764, _, _,
  _, _, 0.1444,
  _, 0.2704, 0.16,
  _, 0.4096, _,
  _, 0.6561, 0.1444,
  0.9409, 0.7921, 0.2809,
  0.5776, 1.0816, 0.2401,
  0.49, 1.1236, 0.2916,
  0.5476, 0.64, 0.16,
  0.6561, 0.5476, 0.2401,
  _, 0.7744, 0.2116,
  _, _, 0.25,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, 0.0361,
  0.4761, 3.2041, 0.3249,
  0.7225, 1.2996, 0.2704,
  0.7056, 1.1025, 0.3025,
  0.2401, 0.7225, 0.2704,
  0.2916, 0.9216, 0.1936,
  0.4225, 1.4641, 0.16,
  0.2704, 0.7744, 0.0961,
  0.2401, 0.7396, 0.0841,
  0.1521, 0.7225, 0.0961,
  0.1296, 0.6561, 0.1089,
  0.1225, 0.7396, 0.1156,
  0.1089, 1.4161, 0.1089,
  0.2304, 1.44, 0.0729,
  0.1936, 0.5329, 0.0576,
  0.2601, 0.5476, 0.0729,
  0.3844, 0.3249, 0.0729,
  0.1521, 0.3481, 0.0729,
  0.2025, _, 0.0841,
  0.25, 0.5041, 0.1024,
  0.1681, _, 0.1296,
  0.1764, _, 0.25,
  _, _, _,
  _, _, _,
  _, _, _,
  0.2116, _, 0.1024,
  0.2116, 0.4761, 0.0841,
  0.2116, _, 0.1369,
  0.09, _, 0.0729,
  0.25, 0.4225, 0.1089,
  0.2704, 1.2769, 0.0961,
  0.3136, 0.4489, 0.1296,
  0.3481, 0.3969, 0.1444,
  0.4356, 0.3721, 0.1444,
  0.5329, 0.4624, 0.1225,
  0.5929, 0.5476, 0.1296,
  0.3969, 0.4489, 0.1225,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0.5329, 0.4489, 0.0961,
  1.1025, 0.4624, 0.1089,
  2.56, 0.6241, 0.1296,
  3.1684, _, 0.2025,
  0.5776, _, 0.25,
  0.7056, 0.5041, 0.1849,
  0.9409, 0.5184, 0.2025,
  0.9604, 0.4225, 0.1764,
  0.8649, 0.49, 0.16,
  0.5041, 0.64, 0.16,
  0.5184, 0.9409, 0.2116,
  0.3136, 0.7744, 0.1024,
  0.6889, _, _,
  0.6084, _, 0.2809,
  0.3969, _, 0.2304,
  0.5184, _, 0.25,
  0.7921, _, 0.1936,
  4.4521, _, 0.2601,
  3.4225, _, 0.2809,
  2.2801, 1.4884, 0.2601,
  0.9216, _, 0.2209,
  1.7956, _, 0.2304,
  0.8649, _, 0.1936,
  0.9216, _, 0.16,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0.8464, 15.7609, 0.5041,
  1.0816, 3.6481, 0.5476,
  5.29, 1.4161, 0.3969,
  1.1881, 2.9241, 0.1849,
  0.7396, 1.69, 0.1849,
  0.3721, 0.7056, 0.1764,
  0.3249, 0.4761, 0.1936,
  0.2601, 0.3136, 0.2025,
  0.3136, 0.2916, 0.2304,
  0.2304, 0.3364, 0.3025,
  0.3249, 0.3969, 0.4225,
  0.5625, 0.5184, 0.5329,
  0.5184, 0.5041, 0.64,
  0.6561, 0.4761, 0.6241,
  0.9604, 0.5184, 0.6241,
  1.0816, 0.5776, 0.7396,
  1.0404, 0.6724, 0.7225,
  0.6889, 0.8464, 0.8281,
  0.8281, 0.8649, 0.6724,
  0.7569, 0.5041, 0.5929,
  0.7396, 0.5184, 0.5929,
  0.7921, 0.5476, 0.6561,
  0.8836, 0.5329, 0.7056,
  0.7396, 0.5776, 0.6561,
  0.64, 0.6084, 0.5929,
  0.7225, 0.5184, 0.4761,
  0.6241, 0.5041, 0.4225,
  0.5041, 0.4096, 0.3364,
  0.3721, 0.3364, 0.2601,
  0.2601, 0.3249, 0.2601,
  0.2704, 0.3481, 0.2401,
  0.2916, 0.3025, 0.2601,
  0.36, 0.2916, 0.2401,
  0.3969, 0.2916, 0.2704,
  0.3364, 0.2704, 0.3025,
  0.3249, 0.2809, 0.25,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0.5184, 0.6889, 0.3249,
  0.4096, 0.8836, 0.3249,
  0.3844, 0.7396, 0.3136,
  0.5184, 0.9604, 0.3481,
  0.81, 1, 0.3025,
  1.0816, 0.7056, 0.3249,
  1.4884, 0.64, 0.36,
  1.2321, 1.0404, 0.3481,
  1, 1.3456, 0.3721,
  0.7056, 1, 0.4624,
  0.8649, 1.0404, 0.5625,
  0.7921, 1.6641, 0.5776,
  1.21, 1.6384, 0.5776,
  1.9044, 1.1025, 0.6561,
  1.9321, 1.44, 0.6241,
  1.8225, 2.1609, 0.5625,
  1.5129, 2.6244, 0.4489,
  1.3456, 2.7556, 0.3969,
  1.1664, 2.4649, 0.3364,
  1.0609, 1.8496, 0.3844,
  0.8464, 1.0201, 0.3136,
  1.2769, 1.2544, 0.2916,
  1.2321, 1.5876, 0.2601,
  1.1025, 0.8836, 0.2401,
  1.1664, 0.5929, 0.16,
  1.1881, 0.6561, 0.1681,
  1.1881, 1.3225, 0.2601,
  _, 1.0816, 0.2809,
  1.2769, 6.6049, 0.6561,
  2.5921, 2.7225, 0.5476,
  1.7689, 0.8281, 0.9409,
  1.6129, 0.8281, 1.21,
  1.4641, 0.6889, 1.3689,
  2.1316, 0.6889, 0.7225,
  0.7056, 0.2704, 0.3364,
  0.3136, 0.3481, 0.1764,
  0.1296, 0.2916, 0.1444,
  0.0961, 0.1089, 0.1681,
  0.1296, 0.1521, 0.1369,
  0.2025, 0.1681, 0.25,
  0.2209, 0.2025, 0.2116,
  0.1849, 0.1849, 0.1681,
  0.16, 0.1444, 0.2116,
  0.2916, 0.1764, 0.16,
  0.2304, 0.1764, 0.1521,
  0.2401, 0.1369, 0.1681,
  0.2916, 0.1764, 0.1849,
  0.1681, 0.2704, 0.1521,
  0.1681, 0.1521, 0.2025,
  0.1936, 0.1764, 0.1444,
  0.1849, 0.2116, 0.1681,
  0.2209, 0.2304, 0.2209,
  0.2401, 0.25, 0.2916,
  0.2209, 0.2401, 0.2025,
  0.2209, 0.3721, 0.2209,
  0.2916, 0.6084, _,
  1.0609, 1.2996, 0.3025,
  2.1904, 1.2544, 0.3481,
  0.6889, 0.8281, 0.4356,
  1.1449, 1.3225, 0.5184,
  0.4356, 0.4761, 0.2401,
  0.4356, 0.7744, 0.3844,
  0.6889, 1.1025, 0.49,
  0.7921, 0.7396, 0.6241,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  1.0404, 1.3225, 0.8464,
  1.0201, 1.1881, 0.81,
  0.8649, 1.1664, 0.7569,
  1.0404, 0.8836, 0.64,
  0.8836, 1.0816, 0.6084,
  0.8836, 1.0816, 0.5625,
  1.1449, 1.1449, 0.5184,
  0.4096, 0.9216, 0.6889,
  0.2401, 0.8281, 0.3844,
  _, 1.2321, _,
  0.4096, 1.1664, 0.1936,
  0.7396, 1.1881, 0.4096,
  0.5929, 1.0404, 0.3481,
  0.6084, 1.0201, 0.3249,
  0.5184, 0.9409, 0.3136,
  1.3225, 0.7225, 0.2116,
  2.3409, 0.6889, 0.16,
  1.3225, 1.5129, 0.1936,
  _, 1.7424, _,
  _, 1.3689, _,
  _, _, 0.1444,
  _, _, 0.0961,
  _, _, _,
  _, _, _,
  _, _, _,
  1.9321, _, _,
  1.7689, _, _,
  _, 0.4761, 0.16,
  _, _, 0.0225,
  _, 0.6084, _,
  0.7569, 0.2809, 0.4356,
  0.2916, 0.1681, 0.5041,
  0.2209, 0.16, 0.4624,
  0.2916, 0.1764, 0.3364,
  0.2304, 0.1764, 0.2809,
  0.2809, 0.1936, 0.5329,
  0.2601, 0.3364, 0.1369,
  0.3721, 0.2809, 0.1521,
  0.3364, 0.3249, 0.3364,
  0.2304, 0.2704, 0.4225,
  0.64, 0.2209, 0.5041,
  0.25, 0.1849, 0.1225,
  0.2304, 0.1936, 0.2116,
  0.3025, 0.2704, 0.36,
  0.3481, 0.36, 0.3481,
  0.2704, 0.3364, 0.2809,
  0.2025, 0.6084, 0.4489,
  0.1764, 0.2601, 0.4225,
  0.1369, 0.1444, 0.3721,
  0.16, 0.1296, 0.2209,
  0.09, 0.1296, 0.1764,
  0.1369, 0.1369, 0.1936,
  0.16, 0.2601, 0.2025,
  0.2601, 0.3249, 0.36,
  0.1225, _, _,
  _, _, _,
  0.4761, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  12.5316, 2.1904, 0.8281,
  14.44, 5.1076, 0.4761,
  3.2041, 0.5041, 0.3481,
  0.9604, 1.5376, 0.3025,
  1.6129, 5.1984, 0.2601,
  1.2996, 3.9601, 0.2025,
  0.2601, 0.3969, 0.1444,
  0.4356, 0.2116, 0.16,
  0.81, 0.2304, 0.1444,
  0.3364, 0.1849, 0.1521,
  0.3481, 0.1764, 0.16,
  0.2401, 0.1936, 0.1849,
  0.1936, 0.1296, 0.1444,
  0.6561, 0.1521, 0.1369,
  0.2116, 0.1369, 0.1369,
  0.1444, 0.2025, 0.1521,
  0.1369, 0.2209, 0.1444,
  0.1296, 0.2116, 0.1296,
  0.1296, 0.1849, 0.1296,
  0.2025, 0.1849, 0.1156,
  0.1156, 0.2209, 0.1369,
  0.1156, 0.2304, 0.1444,
  0.1849, 0.4624, 0.1681,
  0.1936, 0.25, 0.1521,
  0.1444, 0.1225, 0.1369,
  0.1521, 0.1296, 0.1444,
  0.2209, 0.1444, 0.1849,
  0.2916, 0.1764, 0.2025,
  0.3481, 0.1849, 0.2704,
  0.2401, 0.1936, 0.2401,
  0.2916, 0.2704, 0.2116,
  0.25, 0.25, 0.2209,
  0.2116, 0.3136, 0.2704,
  0.2601, 0.2809, 0.2401,
  0.2401, 0.2304, 0.25,
  0.2916, 0.1849, 0.2209,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0.4761, 0.3481, 0.2209,
  0.4489, 0.3481, 0.2401,
  0.3844, 0.3721, 0.2601,
  0.49, 0.2916, 0.25,
  0.5625, 0.3136, 0.2704,
  0.6084, 0.3364, 0.2704,
  0.7744, 0.6889, 0.2916,
  1, 0.49, 0.3025,
  0.7225, 0.5041, 0.3481,
  0.81, 0.7921, 0.3249,
  1.1449, 1.44, 0.7056,
  1.4884, 1.6384, 1.1449,
  1.7161, 1.5376, 1.2769,
  2.3409, 1.3456, 1.2321,
  2.9584, 1.2544, 1.21,
  3.61, 1.1881, 1.1881,
  4, 1.2544, 0.9801,
  2.7889, 1.5129, 0.6889,
  1.0609, 1.3689, 0.4489,
  0.6889, 1.0609, 0.3844,
  1.1881, 1, 0.3364,
  1.1881, 1.1449, 0.3721,
  1.1881, 1.3924, 0.36,
  1.1664, 1.3456, 0.3136,
  0.9801, 1.1664, 0.3136,
  1.0201, 1.1664, 0.3844,
  0.9216, 1.1025, 0.3136,
  0.9604, 0.5625, 0.16,
  0.8836, 1.1025, 0.1764,
  0.36, 1.0816, 0.1369,
  0.7744, 1.0201, 0.16,
  2.7889, 1.3225, 0.1521,
  8.9401, 0.8281, 0.2916,
  1, 0.5329, 0.25,
  0.64, 0.5625, 0.3249,
  0.8836, 0.2704, 0.3481,
  0.6724, 0.3721, 0.25,
  0.5184, 0.4761, 0.3481,
  0.25, 0.2809, 0.4761,
  0.3844, 0.2401, 0.2116,
  0.2704, 0.3481, 0.1681,
  0.2704, 0.5329, 0.1764,
  0.3721, 0.9604, 0.1681,
  0.1369, 0.2809, 0.1156,
  0.1089, 0.1444, 0.1156,
  0.2025, 0.25, 0.1024,
  0.0841, 0.1444, 0.09,
  0.0961, 0.1444, 0.1024,
  0.25, 0.2704, 0.1681,
  0.3721, 0.2916, 0.1521,
  0.1764, 0.1681, 0.1369,
  0.2116, 0.2025, 0.1521,
  0.1521, 0.2209, 0.1764,
  0.1764, 0.2025, 0.1681,
  0.1521, 0.2401, 0.2025,
  0.2304, 0.2809, 0.1225,
  0.1444, 0.2809, 0.1681,
  0.1089, 0.2704, 0.1225,
  0.3136, 0.6241, 0.1444,
  0.1936, 0.2304, 0.1296,
  0.2209, 0.2025, 0.1521,
  0.16, 0.5476, 0.2116,
  0.2401, 0.2304, 0.1369,
  0.5625, 0.2304, 0.16,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0.7225, 0.6889, 0.1024,
  0.7056, 0.7225, 0.1089,
  1.6384, 0.5625, 0.1296,
  1.9321, 0.5625, 0.16,
  0.5041, 0.36, 0.1444,
  _, 0.4761, 0.1936,
  _, 0.8836, 0.2116,
  _, 0.3721, 0.0441,
  _, 0.4225, 0.1681,
  1.1881, 0.5625, 0.2601,
  0.5776, 0.6241, 0.2809,
  0.8281, 0.6561, 0.2601,
  0.6724, 0.49, 0.2025,
  0.6241, 0.64, 0.2304,
  0.8649, 0.64, 0.2401,
  0.6241, 0.4096, 0.2025,
  0.7225, 0.4096, 0.1849,
  1.0201, 0.8649, 0.1849,
  1.5625, 0.7569, 0.2209,
  0.9409, 0.5184, 0.1444,
  0.7744, 0.7225, 0.1225,
  0.64, 0.6561, 0.1444,
  0.4761, 1, 0.1369,
  0.5041, 0.8281, 0.2025,
  0.9409, 0.7921, 0.25,
  _, _, 0.16,
  0.4096, 0.6561, 0.1681,
  _, 0.7056, 0.2304,
  0.3844, 3.0976, 0.2401,
  0.2704, 1.1236, 0.2809,
  0.5625, 3.3856, 0.3136,
  1.2996, 6.8644, 1.96,
  2.2201, 3.0625, 1.7689,
  0.6084, 2.4649, 0.8649,
  0.4761, 1.2996, 0.7744,
  0.3481, 1.5129, 0.8464,
  0.4761, 1.5129, 0.7056,
  0.5329, 1.21, 0.5041,
  0.5041, 1.1664, 0.8464,
  0.5929, 1.0609, 0.9216,
  0.3136, 0.9409, 0.8464,
  0.3025, 1.4161, 0.2916,
  0.3721, 1.6641, 0.6889,
  0.3136, 0.8836, 1.1881,
  0.4225, 1.0404, 0.5329,
  0.16, 0.4761, 0.3721,
  0.1521, 0.2704, 0.25,
  0.1936, 0.4624, 0.36,
  0.2025, 0.1764, 0.4225,
  0.2401, 0.2704, 0.2025,
  0.25, 0.2704, 0.2916,
  0.3364, 0.4761, 0.25,
  0.3364, 0.2401, 0.2116,
  0.2704, 0.3025, 0.3969,
  0.2401, 0.25, 0.3025,
  0.3136, 0.2916, 0.2809,
  0.3481, 0.2601, 0.3721,
  0.4489, 0.3844, 0.3969,
  0.3721, 0.4489, 0.36,
  0.3025, 0.2704, 0.4489,
  0.2916, 0.3844, 0.2401,
  0.25, 0.2601, 0.2116,
  0.4489, 0.5476, 0.3721,
  0.2601, 0.1764, 0.3025,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0.4489, 0.5041, 0.2025,
  0.5184, 0.4489, 0.1936,
  0.5929, 0.6724, 0.2916,
  0.5776, 0.9216, 0.3136,
  0.7056, 0.8464, 0.4489,
  0.64, 0.64, 0.3721,
  0.8649, 0.5041, 0.3249,
  0.7056, 1.0404, 0.3249,
  1.21, 0.5476, 0.2809,
  _, _, _,
  0.3721, _, _,
  0.6889, 0.2601, _,
  1.0201, 0.8649, 0.2025,
  1.5376, 1.4884, 0.2916,
  1.4641, 1.7689, _,
  1.7956, 1.1881, 0.4761,
  1.1881, 0.8464, 0.3721,
  1.1664, 0.9025, 0.3025,
  1.21, 1.4161, 0.2704,
  1.0201, 0.81, 0.2809,
  1.1449, 0.5929, 0.2116,
  1.0404, 0.9216, 0.2304,
  0.5776, 0.5929, 0.1225,
  0.2704, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0.2704, 0.1681, 0.25,
  0.2401, 0.1681, 0.4096,
  0.2304, 0.2304, 0.09,
  0.3025, 0.1849, 0.1089,
  0.2809, 0.2704, 0.1369,
  0.2601, 0.3025, 0.1444,
  0.2809, 0.3136, 0.16,
  0.3136, 0.2304, 0.1444,
  0.36, 0.2304, 0.1444,
  0.7056, 0.3025, 0.2304,
  1.1881, 0.4761, 0.49,
  0.6889, 0.2601, 0.3249,
  0.4225, 0.2601, 0.3364,
  0.2916, 0.1764, 0.4761,
  0.2916, 0.0841, 0.16,
  0.1681, 0.0841, 0.1849,
  0.1849, 0.1089, 0.1369,
  0.25, 0.1089, 0.1444,
  0.2809, 0.1296, 0.1764,
  0.3844, 0.2809, 0.1225,
  0.2809, 0.09, 0.1225,
  0.16, 0.1521, 0.1156,
  0.1936, 0.2601, 0.1444,
  0.2025, 0.2025, 0.1764,
  0.1849, 0.1849, 0.16,
  0.2116, 0.1681, 0.1296,
  0.3364, 0.1521, 0.1156,
  0.2809, 0.2809, 0.2209,
  0.2116, 0.1521, 0.2304,
  0.1936, 0.1936, 0.2401,
  0.2401, 0.16, 0.2601,
  0.81, 0.4356, 0.2809,
  0.7056, 0.5625, 0.4096,
  0.8281, 0.6241, 0.36,
  0.7921, 0.64, 0.2601,
  0.7744, 0.5476, 0.25,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0.8281, 0.64, 0.2704,
  0.5184, 0.6561, 0.3364,
  0.6724, 0.49, 0.2304,
  0.81, 0.6561, 0.2601,
  0.7056, 0.7921, 0.2209,
  0.5041, 0.5184, 0.2304,
  0.3844, 0.3481, 0.2401,
  0.4225, 0.5329, 0.2916,
  0.5184, 0.5929, 0.2916,
  0.6241, 0.4624, 0.1296,
  0.7225, 0.7569, 0.1444,
  0.7225, 0.5041, 0.1681,
  0.6724, 0.5776, 0.2025,
  0.6561, 0.7396, 0.2304,
  0.7056, 0.7921, 0.2025,
  0.7569, 0.7744, 0.2116,
  1.0816, 1.0816, 0.2809,
  1.1025, 2.0449, 0.2916,
  0.8464, 2.1904, 0.3481,
  0.8649, 3.0625, 0.3481,
  0.9216, 3.61, 0.36,
  1.0816, 2.9929, 0.3025,
  0.9604, 1.5876, 0.2601,
  1.1025, 0.9409, 0.2116,
  1.1449, 1.1881, 0.3249,
  0.6889, 0.6561, 0.1936,
  0.6084, _, 0.1225,
  _, _, 0.0841,
  1.0816, 1.44, 0.8649,
  0.6561, 1.4884, 0.8281,
  1.0609, 0.4624, 0.5476,
  0.7569, 0.3364, 1.1236,
  0.3249, 0.2809, 0.2601,
  0.4225, 0.2601, 0.2601,
  0.2209, 0.3136, 0.2304,
  0.1444, 0.1764, 0.1521,
  0.1764, 0.3969, 0.1444,
  0.1225, 0.1521, 0.1225,
  0.1444, 0.1849, 0.1444,
  0.1764, 0.25, 0.1764,
  0.2025, 0.4761, 0.1369,
  0.1156, 0.2209, 0.1156,
  0.09, 0.1681, 0.1156,
  0.0961, 0.1849, 0.1225,
  0.1156, 0.1521, 0.1024,
  0.0841, 0.1681, 0.1024,
  0.1024, 0.1296, 0.1369,
  0.1225, 0.1521, 0.1369,
  0.1156, 0.1521, 0.1444,
  0.1764, 0.2304, 0.1681,
  0.1681, 0.2401, 0.2116,
  0.2116, 0.3481, 0.2304,
  0.2025, 0.4225, 0.4096,
  0.3025, 0.2916, 0.1849,
  0.2916, 0.6724, 0.2304,
  0.5476, 0.2916, 0.2601,
  0.7921, 0.9025, 0.1681,
  0.7056, 0.9216, 0.2025,
  0.5776, 0.6889, 0.2304,
  0.4225, 0.3721, 0.2704,
  0.1521, 0.1369, 0.2304,
  0.7056, 0.7569, 0.2401,
  0.36, 0.4624, 0.2025,
  0.2116, 0.3136, 0.1764,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0.2304, 0.3364, 0.1444,
  0.2601, 0.3364, 0.1296,
  0.2704, 0.64, 0.1296,
  0.3249, 0.2304, 0.1521,
  0.6724, 0.3025, 0.1764,
  0.5929, 0.64, 0.1444,
  0.6241, 0.6241, 0.1764,
  0.6084, 0.4761, 0.1936,
  0.3969, 0.3364, 0.1764,
  0.4489, 0.4624, 0.2025,
  0.3025, 0.4096, 0.3025,
  0.7225, 0.3969, 0.3481,
  0.49, 0.3136, 0.2809,
  0.4096, 0.64, 0.1225,
  0.7569, 0.4489, _,
  2.9241, 0.5184, 0.2809,
  2.4649, 0.6084, 0.2916,
  1.6641, 0.6724, 0.2704,
  1.9321, 0.5476, 0.2401,
  2.1904, 0.5929, 0.2809,
  2.2801, 0.7056, 0.2304,
  1.0201, 0.7396, 0.2304,
  0.7744, 0.81, 0.2401,
  0.6889, 0.6724, 0.1369,
  0.7225, 0.81, 0.1764,
  0.8464, _, 0.3249,
  0.5625, 0.6241, 0.2401,
  _, 0.5776, 0.1521,
  1.3924, 1.2996, 1.5625,
  1.21, 0.9801, 1.1449,
  0.7744, 0.5476, 1.9881,
  0.8464, 0.4624, 1.5376,
  0.81, 0.3136, 0.9801,
  0.7569, 0.2304, 0.6241,
  0.5625, 0.2116, 0.49,
  0.3249, 0.2601, 0.2209,
  0.25, 0.1764, 0.1764,
  0.3969, 0.2025, 0.2401,
  0.4761, 0.4489, 0.4356,
  0.5929, 0.2401, 0.2601,
  0.3136, 0.16, 0.6889,
  0.4761, 0.1089, 0.49,
  0.2601, 0.1089, 0.1849,
  0.2401, 0.2209, 0.7744,
  0.81, 0.3481, 0.8649,
  0.3364, 0.25, 0.7225,
  0.2601, 0.1936, 1.5129,
  0.1681, 0.1444, 0.6561,
  0.1369, 0.1296, 0.2304,
  0.1849, 0.1764, 0.2809,
  0.1296, 0.0961, 0.1369,
  0.1521, 0.0576, 0.1521,
  0.1849, 0.1936, 0.16,
  0.25, 0.1681, 0.1936,
  0.4356, 0.2704, 0.4096,
  0.5041, 0.3025, 0.64,
  0.3364, 0.25, 0.3721,
  0.2601, 0.2025, 0.2304,
  0.2304, 0.1681, 0.1764,
  0.2601, 0.1681, 0.2025,
  0.2704, 0.1681, 0.1849,
  0.2025, 0.1225, 0.2916,
  0.2304, 0.1521, 0.3721,
  0.25, 0.1764, 0.3136,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0.6889, 0.3136, 0.5329,
  0.7569, 0.3249, 0.5476,
  0.9409, 0.3364, 0.5929,
  1.0201, 0.3025, 0.5329,
  1.0816, 0.3721, 0.6241,
  1.1236, 0.3364, 0.7744,
  0.8649, 0.3721, 0.7569,
  1.0816, 0.3969, 0.6084,
  1.2996, 0.4489, 0.4624,
  1.2544, 0.49, _,
  _, 0.4489, 0.1089,
  _, 0.4624, _,
  1.21, 0.5625, _,
  1.6129, 1.5625, 0.1225,
  1.4641, 1.3225, 0.4761,
  1.5625, 2.0736, 0.4356,
  1.5376, 2.6896, 0.4096,
  1.5876, 3.3124, 0.3969,
  1.1881, 2.1609, 0.3969,
  1.1881, 0.9604, 0.49,
  1.1025, 1.3225, 0.5041,
  1.3924, 1.7689, _,
  1.5876, 0.9801, _,
  1.0816, 1.1881, 0.16,
  1.1025, 1.8225, 0.2116,
  1.1236, 1.69, 0.36,
  0.5625, 0.7569, _,
  _, 0.8649, _,
  0.2304, 0.6561, 0.1296,
  0.8649, 0.6561, 0.1444,
  0.4624, 0.7225, 0.1936,
  0.4761, 0.64, 0.1521,
  0.3249, 0.9409, 0.1369,
  0.3364, 1.5129, 0.1764,
  0.3721, 0.36, 0.1936,
  0.49, 0.36, 0.36,
  0.4096, 1.96, 0.3481,
  0.49, 0.4489, 0.4356,
  0.7569, 0.5184, 0.5041,
  0.5184, 0.64, 0.5041,
  0.49, 0.6561, 0.4761,
  0.5625, 0.5041, 0.5041,
  0.6084, 0.49, 0.5476,
  0.49, 0.3364, 0.4624,
  0.4624, 0.4356, 0.5776,
  0.6561, 0.3136, 0.5625,
  0.6889, 0.2304, 0.5329,
  0.8836, 0.7396, 0.64,
  0.6724, 0.5929, 0.6561,
  0.7056, 0.4489, 0.7921,
  0.64, 0.3364, 0.4761,
  0.5184, _, 0.5929,
  0.4225, _, 0.3481,
  0.4225, _, 0.5184,
  _, _, 0.4356,
  _, _, _,
  1.5376, 0.6889, 0.8836,
  1.5376, _, 0.7921,
  0.2704, 0.16, 0.1681,
  1.2996, _, 0.5184,
  0.0961, _, 0.36,
  1.0201, _, 0.5625,
  1.0201, 0.81, 0.6561,
  1.1025, 0.5476, 0.5625,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  1.2321, 0.7396, 0.7569,
  1.2321, 1.3689, 1,
  1.6384, 2.1025, 1.1236,
  2.1316, 2.4649, 1.1664,
  2.6244, 2.5921, 1.1881,
  2.7556, 2.6569, 1.1236,
  2.5281, 2.4964, 1.0404,
  2.1025, 2.4964, 0.9801,
  1.9321, 1.9044, 1,
  2.2201, 1.69, 0.8281,
  2.6569, 0.5776, 0.7225,
  2.8224, _, 0.4624,
  1.3689, _, 0.2601,
  1.7689, 0.3721, 0.4761,
  1.7956, 0.49, 0.4096,
  1.7424, 0.5929, 0.5929,
  1.2769, 1.5876, 0.5929,
  1.0201, 1.3924, 0.5776,
  0.9216, 1.0816, 0.5929,
  0.81, 0.81, 0.5929,
  6.0516, _, 0.6724,
  5.4756, 0.9025, 0.4489,
  4.4521, 1.44, 0.2809,
  4.2849, _, 0.2809,
  4.41, _, 0.2025,
  _, _, 0.1764,
  _, _, 0.1849,
  5.6169, 0.7056, 0.1681,
  0.64, 1.21, 0.49,
  0.8649, 3.8416, 0.7921,
  0.5625, 0.6241, 0.5184,
  1.3924, 0.7744, 0.3025,
  1.3456, 0.7569, 0.3364,
  1.6641, 2.7889, 0.2916,
  0.9025, 0.2916, 0.3844,
  0.7569, 1.3225, 0.4225,
  0.9025, 0.4761, 0.3136,
  0.5929, 0.5041, 0.2809,
  0.5625, 0.5329, 0.25,
  0.2209, 0.7921, 0.2025,
  0.3136, 0.4489, 0.1681,
  0.25, 0.3969, 0.1521,
  0.2304, 0.36, 0.1849,
  0.1764, 0.3481, 0.16,
  0.16, 0.2916, 0.1296,
  0.0961, 0.2704, 0.1089,
  0.1156, 0.2809, 0.1089,
  0.1764, 0.3136, 0.1024,
  0.1156, 0.3721, 0.1024,
  0.0784, 0.3481, 0.1089,
  0.1089, 0.3364, 0.1089,
  0.1225, 0.25, 0.1156,
  0.1089, 0.1764, 0.1296,
  0.1225, 0.1521, 0.1225,
  0.0961, 0.1444, 0.1156,
  0.1296, 0.2025, 0.1225,
  0.1444, 0.5476, 0.1764,
  0.2209, 0.16, 0.3025,
  0.1764, 0.2601, 0.1764,
  0.2025, 0.5041, 0.16,
  0.4489, 2.3409, 0.1681,
  0.1849, 0.2809, 0.1156,
  0.2304, 0.2209, 0.1936,
  0.2601, 0.2304, 0.1849,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0.36, 0.3721, 0.1764,
  0.3249, 0.3025, 0.1764,
  0.36, 0.3721, 0.1764,
  0.3969, 0.5625, 0.1681,
  0.4096, 0.4096, 0.1681,
  0.4356, 0.4624, 0.1681,
  0.4624, 0.7225, 0.1764,
  0.5929, 0.9604, 0.2116,
  1.2996, 0.9025, 0.1764,
  0.4761, 0.5041, 0.2401,
  0.9801, _, 0.3249,
  0.6889, 0.9604, 0.36,
  0.5476, 0.4356, 0.2401,
  0.7396, 0.5625, 0.4356,
  0.8281, 0.6241, 0.3136,
  0.9409, 0.9409, 0.3025,
  0.9409, 1.0816, 0.3136,
  0.6889, 1.1025, 0.3249,
  1.0201, 1.21, 0.2704,
  1.2544, 1.1664, 0.25,
  1.5876, 0.64, 0.2116,
  2.0164, 0.9216, 0.2025,
  1.8496, 1.0201, 0.2025,
  0.8464, 1.0816, 0.2209,
  0.9604, 1.4641, 0.2209,
  1.0816, 1.8225, 0.2025,
  0.7744, 2.3104, 0.25,
  0.8836, 1.3225, 0.3481,
  18.4041, 2.9241, 1.0404,
  1.8769, 15.6025, 0.2704,
  1.9321, 2.9584, 0.2304,
  2.7889, 3.24, 0.1444,
  3.3489, 1.5876, 0.16,
  1.5129, 3.6481, 0.4489,
  1.4884, 1.1881, 0.2916,
  1.1025, 0.6724, 0.4356,
  0.6724, 1.2996, 0.3844,
  0.5329, 0.7225, 0.1936,
  0.5625, 0.3481, 0.2209,
  0.3969, 0.4225, 0.2401,
  0.3481, 0.3844, 0.0961,
  0.3249, 0.2916, 0.1764,
  1.5376, 0.3136, 0.3136,
  1.4161, 0.3721, 0.5625,
  0.6889, 0.3721, 0.7396,
  0.4356, 0.2916, 0.8649,
  0.4761, 0.2704, 0.6241,
  0.5329, 0.2025, 0.25,
  0.3481, 0.1764, 0.1936,
  0.25, 0.2209, 0.2809,
  0.3364, 0.2601, 0.3721,
  0.36, 0.2704, 0.3364,
  0.49, 0.3249, 0.36,
  0.4624, 0.3025, 0.3136,
  0.5329, 0.3364, 0.3721,
  0.5329, 0.2916, 0.3249,
  0.3721, 0.3249, 0.2916,
  0.4096, 0.3721, 0.3481,
  0.64, 0.3721, 0.3969,
  0.49, 0.3136, 0.3249,
  0.3721, 0.3969, 0.4096,
  0.2809, 0.5041, 0.2025,
  1.9881, 0.8281, 0.49,
  1.9881, 0.7396, 0.4489,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  2.2201, 0.6724, 0.4489,
  1.2321, 0.6889, 0.4761,
  1.2321, 0.8281, 0.5476,
  1.5376, 1.3225, 0.6084,
  1.4641, 1.69, 0.6241,
  1.69, 1.4161, 0.6241,
  1.1664, 1.4641, 0.64,
  1.1236, 1.4884, 0.6241,
  1.21, 1.5876, 0.6084,
  1.2996, 1.2769, 0.5184,
  1.7424, _, 0.4624,
  1.1449, 4.3681, 0.3136,
  1.69, 4.3264, 0.5041,
  2.5281, 4, 0.5329,
  1.96, 3.8809, 0.5776,
  1.5625, 3.5344, 0.5625,
  1.2996, 3.7249, 0.5329,
  1.2769, 3.3124, 0.5041,
  1.5376, 2.7556, 0.5184,
  1.1664, 1.2321, 0.3721,
  1.3225, 1.1236, 0.1936,
  0.5776, 0.8649, 0.2304,
  1.1025, 0.9216, 0.3844,
  2.6244, 0.9801, 0.2304,
  1.4884, 1.1881, 0.2025,
  1.96, 2.56, 0.2601,
  1.8496, 3.6864, 0.3136,
  1.5876, 3.5721, 0.4096,
  0.4096, 0.3721, 0.2116,
  0.2601, 0.3844, 0.2401,
  0.3364, 0.7225, 0.2025,
  0.3249, 2.0736, 0.1024,
  0.3481, 2.1904, 0.0576,
  1.1881, 3.1329, 0.09,
  0.7056, 4.5796, 0.6889,
  0.6561, 4.3264, 0.5929,
  0.6084, 4.2436, 0.6724,
  0.6889, 4.9284, 0.5929,
  0.8836, 5.5696, 0.5476,
  0.8649, 5.9536, 0.4761,
  0.9604, 6.8644, 0.3364,
  0.7921, 0.7056, 0.2209,
  0.2601, 0.6084, 0.1089,
  0.1444, 0.5184, 0.0676,
  0.1764, 1.1664, 0.09,
  0.1369, 2.7556, 0.0961,
  0.1225, 2.25, 0.0961,
  0.1681, 0.7569, 0.1225,
  0.3481, 0.49, 0.2916,
  0.3721, _, 0.1089,
  0.1089, 0.3136, 0.0961,
  0.1521, 0.2209, 0.1024,
  0.2025, 0.2916, 0.1156,
  0.2209, 0.2809, 0.1764,
  0.2025, 0.4096, 0.1089,
  0.1936, 0.2025, 0.1225,
  0.1521, 0.2209, 0.1156,
  0.0729, 0.2209, 0.1369,
  0.1764, 0.2116, 0.1521,
  0.3481, 0.5625, 0.16,
  0.3721, 0.8649, 0.2304,
  0.3481, 0.5929, 0.1681,
  0.3481, 0.5776, 0.1681,
  0.3364, 0.6084, 0.1521,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0.3721, 0.64, 0.1369,
  0.5041, 0.6889, 0.2025,
  0.6084, 0.6561, 0.25,
  0.8281, 0.0841, 0.1764,
  0.8281, 0.1936, 0.25,
  0.81, 0.36, 0.3364,
  0.4489, 0.3364, 0.2304,
  0.8281, 0.3364, 0.2304,
  1.2996, 0.3969, 0.2401,
  1.5876, 0.1764, _,
  0.7225, 0.3844, _,
  _, 0.36, _,
  1.5376, 0.3025, 0.1936,
  _, 0.6084, 0.16,
  _, 0.4489, 0.1296,
  _, 0.64, 0.1681,
  0.6084, 0.6241, _,
  0.4624, 0.4096, 0.1369,
  _, 0.4225, 0.2209,
  _, 0.3481, 0.1849,
  0.4356, 0.3844, 0.1089,
  0.49, 0.3844, 0.1024,
  0.5041, 0.4489, 0.1521,
  0.8464, 0.3364, 0.1369,
  0.9409, 0.1849, 0.1369,
  1.8496, _, 0.1024,
  0.8281, 0.3844, 0.1156,
  1.9044, _, 0.0841,
  5.4756, 1.8769, 0.5329,
  5.29, 1.69, 2.4649,
  2.2801, 0.8649, 1.4161,
  2.4336, 2.9241, 1.0609,
  1.9321, 2.0736, 0.9025,
  2.6569, 0.9801, 1.0404,
  2.7556, 0.4225, 0.7056,
  2.6244, 0.5184, 1.0816,
  1.5876, 0.6561, 1.3225,
  1.5129, 0.7569, 2.0164,
  1.9321, 1.5376, 2.3104,
  2.3716, 1.1881, 2.0736,
  2.5921, 1.2321, 2.2201,
  1.6129, 1.1449, 3.2761,
  1.8769, 1.0816, 1.4641,
  0.9604, 0.4225, 0.64,
  0.3721, 0.3721, 0.3025,
  0.3249, 0.3721, 0.36,
  0.4225, 1.3225, 0.36,
  0.4761, 0.49, 0.4624,
  0.5625, 0.6561, 0.2809,
  _, 0.3969, 0.2116,
  _, 0.36, _,
  _, _, _,
  0.5041, _, _,
  0.1089, _, _,
  _, 0.1296, _,
  _, _, _,
  1.0609, 0.4624, 0.2209,
  0.9409, 0.5041, 0.1089,
  0.7056, 0.6724, 0.25,
  0.64, 0.7569, _,
  0.5776, 0.8281, 0.1024,
  0.3721, 0.7569, _,
  0.3249, 0.9025, _,
  0.9025, 1.0201, 0.49,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  1.0816, 1.21, 0.5041,
  1.1025, 1.2996, 0.3844,
  1, 1.1236, 0.2401,
  0.8649, 1.0609, 0.2401,
  0.3969, 0.9409, 0.1521,
  _, 0.6889, _,
  0.2809, 0.7744, _,
  0.4624, 1.5625, 0.3025,
  1.1025, 1.1025, 0.5184,
  0.5776, 1.2544, _,
  _, 0.7921, _,
  _, 0.9409, _,
  _, 1, _,
  _, 1.9321, _,
  0.7056, 2.4336, 0.2601,
  1.3225, 2.1904, 0.6724,
  1.1236, 2.2801, 0.5776,
  0.8464, 2.1904, 0.5929,
  1.0816, 1.0404, 0.7396,
  0.5625, 0.7569, _,
  0.5329, 0.5625, _,
  0.3969, 0.7056, _,
  0.5625, 0.5776, 0.1156,
  0.5476, 0.7056, _,
  _, 0.4624, _,
  _, _, _,
  0.4761, 0.7921, _,
  _, 0.9025, _,
  1.0609, 1.9321, 1.1881,
  0.7569, 0.9409, 0.6561,
  1.0816, 1.0404, 0.7225,
  0.9801, 0.8836, 0.7569,
  1.3689, 0.6561, 1.0816,
  0.7744, 0.8281, 1.3924,
  1.1449, 0.9801, 1.0816,
  0.6724, 1.8225, 0.6889,
  0.3844, 0.4761, 0.8464,
  0.2704, 0.4225, 0.6084,
  0.49, 0.4761, 0.2025,
  0.1156, 0.2916, 0.1849,
  0.1369, 0.2304, 0.2209,
  0.7569, 0.5184, 0.3364,
  0.7569, 2.1316, 0.3844,
  0.5329, 0.49, 0.3969,
  0.2809, 0.2601, 0.4356,
  0.2916, 0.3136, 0.6889,
  0.1849, 0.2025, 0.2916,
  0.2116, 0.2116, 0.4624,
  0.2116, 0.2116, 0.2209,
  0.1296, 0.2116, 0.2304,
  0.1296, _, 0.1156,
  0.1936, 0.2304, 0.16,
  0.1764, 0.2304, 0.2025,
  0.3136, 0.2704, 0.1936,
  0.2025, _, 0.1936,
  _, _, _,
  0.1764, 0.2601, 0.1225,
  0.1681, 0.2809, 0.1089,
  0.5776, 0.8464, 0.1849,
  0.3969, 0.1296, 0.2401,
  1.1025, 1.0816, 0.1369,
  0.9409, 1.0404, 0.2601,
  1.1664, 1.44, 0.1521,
  0.9025, 0.4761, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, 0.9216, 0.1156,
  _, _, _,
  _, 0.3969, _,
  _, 0.5776, _,
  0.3844, 0.6561, 0.1156,
  0.5041, 0.7744, 0.1681,
  0.5041, 0.49, 0.1681,
  0.4356, 0.4356, 0.2601,
  _, _, 0.2401,
  _, _, _,
  _, _, _,
  0.2116, _, _,
  0.4761, _, _,
  0.4761, 0.64, _,
  0.7921, 0.7569, 0.3136,
  1.0816, 1.2544, _,
  _, 1.0609, 0.1764,
  _, 1, _,
  _, 0.6724, 0.2401,
  _, 0.7569, 0.1296,
  0.4096, 0.9409, 0.1444,
  _, _, 0.2209,
  _, 1.5129, _,
  _, _, _,
  0.3721, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  1.7956, 1.9044, 30.9136,
  0.8281, 0.7744, 0.6561,
  0.64, 0.5776, 0.3844,
  0.5929, 0.5041, 0.3249,
  1.0201, 0.4761, 0.3364,
  0.8649, 0.3364, 0.25,
  0.6724, 0.3025, 0.2209,
  0.7225, 0.5041, 0.2209,
  0.3721, 0.1681, 0.2025,
  0.3364, 0.16, 0.4096,
  0.3136, 0.1521, 0.2601,
  0.2209, 0.1936, 0.2209,
  0.2704, 0.1764, 0.3136,
  0.3025, 0.2401, 0.64,
  0.1764, 0.2209, 0.1936,
  0.1369, 0.1156, 0.16,
  0.1156, 0.1024, 0.16,
  0.1521, 0.0961, 0.1681,
  0.3364, 0.1024, 0.1521,
  0.3721, 0.0961, 0.1369,
  0.3136, 0.1089, 0.1156,
  0.3025, 0.1156, 0.1444,
  0.2116, 0.1296, 0.1369,
  0.1764, 0.1369, 0.1225,
  0.16, 0.1225, 0.1296,
  0.1681, 0.1296, 0.1369,
  0.2025, 0.1521, 0.1521,
  0.2025, 0.1521, 0.1764,
  0.2209, 0.1764, 0.2209,
  0.2304, 0.2116, 0.16,
  0.2304, 0.2401, 0.1764,
  0.25, 0.2601, 0.2025,
  0.1849, 0.2116, 0.2025,
  0.3481, 0.1936, 0.2209,
  0.2809, 0.2401, 0.2704,
  0.25, 0.2704, 0.2401,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0.4489, 0.3364, 0.2116,
  0.4489, 0.36, 0.2401,
  0.7569, 0.3025, 0.25,
  0.8464, 0.2916, 0.2209,
  0.8281, 0.3481, 0.2209,
  0.64, 0.49, 0.2601,
  0.6241, 0.9216, 0.3969,
  0.6724, 1.1236, 0.3364,
  0.7056, 1.3225, 0.3481,
  0.9025, 1.2996, 0.3844,
  0.7225, 1.2996, 0.2704,
  0.9409, 1.3225, 0.3844,
  1.1025, 0.9216, 0.4356,
  1.1449, 0.8281, 0.4624,
  1.3456, 1.5129, 0.5776,
  1.0609, 4.6656, 0.3969,
  0.6724, 3.3489, 0.3969,
  0.6561, 2.0164, 0.3364,
  0.7225, 1.5876, 0.3364,
  0.5625, 0.9216, 0.2209,
  0.81, 0.6561, 0.1849,
  0.7921, 1.4161, 0.2116,
  0.8649, 1.4641, 0.1681,
  0.5929, 1.9321, 0.25,
  0.6241, 1.9044, 0.2116,
  0.5625, 1.8496, 0.2304,
  0.6561, 1.5876, 0.1225,
  0.7225, 1.8496, 0.1024,
  2.4336, 2.6244, 0.2916,
  1.5876, 2.2801, 0.8836,
  0.5476, 2.5921, 0.3844,
  1.2544, 1.7424, 0.1521,
  1, 1, 0.2916,
  0.9216, 0.8464, 0.3136,
  0.6889, 0.8649, 0.2304,
  0.3481, 0.3481, 0.16,
  0.3364, 0.3249, 0.1369,
  0.3249, 0.2704, 0.1369,
  0.2916, 0.25, 0.1296,
  0.2916, 0.1936, 0.1156,
  0.2916, 0.1849, 0.1089,
  0.3025, 0.2401, 0.1024,
  0.36, 0.2401, 0.1024,
  0.2025, 0.25, 0.1089,
  0.5329, 0.5476, 0.2916,
  0.6724, 0.7225, 0.4356,
  0.6724, 0.5929, 0.4624,
  0.4761, 0.3481, 0.36,
  0.2809, 0.2601, 0.2401,
  0.2809, 0.2601, 0.2025,
  0.3025, 0.2601, 0.2025,
  0.3025, 0.2601, 0.1849,
  0.5184, 0.3364, 0.2401,
  0.5625, 0.5625, 0.2916,
  0.6561, 0.4225, 0.3025,
  _, _, _,
  3.2761, 0.5476, 0.3249,
  2.3104, 0.6084, 0.3364,
  0.49, 0.5476, 0.3025,
  0.5776, 0.49, 0.4356,
  0.4356, 0.4096, 0.4624,
  0.4225, 0.2809, 0.5184,
  0.5476, 0.3364, 0.3844,
  0.7569, 0.3364, 0.4096,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0.7396, 0.7569, 0.5184,
  1.0609, 0.64, 0.6241,
  1.3456, 0.6241, 0.5929,
  1.4884, 0.8836, 0.6241,
  1.4641, 0.5625, 0.7056,
  1.5376, 0.8464, 0.5476,
  1.3456, 0.8649, 0.4225,
  1.44, 0.6561, 0.2601,
  1.5376, 0.3481, _,
  0.9801, 0.5329, 0.2601,
  1.4161, 0.2916, 0.3364,
  1.7689, _, 0.3481,
  1.7161, _, 0.3969,
  1.2996, _, 0.4624,
  1.3924, 0.8649, 0.5776,
  1.3456, 1.4161, 0.6241,
  1.4641, 2.4964, 0.6724,
  1.2544, 2.5921, 0.5625,
  1.2769, 2.3409, 0.5476,
  1.1025, 3.3489, 0.5184,
  1.6384, 1.7689, 0.4225,
  1.2544, 1.21, 0.5041,
  1.1881, 0.3969, _,
  1.4641, _, _,
  1.8496, _, 0.3721,
  1.5129, 0.2601, 0.3721,
  1.6384, 1.1664, 0.2116,
  1.3225, 1.2321, 0.1849,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  13.1769, _, 0.0324,
  5.1076, 69.5556, 0.2304,
  3.3489, 9, 1,
  8.6436, 14.2884, 0.5041,
  9.3025, _, 3.3489,
  1.8225, 1.1236, 0.6724,
  3.4596, 3.0625, 0.5184,
  3.2761, 2.7225, 0.9216,
  1.96, 1.0404, 0.8649,
  2.0164, 0.7569, 0.8464,
  1.1236, 1.0404, 0.6241,
  1.1025, 1.0404, 0.6724,
  2.1904, 1.0404, 0.4624,
  1.6384, 0.9801, 0.49,
  0.9801, 1.44, 0.5329,
  1.6641, 1.6129, 0.7056,
  1.3456, 2.2201, 0.5184,
  1.4641, 2.6896, 1.1664,
  1.7956, 2.89, 1.2996,
  2.6896, 2.9929, 1.0201,
  3.4596, 2.8561, 1.1664,
  3.3489, 2.8561, 1.5129,
  2.7225, 2.6569, 1.21,
  3.2761, 2.3409, 1.4161,
  1.2544, 3.7249, 2.7556,
  1.3456, 3.5344, 2.7556,
  1.5876, 1.7689, 4.3264,
  1.21, 2.56, 0.7225,
  1.0609, 2.6896, 0.64,
  0.7396, 0.4356, 0.8649,
  0.4624, 0.5329, 0.5329,
  22.7529, 9.8596, 3.4596,
  12.6736, 6.0516, 2.9929,
  0.64, 1.8496, 0.4096,
  15.5236, 7.8961, 3.9601,
  29.9209, 1.44, 0.9801,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  29.0521, 1.21, 2.4964,
  21.9024, 10.24, 2.4964,
  16.9744, 12.6736, 1.2321,
  12.6025, 3.2761, 0.7921,
  11.6964, 6.1009, 0.6561,
  13.2496, 8.5264, 0.7056,
  1.0816, 7.5076, 0.7569,
  1, 6.6564, 0.7921,
  1.2544, _, 0.7225,
  1.2769, _, 0.5776,
  2.0736, 17.5561, 0.64,
  2.56, 3.5344, 0.7056,
  2.3409, 4.7961, 0.7744,
  2.0736, 4, 0.7396,
  1.96, 4.41, 0.7056,
  1.7424, 5.29, 0.6889,
  1.69, 10.4329, 0.6241,
  1.4884, 8.0656, 0.5329,
  1.6641, 4.7961, 0.4624,
  1.3225, 1.2321, 0.2704,
  1.4641, 1.2769, 0.3481,
  1.5376, 1.21, 0.25,
  1.1881, 1.2996, 0.2601,
  1.0201, 1.1881, 0.25,
  0.9216, 1.0816, 0.25,
  _, 0.8649, 0.1764,
  1.7424, _, 0.2209,
  0.7225, _, _,
  0.2601, 0.4761, 0.1849,
  0.1764, 0.5041, 0.2116,
  0.2401, 0.6561, 0.2025,
  0.4489, 0.7056, 0.5041,
  1.3225, 1.1881, 0.25,
  0.9409, 1.6641, 0.0961,
  1.6641, 0.4225, 1,
  1.2544, 0.4489, 0.3481,
  0.9409, 0.4624, 0.5041,
  0.64, 0.5041, 0.9409,
  1.9044, 1.1881, 3.7249,
  0.1296, 1.6384, 0.0961,
  0.1521, 1.8225, 0.09,
  2.4649, 1.3689, 1.9321,
  1.0404, 0.6561, 1.5129,
  0.4096, 0.7921, 0.6241,
  0.4489, 0.8649, 0.7744,
  0.8464, 0.6889, 0.5929,
  0.4761, 0.3721, 0.4225,
  0.3969, 0.3481, 0.2601,
  0.5329, 0.3844, 0.3481,
  0.7396, 0.49, 0.5184,
  1.2769, 0.7396, 0.4761,
  0.7921, 0.64, 0.5929,
  0.5041, 0.4761, 0.4489,
  0.36, 0.64, 0.3844,
  0.3025, 0.2304, 0.2304,
  0.2209, 0.25, 0.1849,
  0.6889, 1.0816, 0.4356,
  0.1849, 0.36, 0.3025,
  0.2916, 0.25, 0.1764,
  0.7921, 1.3225, 0.3249,
  0.4489, 1.0201, 0.3481,
  0.2916, 0.7396, 0.3136,
  0.3721, 0.5184, 0.2916,
  0.3364, 1.2544, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, 0.3481,
  _, 0.8836, 0.5184,
  _, _, 0.2601,
  _, 0.4761, 0.2916,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, 0.1521, _,
  _, _, _,
  _, _, _,
  _, _, 0.16,
  _, _, _,
  _, _, _,
  _, 0.7056, _,
  _, 0.8836, _,
  0.5476, 1.1881, _,
  0.6724, _, _,
  0.3136, _, _,
  0.81, _, _,
  _, _, _,
  _, _, _,
  0.3969, _, _,
  0.9025, _, _,
  1.4161, _, _,
  1.8496, 0.25, _,
  8.1225, 1.1025, 0.16,
  8.1796, 0.8464, 1.3456,
  5.29, 0.81, 1.0201,
  2.25, 0.7396, 0.8464,
  2.1609, 0.9025, 0.9604,
  1.8496, 0.8464, 0.7744,
  2.7225, 1.0816, 0.9216,
  4.6225, 3.2041, 2.4025,
  2.9241, 5.0176, 1.7424,
  1.0201, 0.6241, 0.1764,
  0.3025, 4.7089, 0.1764,
  0.1681, 2.8224, 0.1089,
  1.2321, 1.0404, 0.1681,
  0.9409, 0.5776, 0.1369,
  0.5184, 0.5041, 0.3136,
  0.2401, 0.5184, 0.1936,
  0.2304, 0.1681, 0.0676,
  0.1849, 0.1681, 0.1156,
  0.2209, 0.4761, 0.0784,
  0.49, 0.1681, 0.1089,
  0.1849, _, 0.1024,
  _, _, 0.0841,
  _, _, 0.1024,
  _, 0.1849, 0.0784,
  _, _, 0.0784,
  _, _, 0.0324,
  _, _, 0.0841,
  _, _, 0.0361,
  _, _, 0.0576,
  _, _, 0.0784,
  0.2916, 0.64, 0.1225,
  0.4096, 0.3721, 0.0289,
  0.49, 1.1449, 0.1936,
  1.1025, 0.8464, 0.1521,
  1.2321, 0.5184, 0.16,
  3.7249, 0.36, 0.2304,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  3.7249, 0.9604, 0.1764,
  3.5721, 1.4641, 0.2401,
  0.8281, 0.3249, 0.2025,
  _, _, 0.3025,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, 0.2809,
  _, _, _,
  _, _, 0.1156,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0.3481, 0.9025, 0.2601,
  0.5041, 0.3136, 0.2704,
  0.6084, 0.5625, 0.49,
  0.7396, 0.6889, 1.0609,
  0.6084, 0.6724, 0.9604,
  0.5184, 0.3721, 0.8649,
  0.2601, 0.2601, 0.4225,
  0.4096, 0.3364, 0.8281,
  0.3721, 0.3025, 0.64,
  0.4624, 0.2809, 0.6561,
  0.81, 0.4225, 0.5476,
  0.5041, 0.5625, 0.7744,
  0.2304, 0.2401, 0.2401,
  0.1936, 0.1444, 0.2025,
  0.1849, 0.1521, 0.2916,
  0.2209, 0.1764, 0.3481,
  0.36, 0.1521, 0.2304,
  0.3844, 0.2116, 0.3249,
  0.2704, 0.25, 0.2401,
  0.2401, 0.25, 0.2025,
  0.2209, 0.2601, 0.1936,
  0.3136, 0.25, 0.2025,
  0.2601, 0.2601, 0.2401,
  0.2916, 0.3969, 0.2601,
  0.3844, 0.25, 0.2704,
  0.36, 0.2304, 0.2601,
  0.3364, 0.2809, 0.1296,
  0.2304, _, _,
  1.69, 1.0201, 0.3721,
  2.1025, 0.8836, 0.5041,
  1.4161, 0.8281, 0.3721,
  1.3225, 0.81, 0.3969,
  1.6129, 0.7056, 0.4356,
  0.9409, 0.6241, 0.5329,
  0.7225, 0.3721, 0.4761,
  0.5476, 0.3364, 0.1521,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  0.9409, 0.7744, 0.5776,
  1.0404, 0.9216, 0.5476,
  0.7225, 1.3225, 0.6084,
  1.1664, 0.64, 0.2809,
  0.7921, 0.5476, 0.2209,
  0.9409, _, _,
  1.0404, _, 0.3364,
  _, 0.8836, 0.3721,
  _, 0.5329, 0.3136,
  _, _, 0.49,
  _, _, _,
  _, _, 0.4624,
  _, _, _,
  _, _, _,
  _, _, _,
  _, _, _,
  3.1329, 1.9321, _,
  1.4641, 1.6129, 0.6724,
  1.5376, 2.0736, 0.7569,
  1.8496, 2.7225, 0.7396,
  2.0449, 2.9929, 0.5625,
  2.7225, 2.3104, 0.6241,
  1.96, _, 0.5329,
  _, _, 0.3025,
  _, _, 0.2304,
  1.2321, _, 0.3025,
  1.44, 1.1449, 0.4225,
  0.5776, 0.1849, 0.3844 ;
}
