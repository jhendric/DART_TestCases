netcdf wc13_grd {
dimensions:
	xi_u = 55 ;
	eta_u = 55 ;
	xi_v = 56 ;
	eta_v = 54 ;
	xi_rho = 56 ;
	eta_rho = 55 ;
	xi_psi = 55 ;
	eta_psi = 54 ;
	bath = UNLIMITED ; // (1 currently)
	coast = 12779 ;
variables:
	int spherical ;
		spherical:long_name = "grid type logical switch" ;
		spherical:flag_values = "0, 1" ;
		spherical:flag_meanings = "Cartesian spherical" ;
	double xl ;
		xl:long_name = "domain length in the XI-direction" ;
		xl:units = "meter" ;
	double el ;
		el:long_name = "domain length in the ETA-direction" ;
		el:units = "meter" ;
	double angle(eta_rho, xi_rho) ;
		angle:long_name = "angle between xi axis and east" ;
		angle:units = "radians" ;
		angle:coordinates = "lon_rho lat_rho" ;
	double h(eta_rho, xi_rho) ;
		h:long_name = "Final bathymetry at RHO-points" ;
		h:units = "meter" ;
		h:coordinates = "lon_rho lat_rho" ;
	double hraw(bath, eta_rho, xi_rho) ;
		hraw:long_name = "Working bathymetry at RHO-points" ;
		hraw:units = "meter" ;
		hraw:coordinates = "lon_rho lat_rho bath" ;
	double alpha(eta_rho, xi_rho) ;
		alpha:long_name = "Weights between coarse and fine grids at RHO-points" ;
		alpha:coordinates = "lon_rho lat_rho" ;
	double f(eta_rho, xi_rho) ;
		f:long_name = "Coriolis parameter at RHO-points" ;
		f:units = "second-1" ;
		f:coordinates = "lon_rho lat_rho" ;
	double pm(eta_rho, xi_rho) ;
		pm:long_name = "curvilinear coordinate metric in XI" ;
		pm:units = "meter-1" ;
		pm:coordinates = "lon_rho lat_rho" ;
	double pn(eta_rho, xi_rho) ;
		pn:long_name = "curvilinear coordinate metric in ETA" ;
		pn:units = "meter-1" ;
		pn:coordinates = "lon_rho lat_rho" ;
	double dndx(eta_rho, xi_rho) ;
		dndx:long_name = "xi derivative of inverse metric factor pn" ;
		dndx:units = "meter" ;
		dndx:coordinates = "lon_rho lat_rho" ;
	double dmde(eta_rho, xi_rho) ;
		dmde:long_name = "eta derivative of inverse metric factor pm" ;
		dmde:units = "meter" ;
		dmde:coordinates = "lon_rho lat_rho" ;
	double x_rho(eta_rho, xi_rho) ;
		x_rho:long_name = "x location of RHO-points" ;
		x_rho:units = "meter" ;
	double x_u(eta_u, xi_u) ;
		x_u:long_name = "x location of U-points" ;
		x_u:units = "meter" ;
	double x_v(eta_v, xi_v) ;
		x_v:long_name = "x location of V-points" ;
		x_v:units = "meter" ;
	double x_psi(eta_psi, xi_psi) ;
		x_psi:long_name = "x location of PSI-points" ;
		x_psi:units = "meter" ;
	double y_rho(eta_rho, xi_rho) ;
		y_rho:long_name = "y location of RHO-points" ;
		y_rho:units = "meter" ;
	double y_u(eta_u, xi_u) ;
		y_u:long_name = "y location of U-points" ;
		y_u:units = "meter" ;
	double y_v(eta_v, xi_v) ;
		y_v:long_name = "y location of V-points" ;
		y_v:units = "meter" ;
	double y_psi(eta_psi, xi_psi) ;
		y_psi:long_name = "y location of PSI-points" ;
		y_psi:units = "meter" ;
	double lon_rho(eta_rho, xi_rho) ;
		lon_rho:long_name = "longitude of RHO-points" ;
		lon_rho:units = "degree_east" ;
		lon_rho:standard_name = "longitude" ;
	double lon_u(eta_u, xi_u) ;
		lon_u:long_name = "longitude of U-points" ;
		lon_u:units = "degree_east" ;
		lon_u:standard_name = "longitude" ;
	double lon_v(eta_v, xi_v) ;
		lon_v:long_name = "longitude of V-points" ;
		lon_v:units = "degree_east" ;
		lon_v:standard_name = "longitude" ;
	double lon_psi(eta_psi, xi_psi) ;
		lon_psi:long_name = "longitude of PSI-points" ;
		lon_psi:units = "degree_east" ;
		lon_psi:standard_name = "longitude" ;
	double lat_rho(eta_rho, xi_rho) ;
		lat_rho:long_name = "latitude of RHO-points" ;
		lat_rho:units = "degree_north" ;
		lat_rho:standard_name = "latitude" ;
	double lat_u(eta_u, xi_u) ;
		lat_u:long_name = "latitude of U-points" ;
		lat_u:units = "degree_north" ;
		lat_u:standard_name = "latitude" ;
	double lat_v(eta_v, xi_v) ;
		lat_v:long_name = "latitude of V-points" ;
		lat_v:units = "degree_north" ;
		lat_v:standard_name = "latitude" ;
	double lat_psi(eta_psi, xi_psi) ;
		lat_psi:long_name = "latitude of PSI-points" ;
		lat_psi:units = "degree_north" ;
		lat_psi:standard_name = "latitude" ;
	double mask_rho(eta_rho, xi_rho) ;
		mask_rho:long_name = "mask on RHO-points" ;
		mask_rho:flag_values = 0., 1. ;
		mask_rho:flag_meanings = "land water" ;
		mask_rho:coordinates = "lon_rho lat_rho" ;
	double mask_u(eta_u, xi_u) ;
		mask_u:long_name = "mask on U-points" ;
		mask_u:flag_values = 0., 1. ;
		mask_u:flag_meanings = "land water" ;
		mask_u:coordinates = "lon_u lat_u" ;
	double mask_v(eta_v, xi_v) ;
		mask_v:long_name = "mask on V-points" ;
		mask_v:flag_values = 0., 1. ;
		mask_v:flag_meanings = "land water" ;
		mask_v:coordinates = "lon_rho lat_rho" ;
	double mask_psi(eta_psi, xi_psi) ;
		mask_psi:long_name = "mask on PSI-points" ;
		mask_psi:flag_values = 0., 1. ;
		mask_psi:flag_meanings = "land water" ;
		mask_psi:coordinates = "lon_psi lat_psi" ;
	double lon_coast(coast) ;
		lon_coast:long_name = "Coastline longitude" ;
		lon_coast:units = "degree_east" ;
	double lat_coast(coast) ;
		lat_coast:long_name = "Coastline latitude" ;
		lat_coast:units = "degree_north" ;

// global attributes:
		:type = "ROMS grid file" ;
		:title = "California Current System, 1/3 degree resolution (WC13)" ;
		:history = "Monday - December 11, 2006 - 11:00:00 AM" ;
data:

 spherical = 1 ;

 xl = 1764470.21024891 ;

 el = 2000391.13969695 ;

 angle =
  0.001454444122029, 0.001454444122029, 0.001454444122029, 
    0.00145444412202878, 0.001454444122029, 0.001454444122029, 
    0.00145444412202878, 0.001454444122029, 0.001454444122029, 
    0.00145444412202878, 0.001454444122029, 0.001454444122029, 
    0.00145444412202878, 0.001454444122029, 0.001454444122029, 
    0.00145444412202878, 0.001454444122029, 0.001454444122029, 
    0.00145444412202878, 0.001454444122029, 0.00145444412202878, 
    0.001454444122029, 0.00145444412202878, 0.001454444122029, 
    0.001454444122029, 0.001454444122029, 0.001454444122029, 
    0.001454444122029, 0.00145444412202878, 0.001454444122029, 
    0.001454444122029, 0.001454444122029, 0.00145444412202878, 
    0.001454444122029, 0.00145444412202878, 0.001454444122029, 
    0.001454444122029, 0.00145444412202878, 0.001454444122029, 
    0.001454444122029, 0.001454444122029, 0.00145444412202878, 
    0.001454444122029, 0.001454444122029, 0.00145444412202878, 
    0.001454444122029, 0.001454444122029, 0.00145444412202878, 
    0.001454444122029, 0.00145444412202878, 0.001454444122029, 
    0.001454444122029, 0.001454444122029, 0.001454444122029, 
    0.001454444122029, 0.001454444122029,
  0.00146907534809437, 0.00146907534809437, 0.00146907534809437, 
    0.00146907534809415, 0.00146907534809437, 0.00146907534809437, 
    0.00146907534809415, 0.00146907534809437, 0.00146907534809437, 
    0.00146907534809415, 0.00146907534809437, 0.00146907534809437, 
    0.00146907534809415, 0.00146907534809437, 0.00146907534809437, 
    0.00146907534809415, 0.00146907534809437, 0.00146907534809437, 
    0.00146907534809415, 0.00146907534809437, 0.00146907534809415, 
    0.00146907534809437, 0.00146907534809415, 0.00146907534809437, 
    0.00146907534809437, 0.00146907534809437, 0.00146907534809437, 
    0.00146907534809437, 0.00146907534809415, 0.00146907534809437, 
    0.00146907534809437, 0.00146907534809437, 0.00146907534809415, 
    0.00146907534809437, 0.00146907534809415, 0.00146907534809437, 
    0.00146907534809437, 0.00146907534809415, 0.00146907534809437, 
    0.00146907534809437, 0.00146907534809437, 0.00146907534809415, 
    0.00146907534809437, 0.00146907534809437, 0.00146907534809415, 
    0.00146907534809437, 0.00146907534809437, 0.00146907534809415, 
    0.00146907534809437, 0.00146907534809415, 0.00146907534809437, 
    0.00146907534809437, 0.00146907534809437, 0.00146907534809437, 
    0.00146907534809437, 0.00146907534809437,
  0.00148365685086094, 0.00148365685086094, 0.00148365685086094, 
    0.00148365685086072, 0.00148365685086094, 0.00148365685086094, 
    0.00148365685086072, 0.00148365685086094, 0.00148365685086094, 
    0.00148365685086072, 0.00148365685086094, 0.00148365685086094, 
    0.00148365685086072, 0.00148365685086094, 0.00148365685086094, 
    0.00148365685086072, 0.00148365685086094, 0.00148365685086094, 
    0.00148365685086072, 0.00148365685086094, 0.00148365685086072, 
    0.00148365685086094, 0.00148365685086072, 0.00148365685086094, 
    0.00148365685086094, 0.00148365685086094, 0.00148365685086094, 
    0.00148365685086094, 0.00148365685086072, 0.00148365685086094, 
    0.00148365685086094, 0.00148365685086094, 0.00148365685086072, 
    0.00148365685086094, 0.00148365685086072, 0.00148365685086094, 
    0.00148365685086094, 0.00148365685086072, 0.00148365685086094, 
    0.00148365685086094, 0.00148365685086094, 0.00148365685086072, 
    0.00148365685086094, 0.00148365685086094, 0.00148365685086072, 
    0.00148365685086094, 0.00148365685086094, 0.00148365685086072, 
    0.00148365685086094, 0.00148365685086072, 0.00148365685086094, 
    0.00148365685086094, 0.00148365685086094, 0.00148365685086094, 
    0.00148365685086094, 0.00148365685086094,
  0.00149818813682301, 0.00149818813682301, 0.00149818813682301, 
    0.00149818813682256, 0.00149818813682301, 0.00149818813682279, 
    0.00149818813682279, 0.00149818813682301, 0.00149818813682279, 
    0.00149818813682279, 0.00149818813682279, 0.00149818813682301, 
    0.00149818813682256, 0.00149818813682279, 0.00149818813682301, 
    0.00149818813682256, 0.00149818813682301, 0.00149818813682301, 
    0.00149818813682279, 0.00149818813682279, 0.00149818813682279, 
    0.00149818813682301, 0.00149818813682279, 0.00149818813682279, 
    0.00149818813682279, 0.00149818813682279, 0.00149818813682279, 
    0.00149818813682279, 0.00149818813682279, 0.00149818813682279, 
    0.00149818813682279, 0.00149818813682279, 0.00149818813682279, 
    0.00149818813682301, 0.00149818813682279, 0.00149818813682279, 
    0.00149818813682301, 0.00149818813682279, 0.00149818813682279, 
    0.00149818813682279, 0.00149818813682279, 0.00149818813682279, 
    0.00149818813682279, 0.00149818813682279, 0.00149818813682279, 
    0.00149818813682301, 0.00149818813682279, 0.00149818813682279, 
    0.00149818813682301, 0.00149818813682279, 0.00149818813682279, 
    0.00149818813682279, 0.00149818813682279, 0.00149818813682279, 
    0.00149818813682279, 0.00149818813682279,
  0.00151266871408717, 0.00151266871408717, 0.00151266871408717, 
    0.00151266871408695, 0.00151266871408717, 0.00151266871408717, 
    0.00151266871408695, 0.00151266871408717, 0.00151266871408717, 
    0.00151266871408695, 0.00151266871408717, 0.00151266871408717, 
    0.00151266871408695, 0.00151266871408717, 0.00151266871408717, 
    0.00151266871408695, 0.00151266871408717, 0.00151266871408717, 
    0.00151266871408695, 0.00151266871408717, 0.00151266871408695, 
    0.00151266871408717, 0.00151266871408695, 0.00151266871408717, 
    0.00151266871408717, 0.00151266871408717, 0.00151266871408717, 
    0.00151266871408717, 0.00151266871408695, 0.00151266871408717, 
    0.00151266871408717, 0.00151266871408717, 0.00151266871408695, 
    0.00151266871408717, 0.00151266871408695, 0.00151266871408717, 
    0.00151266871408717, 0.00151266871408695, 0.00151266871408717, 
    0.00151266871408717, 0.00151266871408717, 0.00151266871408695, 
    0.00151266871408717, 0.00151266871408717, 0.00151266871408695, 
    0.00151266871408717, 0.00151266871408717, 0.00151266871408695, 
    0.00151266871408717, 0.00151266871408695, 0.00151266871408717, 
    0.00151266871408717, 0.00151266871408717, 0.00151266871408717, 
    0.00151266871408717, 0.00151266871408717,
  0.00152709809263119, 0.00152709809263119, 0.00152709809263119, 
    0.00152709809263074, 0.00152709809263119, 0.00152709809263096, 
    0.00152709809263096, 0.00152709809263119, 0.00152709809263096, 
    0.00152709809263096, 0.00152709809263096, 0.00152709809263119, 
    0.00152709809263074, 0.00152709809263096, 0.00152709809263119, 
    0.00152709809263074, 0.00152709809263119, 0.00152709809263119, 
    0.00152709809263096, 0.00152709809263096, 0.00152709809263096, 
    0.00152709809263119, 0.00152709809263096, 0.00152709809263096, 
    0.00152709809263096, 0.00152709809263096, 0.00152709809263096, 
    0.00152709809263096, 0.00152709809263096, 0.00152709809263096, 
    0.00152709809263096, 0.00152709809263096, 0.00152709809263096, 
    0.00152709809263119, 0.00152709809263096, 0.00152709809263096, 
    0.00152709809263119, 0.00152709809263096, 0.00152709809263096, 
    0.00152709809263096, 0.00152709809263096, 0.00152709809263096, 
    0.00152709809263096, 0.00152709809263096, 0.00152709809263096, 
    0.00152709809263119, 0.00152709809263096, 0.00152709809263096, 
    0.00152709809263119, 0.00152709809263096, 0.00152709809263096, 
    0.00152709809263096, 0.00152709809263096, 0.00152709809263096, 
    0.00152709809263096, 0.00152709809263096,
  0.00154147578395847, 0.00154147578395847, 0.00154147578395847, 
    0.00154147578395825, 0.00154147578395847, 0.00154147578395847, 
    0.00154147578395825, 0.00154147578395847, 0.00154147578395847, 
    0.00154147578395825, 0.00154147578395847, 0.00154147578395847, 
    0.00154147578395825, 0.00154147578395847, 0.00154147578395847, 
    0.00154147578395825, 0.00154147578395847, 0.00154147578395847, 
    0.00154147578395825, 0.00154147578395847, 0.00154147578395825, 
    0.00154147578395847, 0.00154147578395825, 0.00154147578395847, 
    0.00154147578395847, 0.00154147578395847, 0.00154147578395847, 
    0.00154147578395847, 0.00154147578395825, 0.00154147578395847, 
    0.00154147578395847, 0.00154147578395847, 0.00154147578395825, 
    0.00154147578395847, 0.00154147578395825, 0.00154147578395847, 
    0.00154147578395847, 0.00154147578395825, 0.00154147578395847, 
    0.00154147578395847, 0.00154147578395847, 0.00154147578395825, 
    0.00154147578395847, 0.00154147578395847, 0.00154147578395825, 
    0.00154147578395847, 0.00154147578395847, 0.00154147578395825, 
    0.00154147578395847, 0.00154147578395825, 0.00154147578395847, 
    0.00154147578395847, 0.00154147578395847, 0.00154147578395847, 
    0.00154147578395847, 0.00154147578395847,
  0.00155580130157773, 0.00155580130157773, 0.00155580130157773, 
    0.00155580130157729, 0.00155580130157773, 0.00155580130157751, 
    0.00155580130157751, 0.00155580130157773, 0.00155580130157751, 
    0.00155580130157751, 0.00155580130157751, 0.00155580130157773, 
    0.00155580130157729, 0.00155580130157751, 0.00155580130157773, 
    0.00155580130157729, 0.00155580130157773, 0.00155580130157773, 
    0.00155580130157751, 0.00155580130157751, 0.00155580130157751, 
    0.00155580130157773, 0.00155580130157751, 0.00155580130157751, 
    0.00155580130157751, 0.00155580130157751, 0.00155580130157751, 
    0.00155580130157751, 0.00155580130157751, 0.00155580130157751, 
    0.00155580130157751, 0.00155580130157751, 0.00155580130157751, 
    0.00155580130157773, 0.00155580130157751, 0.00155580130157751, 
    0.00155580130157773, 0.00155580130157751, 0.00155580130157751, 
    0.00155580130157751, 0.00155580130157751, 0.00155580130157751, 
    0.00155580130157751, 0.00155580130157751, 0.00155580130157751, 
    0.00155580130157773, 0.00155580130157751, 0.00155580130157751, 
    0.00155580130157773, 0.00155580130157751, 0.00155580130157751, 
    0.00155580130157751, 0.00155580130157751, 0.00155580130157751, 
    0.00155580130157751, 0.00155580130157751,
  0.00157007416050425, 0.00157007416050425, 0.00157007416050425, 
    0.00157007416050403, 0.00157007416050425, 0.00157007416050425, 
    0.00157007416050403, 0.00157007416050425, 0.00157007416050425, 
    0.00157007416050403, 0.00157007416050425, 0.00157007416050425, 
    0.00157007416050403, 0.00157007416050425, 0.00157007416050425, 
    0.00157007416050403, 0.00157007416050425, 0.00157007416050425, 
    0.00157007416050403, 0.00157007416050425, 0.00157007416050403, 
    0.00157007416050425, 0.00157007416050403, 0.00157007416050425, 
    0.00157007416050425, 0.00157007416050425, 0.00157007416050425, 
    0.00157007416050425, 0.00157007416050403, 0.00157007416050425, 
    0.00157007416050425, 0.00157007416050425, 0.00157007416050403, 
    0.00157007416050425, 0.00157007416050403, 0.00157007416050425, 
    0.00157007416050425, 0.00157007416050403, 0.00157007416050425, 
    0.00157007416050425, 0.00157007416050425, 0.00157007416050403, 
    0.00157007416050425, 0.00157007416050425, 0.00157007416050403, 
    0.00157007416050425, 0.00157007416050425, 0.00157007416050403, 
    0.00157007416050425, 0.00157007416050403, 0.00157007416050425, 
    0.00157007416050425, 0.00157007416050425, 0.00157007416050425, 
    0.00157007416050425, 0.00157007416050425,
  0.00158429387772019, 0.00158429387772019, 0.00158429387772019, 
    0.00158429387771974, 0.00158429387772019, 0.00158429387771997, 
    0.00158429387771997, 0.00158429387772019, 0.00158429387771997, 
    0.00158429387771997, 0.00158429387771997, 0.00158429387772019, 
    0.00158429387771974, 0.00158429387771997, 0.00158429387772019, 
    0.00158429387771974, 0.00158429387772019, 0.00158429387772019, 
    0.00158429387771997, 0.00158429387771997, 0.00158429387771997, 
    0.00158429387772019, 0.00158429387771997, 0.00158429387771997, 
    0.00158429387771997, 0.00158429387771997, 0.00158429387771997, 
    0.00158429387771997, 0.00158429387771997, 0.00158429387771997, 
    0.00158429387771997, 0.00158429387771997, 0.00158429387771997, 
    0.00158429387772019, 0.00158429387771997, 0.00158429387771997, 
    0.00158429387772019, 0.00158429387771997, 0.00158429387771997, 
    0.00158429387771997, 0.00158429387771997, 0.00158429387771997, 
    0.00158429387771997, 0.00158429387771997, 0.00158429387771997, 
    0.00158429387772019, 0.00158429387771997, 0.00158429387771997, 
    0.00158429387772019, 0.00158429387771997, 0.00158429387771997, 
    0.00158429387771997, 0.00158429387771997, 0.00158429387771997, 
    0.00158429387771997, 0.00158429387771997,
  0.00159845997192432, 0.00159845997192432, 0.00159845997192432, 
    0.00159845997192387, 0.00159845997192432, 0.00159845997192409, 
    0.00159845997192409, 0.00159845997192432, 0.00159845997192409, 
    0.00159845997192409, 0.00159845997192409, 0.00159845997192432, 
    0.00159845997192387, 0.00159845997192409, 0.00159845997192432, 
    0.00159845997192387, 0.00159845997192432, 0.00159845997192432, 
    0.00159845997192409, 0.00159845997192409, 0.00159845997192409, 
    0.00159845997192432, 0.00159845997192409, 0.00159845997192409, 
    0.00159845997192409, 0.00159845997192409, 0.00159845997192409, 
    0.00159845997192409, 0.00159845997192409, 0.00159845997192409, 
    0.00159845997192409, 0.00159845997192409, 0.00159845997192409, 
    0.00159845997192432, 0.00159845997192409, 0.00159845997192409, 
    0.00159845997192432, 0.00159845997192409, 0.00159845997192409, 
    0.00159845997192409, 0.00159845997192409, 0.00159845997192409, 
    0.00159845997192409, 0.00159845997192409, 0.00159845997192409, 
    0.00159845997192432, 0.00159845997192409, 0.00159845997192409, 
    0.00159845997192432, 0.00159845997192409, 0.00159845997192409, 
    0.00159845997192409, 0.00159845997192409, 0.00159845997192409, 
    0.00159845997192409, 0.00159845997192409,
  0.00161257196366749, 0.00161257196366749, 0.00161257196366749, 
    0.00161257196366704, 0.00161257196366749, 0.00161257196366726, 
    0.00161257196366726, 0.00161257196366749, 0.00161257196366726, 
    0.00161257196366726, 0.00161257196366726, 0.00161257196366749, 
    0.00161257196366704, 0.00161257196366726, 0.00161257196366749, 
    0.00161257196366704, 0.00161257196366749, 0.00161257196366749, 
    0.00161257196366726, 0.00161257196366726, 0.00161257196366726, 
    0.00161257196366749, 0.00161257196366726, 0.00161257196366726, 
    0.00161257196366726, 0.00161257196366726, 0.00161257196366726, 
    0.00161257196366726, 0.00161257196366726, 0.00161257196366726, 
    0.00161257196366726, 0.00161257196366726, 0.00161257196366726, 
    0.00161257196366749, 0.00161257196366726, 0.00161257196366726, 
    0.00161257196366749, 0.00161257196366726, 0.00161257196366726, 
    0.00161257196366726, 0.00161257196366726, 0.00161257196366726, 
    0.00161257196366726, 0.00161257196366726, 0.00161257196366726, 
    0.00161257196366749, 0.00161257196366726, 0.00161257196366726, 
    0.00161257196366749, 0.00161257196366726, 0.00161257196366726, 
    0.00161257196366726, 0.00161257196366726, 0.00161257196366726, 
    0.00161257196366726, 0.00161257196366726,
  0.00162662937527513, 0.00162662937527513, 0.00162662937527513, 
    0.00162662937527469, 0.00162662937527513, 0.00162662937527491, 
    0.00162662937527491, 0.00162662937527513, 0.00162662937527491, 
    0.00162662937527491, 0.00162662937527491, 0.00162662937527513, 
    0.00162662937527469, 0.00162662937527491, 0.00162662937527513, 
    0.00162662937527469, 0.00162662937527513, 0.00162662937527513, 
    0.00162662937527491, 0.00162662937527491, 0.00162662937527491, 
    0.00162662937527513, 0.00162662937527491, 0.00162662937527491, 
    0.00162662937527491, 0.00162662937527491, 0.00162662937527491, 
    0.00162662937527491, 0.00162662937527491, 0.00162662937527491, 
    0.00162662937527491, 0.00162662937527491, 0.00162662937527491, 
    0.00162662937527513, 0.00162662937527491, 0.00162662937527491, 
    0.00162662937527513, 0.00162662937527491, 0.00162662937527491, 
    0.00162662937527491, 0.00162662937527491, 0.00162662937527491, 
    0.00162662937527491, 0.00162662937527491, 0.00162662937527491, 
    0.00162662937527513, 0.00162662937527491, 0.00162662937527491, 
    0.00162662937527513, 0.00162662937527491, 0.00162662937527491, 
    0.00162662937527491, 0.00162662937527491, 0.00162662937527491, 
    0.00162662937527491, 0.00162662937527491,
  0.00164063173096207, 0.00164063173096207, 0.00164063173096207, 
    0.00164063173096185, 0.00164063173096207, 0.00164063173096207, 
    0.00164063173096185, 0.00164063173096207, 0.00164063173096207, 
    0.00164063173096185, 0.00164063173096207, 0.00164063173096207, 
    0.00164063173096185, 0.00164063173096207, 0.00164063173096207, 
    0.00164063173096185, 0.00164063173096207, 0.00164063173096207, 
    0.00164063173096185, 0.00164063173096207, 0.00164063173096185, 
    0.00164063173096207, 0.00164063173096185, 0.00164063173096207, 
    0.00164063173096207, 0.00164063173096207, 0.00164063173096207, 
    0.00164063173096207, 0.00164063173096185, 0.00164063173096207, 
    0.00164063173096207, 0.00164063173096207, 0.00164063173096185, 
    0.00164063173096207, 0.00164063173096185, 0.00164063173096207, 
    0.00164063173096207, 0.00164063173096185, 0.00164063173096207, 
    0.00164063173096207, 0.00164063173096207, 0.00164063173096185, 
    0.00164063173096207, 0.00164063173096207, 0.00164063173096185, 
    0.00164063173096207, 0.00164063173096207, 0.00164063173096185, 
    0.00164063173096207, 0.00164063173096185, 0.00164063173096207, 
    0.00164063173096207, 0.00164063173096207, 0.00164063173096207, 
    0.00164063173096207, 0.00164063173096207,
  0.00165457855685225, 0.00165457855685225, 0.00165457855685225, 
    0.0016545785568518, 0.00165457855685225, 0.00165457855685203, 
    0.00165457855685203, 0.00165457855685225, 0.00165457855685203, 
    0.00165457855685203, 0.00165457855685203, 0.00165457855685225, 
    0.0016545785568518, 0.00165457855685203, 0.00165457855685225, 
    0.0016545785568518, 0.00165457855685225, 0.00165457855685225, 
    0.00165457855685203, 0.00165457855685203, 0.00165457855685203, 
    0.00165457855685225, 0.00165457855685203, 0.00165457855685203, 
    0.00165457855685203, 0.00165457855685203, 0.00165457855685203, 
    0.00165457855685203, 0.00165457855685203, 0.00165457855685203, 
    0.00165457855685203, 0.00165457855685203, 0.00165457855685203, 
    0.00165457855685225, 0.00165457855685203, 0.00165457855685203, 
    0.00165457855685225, 0.00165457855685203, 0.00165457855685203, 
    0.00165457855685203, 0.00165457855685203, 0.00165457855685203, 
    0.00165457855685203, 0.00165457855685203, 0.00165457855685203, 
    0.00165457855685225, 0.00165457855685203, 0.00165457855685203, 
    0.00165457855685225, 0.00165457855685203, 0.00165457855685203, 
    0.00165457855685203, 0.00165457855685203, 0.00165457855685203, 
    0.00165457855685203, 0.00165457855685203,
  0.00166846938086262, 0.00166846938086262, 0.00166846938086262, 
    0.0016684693808624, 0.00166846938086262, 0.00166846938086262, 
    0.0016684693808624, 0.00166846938086262, 0.00166846938086262, 
    0.0016684693808624, 0.00166846938086262, 0.00166846938086262, 
    0.0016684693808624, 0.00166846938086262, 0.00166846938086262, 
    0.0016684693808624, 0.00166846938086262, 0.00166846938086262, 
    0.0016684693808624, 0.00166846938086262, 0.0016684693808624, 
    0.00166846938086262, 0.0016684693808624, 0.00166846938086262, 
    0.00166846938086262, 0.00166846938086262, 0.00166846938086262, 
    0.00166846938086262, 0.0016684693808624, 0.00166846938086262, 
    0.00166846938086262, 0.00166846938086262, 0.0016684693808624, 
    0.00166846938086262, 0.0016684693808624, 0.00166846938086262, 
    0.00166846938086262, 0.0016684693808624, 0.00166846938086262, 
    0.00166846938086262, 0.00166846938086262, 0.0016684693808624, 
    0.00166846938086262, 0.00166846938086262, 0.0016684693808624, 
    0.00166846938086262, 0.00166846938086262, 0.0016684693808624, 
    0.00166846938086262, 0.0016684693808624, 0.00166846938086262, 
    0.00166846938086262, 0.00166846938086262, 0.00166846938086262, 
    0.00166846938086262, 0.00166846938086262,
  0.00168230373285794, 0.00168230373285794, 0.00168230373285794, 
    0.00168230373285749, 0.00168230373285794, 0.00168230373285772, 
    0.00168230373285772, 0.00168230373285794, 0.00168230373285772, 
    0.00168230373285772, 0.00168230373285772, 0.00168230373285794, 
    0.00168230373285749, 0.00168230373285772, 0.00168230373285794, 
    0.00168230373285749, 0.00168230373285794, 0.00168230373285794, 
    0.00168230373285772, 0.00168230373285772, 0.00168230373285772, 
    0.00168230373285794, 0.00168230373285772, 0.00168230373285772, 
    0.00168230373285772, 0.00168230373285772, 0.00168230373285772, 
    0.00168230373285772, 0.00168230373285772, 0.00168230373285772, 
    0.00168230373285772, 0.00168230373285772, 0.00168230373285772, 
    0.00168230373285794, 0.00168230373285772, 0.00168230373285772, 
    0.00168230373285794, 0.00168230373285772, 0.00168230373285772, 
    0.00168230373285772, 0.00168230373285772, 0.00168230373285772, 
    0.00168230373285772, 0.00168230373285772, 0.00168230373285772, 
    0.00168230373285794, 0.00168230373285772, 0.00168230373285772, 
    0.00168230373285794, 0.00168230373285772, 0.00168230373285772, 
    0.00168230373285772, 0.00168230373285772, 0.00168230373285772, 
    0.00168230373285772, 0.00168230373285772,
  0.00169608114455322, 0.00169608114455322, 0.00169608114455322, 
    0.00169608114455277, 0.00169608114455322, 0.001696081144553, 
    0.001696081144553, 0.00169608114455322, 0.001696081144553, 
    0.001696081144553, 0.001696081144553, 0.00169608114455322, 
    0.00169608114455277, 0.001696081144553, 0.00169608114455322, 
    0.00169608114455277, 0.00169608114455322, 0.00169608114455322, 
    0.001696081144553, 0.001696081144553, 0.001696081144553, 
    0.00169608114455322, 0.001696081144553, 0.001696081144553, 
    0.001696081144553, 0.001696081144553, 0.001696081144553, 
    0.001696081144553, 0.001696081144553, 0.001696081144553, 
    0.001696081144553, 0.001696081144553, 0.001696081144553, 
    0.00169608114455322, 0.001696081144553, 0.001696081144553, 
    0.00169608114455322, 0.001696081144553, 0.001696081144553, 
    0.001696081144553, 0.001696081144553, 0.001696081144553, 
    0.001696081144553, 0.001696081144553, 0.001696081144553, 
    0.00169608114455322, 0.001696081144553, 0.001696081144553, 
    0.00169608114455322, 0.001696081144553, 0.001696081144553, 
    0.001696081144553, 0.001696081144553, 0.001696081144553, 
    0.001696081144553, 0.001696081144553,
  0.00170980114970609, 0.00170980114970609, 0.00170980114970609, 
    0.00170980114970587, 0.00170980114970609, 0.00170980114970609, 
    0.00170980114970587, 0.00170980114970609, 0.00170980114970609, 
    0.00170980114970587, 0.00170980114970609, 0.00170980114970609, 
    0.00170980114970587, 0.00170980114970609, 0.00170980114970609, 
    0.00170980114970587, 0.00170980114970609, 0.00170980114970609, 
    0.00170980114970587, 0.00170980114970609, 0.00170980114970587, 
    0.00170980114970609, 0.00170980114970587, 0.00170980114970609, 
    0.00170980114970609, 0.00170980114970609, 0.00170980114970609, 
    0.00170980114970609, 0.00170980114970587, 0.00170980114970609, 
    0.00170980114970609, 0.00170980114970609, 0.00170980114970587, 
    0.00170980114970609, 0.00170980114970587, 0.00170980114970609, 
    0.00170980114970609, 0.00170980114970587, 0.00170980114970609, 
    0.00170980114970609, 0.00170980114970609, 0.00170980114970587, 
    0.00170980114970609, 0.00170980114970609, 0.00170980114970587, 
    0.00170980114970609, 0.00170980114970609, 0.00170980114970587, 
    0.00170980114970609, 0.00170980114970587, 0.00170980114970609, 
    0.00170980114970609, 0.00170980114970609, 0.00170980114970609, 
    0.00170980114970609, 0.00170980114970609,
  0.00172346328388762, 0.00172346328388762, 0.00172346328388762, 
    0.00172346328388717, 0.00172346328388762, 0.00172346328388739, 
    0.00172346328388739, 0.00172346328388762, 0.00172346328388739, 
    0.00172346328388739, 0.00172346328388739, 0.00172346328388762, 
    0.00172346328388717, 0.00172346328388739, 0.00172346328388762, 
    0.00172346328388717, 0.00172346328388762, 0.00172346328388762, 
    0.00172346328388739, 0.00172346328388739, 0.00172346328388739, 
    0.00172346328388762, 0.00172346328388739, 0.00172346328388739, 
    0.00172346328388739, 0.00172346328388739, 0.00172346328388739, 
    0.00172346328388739, 0.00172346328388739, 0.00172346328388739, 
    0.00172346328388739, 0.00172346328388739, 0.00172346328388739, 
    0.00172346328388762, 0.00172346328388739, 0.00172346328388739, 
    0.00172346328388762, 0.00172346328388739, 0.00172346328388739, 
    0.00172346328388739, 0.00172346328388739, 0.00172346328388739, 
    0.00172346328388739, 0.00172346328388739, 0.00172346328388739, 
    0.00172346328388762, 0.00172346328388739, 0.00172346328388739, 
    0.00172346328388762, 0.00172346328388739, 0.00172346328388739, 
    0.00172346328388739, 0.00172346328388739, 0.00172346328388739, 
    0.00172346328388739, 0.00172346328388739,
  0.0017370670847483, 0.0017370670847483, 0.0017370670847483, 
    0.00173706708474808, 0.0017370670847483, 0.0017370670847483, 
    0.00173706708474808, 0.0017370670847483, 0.0017370670847483, 
    0.00173706708474808, 0.0017370670847483, 0.0017370670847483, 
    0.00173706708474808, 0.0017370670847483, 0.0017370670847483, 
    0.00173706708474808, 0.0017370670847483, 0.0017370670847483, 
    0.00173706708474808, 0.0017370670847483, 0.00173706708474808, 
    0.0017370670847483, 0.00173706708474808, 0.0017370670847483, 
    0.0017370670847483, 0.0017370670847483, 0.0017370670847483, 
    0.0017370670847483, 0.00173706708474808, 0.0017370670847483, 
    0.0017370670847483, 0.0017370670847483, 0.00173706708474808, 
    0.0017370670847483, 0.00173706708474808, 0.0017370670847483, 
    0.0017370670847483, 0.00173706708474808, 0.0017370670847483, 
    0.0017370670847483, 0.0017370670847483, 0.00173706708474808, 
    0.0017370670847483, 0.0017370670847483, 0.00173706708474808, 
    0.0017370670847483, 0.0017370670847483, 0.00173706708474808, 
    0.0017370670847483, 0.00173706708474808, 0.0017370670847483, 
    0.0017370670847483, 0.0017370670847483, 0.0017370670847483, 
    0.0017370670847483, 0.0017370670847483,
  0.00175061209179073, 0.00175061209179073, 0.00175061209179073, 
    0.00175061209179028, 0.00175061209179073, 0.0017506120917905, 
    0.0017506120917905, 0.00175061209179073, 0.0017506120917905, 
    0.0017506120917905, 0.0017506120917905, 0.00175061209179073, 
    0.00175061209179028, 0.0017506120917905, 0.00175061209179073, 
    0.00175061209179028, 0.00175061209179073, 0.00175061209179073, 
    0.0017506120917905, 0.0017506120917905, 0.0017506120917905, 
    0.00175061209179073, 0.0017506120917905, 0.0017506120917905, 
    0.0017506120917905, 0.0017506120917905, 0.0017506120917905, 
    0.0017506120917905, 0.0017506120917905, 0.0017506120917905, 
    0.0017506120917905, 0.0017506120917905, 0.0017506120917905, 
    0.00175061209179073, 0.0017506120917905, 0.0017506120917905, 
    0.00175061209179073, 0.0017506120917905, 0.0017506120917905, 
    0.0017506120917905, 0.0017506120917905, 0.0017506120917905, 
    0.0017506120917905, 0.0017506120917905, 0.0017506120917905, 
    0.00175061209179073, 0.0017506120917905, 0.0017506120917905, 
    0.00175061209179073, 0.0017506120917905, 0.0017506120917905, 
    0.0017506120917905, 0.0017506120917905, 0.0017506120917905, 
    0.0017506120917905, 0.0017506120917905,
  0.00176409784661624, 0.00176409784661624, 0.00176409784661624, 
    0.0017640978466158, 0.00176409784661624, 0.00176409784661624, 
    0.00176409784661602, 0.00176409784661624, 0.00176409784661624, 
    0.00176409784661602, 0.00176409784661624, 0.00176409784661624, 
    0.0017640978466158, 0.00176409784661624, 0.00176409784661624, 
    0.0017640978466158, 0.00176409784661624, 0.00176409784661624, 
    0.00176409784661602, 0.00176409784661624, 0.00176409784661602, 
    0.00176409784661624, 0.00176409784661602, 0.00176409784661624, 
    0.00176409784661624, 0.00176409784661624, 0.00176409784661624, 
    0.00176409784661624, 0.00176409784661602, 0.00176409784661624, 
    0.00176409784661624, 0.00176409784661624, 0.00176409784661602, 
    0.00176409784661624, 0.00176409784661602, 0.00176409784661624, 
    0.00176409784661624, 0.00176409784661602, 0.00176409784661624, 
    0.00176409784661624, 0.00176409784661624, 0.00176409784661602, 
    0.00176409784661624, 0.00176409784661624, 0.00176409784661602, 
    0.00176409784661624, 0.00176409784661624, 0.00176409784661602, 
    0.00176409784661624, 0.00176409784661602, 0.00176409784661624, 
    0.00176409784661624, 0.00176409784661624, 0.00176409784661624, 
    0.00176409784661624, 0.00176409784661624,
  0.00177752389275421, 0.00177752389275421, 0.00177752389275421, 
    0.00177752389275376, 0.00177752389275421, 0.00177752389275398, 
    0.00177752389275376, 0.00177752389275421, 0.00177752389275398, 
    0.00177752389275376, 0.00177752389275398, 0.00177752389275421, 
    0.00177752389275376, 0.00177752389275398, 0.00177752389275421, 
    0.00177752389275376, 0.00177752389275421, 0.00177752389275421, 
    0.00177752389275376, 0.00177752389275398, 0.00177752389275376, 
    0.00177752389275421, 0.00177752389275376, 0.00177752389275398, 
    0.00177752389275398, 0.00177752389275398, 0.00177752389275398, 
    0.00177752389275398, 0.00177752389275376, 0.00177752389275398, 
    0.00177752389275398, 0.00177752389275398, 0.00177752389275376, 
    0.00177752389275421, 0.00177752389275376, 0.00177752389275398, 
    0.00177752389275421, 0.00177752389275376, 0.00177752389275398, 
    0.00177752389275398, 0.00177752389275398, 0.00177752389275376, 
    0.00177752389275398, 0.00177752389275398, 0.00177752389275376, 
    0.00177752389275421, 0.00177752389275398, 0.00177752389275376, 
    0.00177752389275421, 0.00177752389275376, 0.00177752389275398, 
    0.00177752389275398, 0.00177752389275398, 0.00177752389275398, 
    0.00177752389275398, 0.00177752389275398,
  0.00179088977585207, 0.00179088977585207, 0.00179088977585207, 
    0.00179088977585162, 0.00179088977585207, 0.00179088977585184, 
    0.00179088977585162, 0.00179088977585207, 0.00179088977585184, 
    0.00179088977585162, 0.00179088977585184, 0.00179088977585207, 
    0.00179088977585162, 0.00179088977585184, 0.00179088977585207, 
    0.00179088977585162, 0.00179088977585207, 0.00179088977585207, 
    0.00179088977585162, 0.00179088977585184, 0.00179088977585162, 
    0.00179088977585207, 0.00179088977585162, 0.00179088977585184, 
    0.00179088977585184, 0.00179088977585184, 0.00179088977585184, 
    0.00179088977585184, 0.00179088977585162, 0.00179088977585184, 
    0.00179088977585184, 0.00179088977585184, 0.00179088977585162, 
    0.00179088977585207, 0.00179088977585162, 0.00179088977585184, 
    0.00179088977585207, 0.00179088977585162, 0.00179088977585184, 
    0.00179088977585184, 0.00179088977585184, 0.00179088977585162, 
    0.00179088977585184, 0.00179088977585184, 0.00179088977585162, 
    0.00179088977585207, 0.00179088977585184, 0.00179088977585162, 
    0.00179088977585207, 0.00179088977585162, 0.00179088977585184, 
    0.00179088977585184, 0.00179088977585184, 0.00179088977585184, 
    0.00179088977585184, 0.00179088977585184,
  0.00180419504342777, 0.00180419504342777, 0.00180419504342777, 
    0.00180419504342733, 0.00180419504342777, 0.00180419504342755, 
    0.00180419504342733, 0.00180419504342777, 0.00180419504342755, 
    0.00180419504342733, 0.00180419504342755, 0.00180419504342777, 
    0.00180419504342733, 0.00180419504342755, 0.00180419504342777, 
    0.00180419504342733, 0.00180419504342777, 0.00180419504342777, 
    0.00180419504342733, 0.00180419504342755, 0.00180419504342733, 
    0.00180419504342777, 0.00180419504342733, 0.00180419504342755, 
    0.00180419504342755, 0.00180419504342755, 0.00180419504342755, 
    0.00180419504342755, 0.00180419504342733, 0.00180419504342755, 
    0.00180419504342755, 0.00180419504342755, 0.00180419504342733, 
    0.00180419504342777, 0.00180419504342733, 0.00180419504342755, 
    0.00180419504342777, 0.00180419504342733, 0.00180419504342755, 
    0.00180419504342755, 0.00180419504342755, 0.00180419504342733, 
    0.00180419504342755, 0.00180419504342755, 0.00180419504342733, 
    0.00180419504342777, 0.00180419504342755, 0.00180419504342733, 
    0.00180419504342777, 0.00180419504342733, 0.00180419504342755, 
    0.00180419504342755, 0.00180419504342755, 0.00180419504342755, 
    0.00180419504342755, 0.00180419504342755,
  0.00181743924519417, 0.00181743924519417, 0.00181743924519417, 
    0.00181743924519373, 0.00181743924519417, 0.00181743924519395, 
    0.00181743924519373, 0.00181743924519417, 0.00181743924519395, 
    0.00181743924519373, 0.00181743924519395, 0.00181743924519417, 
    0.00181743924519373, 0.00181743924519395, 0.00181743924519417, 
    0.00181743924519373, 0.00181743924519417, 0.00181743924519417, 
    0.00181743924519373, 0.00181743924519395, 0.00181743924519373, 
    0.00181743924519417, 0.00181743924519373, 0.00181743924519395, 
    0.00181743924519395, 0.00181743924519395, 0.00181743924519395, 
    0.00181743924519395, 0.00181743924519373, 0.00181743924519395, 
    0.00181743924519395, 0.00181743924519395, 0.00181743924519373, 
    0.00181743924519417, 0.00181743924519373, 0.00181743924519395, 
    0.00181743924519417, 0.00181743924519373, 0.00181743924519395, 
    0.00181743924519395, 0.00181743924519395, 0.00181743924519373, 
    0.00181743924519395, 0.00181743924519395, 0.00181743924519373, 
    0.00181743924519417, 0.00181743924519395, 0.00181743924519373, 
    0.00181743924519417, 0.00181743924519373, 0.00181743924519395, 
    0.00181743924519395, 0.00181743924519395, 0.00181743924519395, 
    0.00181743924519395, 0.00181743924519395,
  0.00183062193290584, 0.00183062193290584, 0.00183062193290584, 
    0.00183062193290562, 0.00183062193290584, 0.00183062193290584, 
    0.00183062193290562, 0.00183062193290584, 0.00183062193290584, 
    0.00183062193290562, 0.00183062193290584, 0.00183062193290584, 
    0.00183062193290562, 0.00183062193290584, 0.00183062193290584, 
    0.00183062193290562, 0.00183062193290584, 0.00183062193290584, 
    0.00183062193290562, 0.00183062193290584, 0.00183062193290562, 
    0.00183062193290584, 0.00183062193290562, 0.00183062193290584, 
    0.00183062193290584, 0.00183062193290584, 0.00183062193290584, 
    0.00183062193290584, 0.00183062193290562, 0.00183062193290584, 
    0.00183062193290584, 0.00183062193290584, 0.00183062193290562, 
    0.00183062193290584, 0.00183062193290562, 0.00183062193290584, 
    0.00183062193290584, 0.00183062193290562, 0.00183062193290584, 
    0.00183062193290584, 0.00183062193290584, 0.00183062193290562, 
    0.00183062193290584, 0.00183062193290584, 0.00183062193290562, 
    0.00183062193290584, 0.00183062193290584, 0.00183062193290562, 
    0.00183062193290584, 0.00183062193290562, 0.00183062193290584, 
    0.00183062193290584, 0.00183062193290584, 0.00183062193290584, 
    0.00183062193290584, 0.00183062193290584,
  0.00184374266037923, 0.00184374266037923, 0.00184374266037923, 
    0.00184374266037879, 0.00184374266037923, 0.00184374266037901, 
    0.00184374266037901, 0.00184374266037923, 0.00184374266037901, 
    0.00184374266037901, 0.00184374266037901, 0.00184374266037923, 
    0.00184374266037879, 0.00184374266037901, 0.00184374266037923, 
    0.00184374266037879, 0.00184374266037923, 0.00184374266037923, 
    0.00184374266037901, 0.00184374266037901, 0.00184374266037901, 
    0.00184374266037923, 0.00184374266037901, 0.00184374266037901, 
    0.00184374266037901, 0.00184374266037901, 0.00184374266037901, 
    0.00184374266037901, 0.00184374266037901, 0.00184374266037901, 
    0.00184374266037901, 0.00184374266037901, 0.00184374266037901, 
    0.00184374266037923, 0.00184374266037901, 0.00184374266037901, 
    0.00184374266037923, 0.00184374266037901, 0.00184374266037901, 
    0.00184374266037901, 0.00184374266037901, 0.00184374266037901, 
    0.00184374266037901, 0.00184374266037901, 0.00184374266037901, 
    0.00184374266037923, 0.00184374266037901, 0.00184374266037901, 
    0.00184374266037923, 0.00184374266037901, 0.00184374266037901, 
    0.00184374266037901, 0.00184374266037901, 0.00184374266037901, 
    0.00184374266037901, 0.00184374266037901,
  0.00185680098351027, 0.00185680098351027, 0.00185680098351027, 
    0.00185680098350982, 0.00185680098351027, 0.00185680098351004, 
    0.00185680098351004, 0.00185680098351027, 0.00185680098351004, 
    0.00185680098351004, 0.00185680098351004, 0.00185680098351027, 
    0.00185680098350982, 0.00185680098351004, 0.00185680098351027, 
    0.00185680098350982, 0.00185680098351027, 0.00185680098351027, 
    0.00185680098351004, 0.00185680098351004, 0.00185680098351004, 
    0.00185680098351027, 0.00185680098351004, 0.00185680098351004, 
    0.00185680098351004, 0.00185680098351004, 0.00185680098351004, 
    0.00185680098351004, 0.00185680098351004, 0.00185680098351004, 
    0.00185680098351004, 0.00185680098351004, 0.00185680098351004, 
    0.00185680098351027, 0.00185680098351004, 0.00185680098351004, 
    0.00185680098351027, 0.00185680098351004, 0.00185680098351004, 
    0.00185680098351004, 0.00185680098351004, 0.00185680098351004, 
    0.00185680098351004, 0.00185680098351004, 0.00185680098351004, 
    0.00185680098351027, 0.00185680098351004, 0.00185680098351004, 
    0.00185680098351027, 0.00185680098351004, 0.00185680098351004, 
    0.00185680098351004, 0.00185680098351004, 0.00185680098351004, 
    0.00185680098351004, 0.00185680098351004,
  0.00186979646035179, 0.00186979646035179, 0.00186979646035179, 
    0.00186979646035135, 0.00186979646035179, 0.00186979646035179, 
    0.00186979646035157, 0.00186979646035179, 0.00186979646035179, 
    0.00186979646035157, 0.00186979646035179, 0.00186979646035179, 
    0.00186979646035135, 0.00186979646035179, 0.00186979646035179, 
    0.00186979646035135, 0.00186979646035179, 0.00186979646035179, 
    0.00186979646035157, 0.00186979646035179, 0.00186979646035157, 
    0.00186979646035179, 0.00186979646035157, 0.00186979646035179, 
    0.00186979646035179, 0.00186979646035179, 0.00186979646035179, 
    0.00186979646035179, 0.00186979646035157, 0.00186979646035179, 
    0.00186979646035179, 0.00186979646035179, 0.00186979646035157, 
    0.00186979646035179, 0.00186979646035157, 0.00186979646035179, 
    0.00186979646035179, 0.00186979646035157, 0.00186979646035179, 
    0.00186979646035179, 0.00186979646035179, 0.00186979646035157, 
    0.00186979646035179, 0.00186979646035179, 0.00186979646035157, 
    0.00186979646035179, 0.00186979646035179, 0.00186979646035157, 
    0.00186979646035179, 0.00186979646035157, 0.00186979646035179, 
    0.00186979646035179, 0.00186979646035179, 0.00186979646035179, 
    0.00186979646035179, 0.00186979646035179,
  0.00188272865105632, 0.00188272865105632, 0.00188272865105632, 
    0.00188272865105588, 0.00188272865105632, 0.0018827286510561, 
    0.00188272865105588, 0.00188272865105632, 0.0018827286510561, 
    0.00188272865105588, 0.0018827286510561, 0.00188272865105632, 
    0.00188272865105588, 0.0018827286510561, 0.00188272865105632, 
    0.00188272865105588, 0.00188272865105632, 0.00188272865105632, 
    0.00188272865105588, 0.0018827286510561, 0.00188272865105588, 
    0.00188272865105632, 0.00188272865105588, 0.0018827286510561, 
    0.0018827286510561, 0.0018827286510561, 0.0018827286510561, 
    0.0018827286510561, 0.00188272865105588, 0.0018827286510561, 
    0.0018827286510561, 0.0018827286510561, 0.00188272865105588, 
    0.00188272865105632, 0.00188272865105588, 0.0018827286510561, 
    0.00188272865105632, 0.00188272865105588, 0.0018827286510561, 
    0.0018827286510561, 0.0018827286510561, 0.00188272865105588, 
    0.0018827286510561, 0.0018827286510561, 0.00188272865105588, 
    0.00188272865105632, 0.0018827286510561, 0.00188272865105588, 
    0.00188272865105632, 0.00188272865105588, 0.0018827286510561, 
    0.0018827286510561, 0.0018827286510561, 0.0018827286510561, 
    0.0018827286510561, 0.0018827286510561,
  0.00189559711795129, 0.00189559711795129, 0.00189559711795129, 
    0.00189559711795084, 0.00189559711795129, 0.00189559711795106, 
    0.00189559711795084, 0.00189559711795129, 0.00189559711795106, 
    0.00189559711795084, 0.00189559711795106, 0.00189559711795129, 
    0.00189559711795084, 0.00189559711795106, 0.00189559711795129, 
    0.00189559711795084, 0.00189559711795129, 0.00189559711795129, 
    0.00189559711795084, 0.00189559711795106, 0.00189559711795084, 
    0.00189559711795129, 0.00189559711795084, 0.00189559711795106, 
    0.00189559711795106, 0.00189559711795106, 0.00189559711795106, 
    0.00189559711795106, 0.00189559711795084, 0.00189559711795106, 
    0.00189559711795106, 0.00189559711795106, 0.00189559711795084, 
    0.00189559711795129, 0.00189559711795084, 0.00189559711795106, 
    0.00189559711795129, 0.00189559711795084, 0.00189559711795106, 
    0.00189559711795106, 0.00189559711795106, 0.00189559711795084, 
    0.00189559711795106, 0.00189559711795106, 0.00189559711795084, 
    0.00189559711795129, 0.00189559711795106, 0.00189559711795084, 
    0.00189559711795129, 0.00189559711795084, 0.00189559711795106, 
    0.00189559711795106, 0.00189559711795106, 0.00189559711795106, 
    0.00189559711795106, 0.00189559711795106,
  0.00190840142538762, 0.00190840142538762, 0.00190840142538762, 
    0.00190840142538717, 0.00190840142538762, 0.00190840142538762, 
    0.0019084014253874, 0.00190840142538762, 0.00190840142538762, 
    0.0019084014253874, 0.00190840142538762, 0.00190840142538762, 
    0.00190840142538717, 0.00190840142538762, 0.00190840142538762, 
    0.00190840142538717, 0.00190840142538762, 0.00190840142538762, 
    0.0019084014253874, 0.00190840142538762, 0.0019084014253874, 
    0.00190840142538762, 0.0019084014253874, 0.00190840142538762, 
    0.00190840142538762, 0.00190840142538762, 0.00190840142538762, 
    0.00190840142538762, 0.0019084014253874, 0.00190840142538762, 
    0.00190840142538762, 0.00190840142538762, 0.0019084014253874, 
    0.00190840142538762, 0.0019084014253874, 0.00190840142538762, 
    0.00190840142538762, 0.0019084014253874, 0.00190840142538762, 
    0.00190840142538762, 0.00190840142538762, 0.0019084014253874, 
    0.00190840142538762, 0.00190840142538762, 0.0019084014253874, 
    0.00190840142538762, 0.00190840142538762, 0.0019084014253874, 
    0.00190840142538762, 0.0019084014253874, 0.00190840142538762, 
    0.00190840142538762, 0.00190840142538762, 0.00190840142538762, 
    0.00190840142538762, 0.00190840142538762,
  0.00192114114012121, 0.00192114114012121, 0.00192114114012121, 
    0.00192114114012076, 0.00192114114012121, 0.00192114114012099, 
    0.00192114114012076, 0.00192114114012121, 0.00192114114012099, 
    0.00192114114012076, 0.00192114114012099, 0.00192114114012121, 
    0.00192114114012076, 0.00192114114012099, 0.00192114114012121, 
    0.00192114114012076, 0.00192114114012121, 0.00192114114012121, 
    0.00192114114012076, 0.00192114114012099, 0.00192114114012076, 
    0.00192114114012121, 0.00192114114012076, 0.00192114114012099, 
    0.00192114114012099, 0.00192114114012099, 0.00192114114012099, 
    0.00192114114012099, 0.00192114114012076, 0.00192114114012099, 
    0.00192114114012099, 0.00192114114012099, 0.00192114114012076, 
    0.00192114114012121, 0.00192114114012076, 0.00192114114012099, 
    0.00192114114012121, 0.00192114114012076, 0.00192114114012099, 
    0.00192114114012099, 0.00192114114012099, 0.00192114114012076, 
    0.00192114114012099, 0.00192114114012099, 0.00192114114012076, 
    0.00192114114012121, 0.00192114114012099, 0.00192114114012076, 
    0.00192114114012121, 0.00192114114012076, 0.00192114114012099, 
    0.00192114114012099, 0.00192114114012099, 0.00192114114012099, 
    0.00192114114012099, 0.00192114114012099,
  0.00193381583085395, 0.00193381583085395, 0.00193381583085395, 
    0.0019338158308535, 0.00193381583085395, 0.00193381583085372, 
    0.0019338158308535, 0.00193381583085395, 0.00193381583085372, 
    0.0019338158308535, 0.00193381583085372, 0.00193381583085395, 
    0.0019338158308535, 0.00193381583085372, 0.00193381583085395, 
    0.0019338158308535, 0.00193381583085395, 0.00193381583085395, 
    0.0019338158308535, 0.00193381583085372, 0.0019338158308535, 
    0.00193381583085395, 0.0019338158308535, 0.00193381583085372, 
    0.00193381583085372, 0.00193381583085372, 0.00193381583085372, 
    0.00193381583085372, 0.0019338158308535, 0.00193381583085372, 
    0.00193381583085372, 0.00193381583085372, 0.0019338158308535, 
    0.00193381583085395, 0.0019338158308535, 0.00193381583085372, 
    0.00193381583085395, 0.0019338158308535, 0.00193381583085372, 
    0.00193381583085372, 0.00193381583085372, 0.0019338158308535, 
    0.00193381583085372, 0.00193381583085372, 0.0019338158308535, 
    0.00193381583085395, 0.00193381583085372, 0.0019338158308535, 
    0.00193381583085395, 0.0019338158308535, 0.00193381583085372, 
    0.00193381583085372, 0.00193381583085372, 0.00193381583085372, 
    0.00193381583085372, 0.00193381583085372,
  0.0019464250686545, 0.0019464250686545, 0.0019464250686545, 
    0.00194642506865406, 0.0019464250686545, 0.00194642506865428, 
    0.00194642506865428, 0.0019464250686545, 0.00194642506865428, 
    0.00194642506865428, 0.00194642506865428, 0.0019464250686545, 
    0.00194642506865406, 0.00194642506865428, 0.0019464250686545, 
    0.00194642506865406, 0.0019464250686545, 0.0019464250686545, 
    0.00194642506865428, 0.00194642506865428, 0.00194642506865428, 
    0.0019464250686545, 0.00194642506865428, 0.00194642506865428, 
    0.00194642506865428, 0.00194642506865428, 0.00194642506865428, 
    0.00194642506865428, 0.00194642506865428, 0.00194642506865428, 
    0.00194642506865428, 0.00194642506865428, 0.00194642506865428, 
    0.0019464250686545, 0.00194642506865428, 0.00194642506865428, 
    0.0019464250686545, 0.00194642506865428, 0.00194642506865428, 
    0.00194642506865428, 0.00194642506865428, 0.00194642506865428, 
    0.00194642506865428, 0.00194642506865428, 0.00194642506865428, 
    0.0019464250686545, 0.00194642506865428, 0.00194642506865428, 
    0.0019464250686545, 0.00194642506865428, 0.00194642506865428, 
    0.00194642506865428, 0.00194642506865428, 0.00194642506865428, 
    0.00194642506865428, 0.00194642506865428,
  0.00195896842680554, 0.00195896842680554, 0.00195896842680554, 
    0.0019589684268051, 0.00195896842680554, 0.00195896842680532, 
    0.00195896842680532, 0.00195896842680554, 0.00195896842680532, 
    0.00195896842680532, 0.00195896842680532, 0.00195896842680554, 
    0.0019589684268051, 0.00195896842680532, 0.00195896842680554, 
    0.0019589684268051, 0.00195896842680554, 0.00195896842680554, 
    0.00195896842680532, 0.00195896842680532, 0.00195896842680532, 
    0.00195896842680554, 0.00195896842680532, 0.00195896842680532, 
    0.00195896842680532, 0.00195896842680532, 0.00195896842680532, 
    0.00195896842680532, 0.00195896842680532, 0.00195896842680532, 
    0.00195896842680532, 0.00195896842680532, 0.00195896842680532, 
    0.00195896842680554, 0.00195896842680532, 0.00195896842680532, 
    0.00195896842680554, 0.00195896842680532, 0.00195896842680532, 
    0.00195896842680532, 0.00195896842680532, 0.00195896842680532, 
    0.00195896842680532, 0.00195896842680532, 0.00195896842680532, 
    0.00195896842680554, 0.00195896842680532, 0.00195896842680532, 
    0.00195896842680554, 0.00195896842680532, 0.00195896842680532, 
    0.00195896842680532, 0.00195896842680532, 0.00195896842680532, 
    0.00195896842680532, 0.00195896842680532,
  0.00197144548063166, 0.00197144548063166, 0.00197144548063166, 
    0.00197144548063122, 0.00197144548063166, 0.00197144548063144, 
    0.00197144548063144, 0.00197144548063166, 0.00197144548063144, 
    0.00197144548063144, 0.00197144548063144, 0.00197144548063166, 
    0.00197144548063122, 0.00197144548063144, 0.00197144548063166, 
    0.00197144548063122, 0.00197144548063166, 0.00197144548063166, 
    0.00197144548063144, 0.00197144548063144, 0.00197144548063144, 
    0.00197144548063166, 0.00197144548063144, 0.00197144548063144, 
    0.00197144548063144, 0.00197144548063144, 0.00197144548063144, 
    0.00197144548063144, 0.00197144548063144, 0.00197144548063144, 
    0.00197144548063144, 0.00197144548063144, 0.00197144548063144, 
    0.00197144548063166, 0.00197144548063144, 0.00197144548063144, 
    0.00197144548063166, 0.00197144548063144, 0.00197144548063144, 
    0.00197144548063144, 0.00197144548063144, 0.00197144548063144, 
    0.00197144548063144, 0.00197144548063144, 0.00197144548063144, 
    0.00197144548063166, 0.00197144548063144, 0.00197144548063144, 
    0.00197144548063166, 0.00197144548063144, 0.00197144548063144, 
    0.00197144548063144, 0.00197144548063144, 0.00197144548063144, 
    0.00197144548063144, 0.00197144548063144,
  0.00198385580797655, 0.00198385580797655, 0.00198385580797655, 
    0.00198385580797611, 0.00198385580797655, 0.00198385580797655, 
    0.00198385580797633, 0.00198385580797655, 0.00198385580797655, 
    0.00198385580797633, 0.00198385580797655, 0.00198385580797655, 
    0.00198385580797611, 0.00198385580797655, 0.00198385580797655, 
    0.00198385580797611, 0.00198385580797655, 0.00198385580797655, 
    0.00198385580797633, 0.00198385580797655, 0.00198385580797633, 
    0.00198385580797655, 0.00198385580797633, 0.00198385580797655, 
    0.00198385580797655, 0.00198385580797655, 0.00198385580797655, 
    0.00198385580797655, 0.00198385580797633, 0.00198385580797655, 
    0.00198385580797655, 0.00198385580797655, 0.00198385580797633, 
    0.00198385580797655, 0.00198385580797633, 0.00198385580797655, 
    0.00198385580797655, 0.00198385580797633, 0.00198385580797655, 
    0.00198385580797655, 0.00198385580797655, 0.00198385580797633, 
    0.00198385580797655, 0.00198385580797655, 0.00198385580797633, 
    0.00198385580797655, 0.00198385580797655, 0.00198385580797633, 
    0.00198385580797655, 0.00198385580797633, 0.00198385580797655, 
    0.00198385580797655, 0.00198385580797655, 0.00198385580797655, 
    0.00198385580797655, 0.00198385580797655,
  0.00199619898874537, 0.00199619898874537, 0.00199619898874537, 
    0.00199619898874492, 0.00199619898874537, 0.00199619898874515, 
    0.00199619898874492, 0.00199619898874537, 0.00199619898874515, 
    0.00199619898874492, 0.00199619898874515, 0.00199619898874537, 
    0.00199619898874492, 0.00199619898874515, 0.00199619898874537, 
    0.00199619898874492, 0.00199619898874537, 0.00199619898874537, 
    0.00199619898874492, 0.00199619898874515, 0.00199619898874492, 
    0.00199619898874537, 0.00199619898874492, 0.00199619898874515, 
    0.00199619898874515, 0.00199619898874515, 0.00199619898874515, 
    0.00199619898874515, 0.00199619898874492, 0.00199619898874515, 
    0.00199619898874515, 0.00199619898874515, 0.00199619898874492, 
    0.00199619898874537, 0.00199619898874492, 0.00199619898874515, 
    0.00199619898874537, 0.00199619898874492, 0.00199619898874515, 
    0.00199619898874515, 0.00199619898874515, 0.00199619898874492, 
    0.00199619898874515, 0.00199619898874515, 0.00199619898874492, 
    0.00199619898874537, 0.00199619898874515, 0.00199619898874492, 
    0.00199619898874537, 0.00199619898874492, 0.00199619898874515, 
    0.00199619898874515, 0.00199619898874515, 0.00199619898874515, 
    0.00199619898874515, 0.00199619898874515,
  0.00200847460511366, 0.00200847460511366, 0.00200847460511366, 
    0.00200847460511322, 0.00200847460511366, 0.00200847460511366, 
    0.00200847460511344, 0.00200847460511366, 0.00200847460511366, 
    0.00200847460511344, 0.00200847460511366, 0.00200847460511366, 
    0.00200847460511322, 0.00200847460511366, 0.00200847460511366, 
    0.00200847460511322, 0.00200847460511366, 0.00200847460511366, 
    0.00200847460511344, 0.00200847460511366, 0.00200847460511344, 
    0.00200847460511366, 0.00200847460511344, 0.00200847460511366, 
    0.00200847460511366, 0.00200847460511366, 0.00200847460511366, 
    0.00200847460511366, 0.00200847460511344, 0.00200847460511366, 
    0.00200847460511366, 0.00200847460511366, 0.00200847460511344, 
    0.00200847460511366, 0.00200847460511344, 0.00200847460511366, 
    0.00200847460511366, 0.00200847460511344, 0.00200847460511366, 
    0.00200847460511366, 0.00200847460511366, 0.00200847460511344, 
    0.00200847460511366, 0.00200847460511366, 0.00200847460511344, 
    0.00200847460511366, 0.00200847460511366, 0.00200847460511344, 
    0.00200847460511366, 0.00200847460511344, 0.00200847460511366, 
    0.00200847460511366, 0.00200847460511366, 0.00200847460511366, 
    0.00200847460511366, 0.00200847460511366,
  0.0020206822416815, 0.0020206822416815, 0.0020206822416815, 
    0.00202068224168106, 0.0020206822416815, 0.0020206822416815, 
    0.00202068224168128, 0.0020206822416815, 0.0020206822416815, 
    0.00202068224168128, 0.0020206822416815, 0.0020206822416815, 
    0.00202068224168106, 0.0020206822416815, 0.0020206822416815, 
    0.00202068224168106, 0.0020206822416815, 0.0020206822416815, 
    0.00202068224168128, 0.0020206822416815, 0.00202068224168128, 
    0.0020206822416815, 0.00202068224168128, 0.0020206822416815, 
    0.0020206822416815, 0.0020206822416815, 0.0020206822416815, 
    0.0020206822416815, 0.00202068224168128, 0.0020206822416815, 
    0.0020206822416815, 0.0020206822416815, 0.00202068224168128, 
    0.0020206822416815, 0.00202068224168128, 0.0020206822416815, 
    0.0020206822416815, 0.00202068224168128, 0.0020206822416815, 
    0.0020206822416815, 0.0020206822416815, 0.00202068224168128, 
    0.0020206822416815, 0.0020206822416815, 0.00202068224168128, 
    0.0020206822416815, 0.0020206822416815, 0.00202068224168128, 
    0.0020206822416815, 0.00202068224168128, 0.0020206822416815, 
    0.0020206822416815, 0.0020206822416815, 0.0020206822416815, 
    0.0020206822416815, 0.0020206822416815,
  0.00203282148530071, 0.00203282148530071, 0.00203282148530071, 
    0.00203282148530026, 0.00203282148530071, 0.00203282148530048, 
    0.00203282148530026, 0.00203282148530071, 0.00203282148530048, 
    0.00203282148530026, 0.00203282148530048, 0.00203282148530071, 
    0.00203282148530026, 0.00203282148530048, 0.00203282148530071, 
    0.00203282148530026, 0.00203282148530071, 0.00203282148530071, 
    0.00203282148530026, 0.00203282148530048, 0.00203282148530026, 
    0.00203282148530071, 0.00203282148530026, 0.00203282148530048, 
    0.00203282148530048, 0.00203282148530048, 0.00203282148530048, 
    0.00203282148530048, 0.00203282148530026, 0.00203282148530048, 
    0.00203282148530048, 0.00203282148530048, 0.00203282148530026, 
    0.00203282148530071, 0.00203282148530026, 0.00203282148530048, 
    0.00203282148530071, 0.00203282148530026, 0.00203282148530048, 
    0.00203282148530048, 0.00203282148530048, 0.00203282148530026, 
    0.00203282148530048, 0.00203282148530048, 0.00203282148530026, 
    0.00203282148530071, 0.00203282148530048, 0.00203282148530026, 
    0.00203282148530071, 0.00203282148530026, 0.00203282148530048, 
    0.00203282148530048, 0.00203282148530048, 0.00203282148530048, 
    0.00203282148530048, 0.00203282148530048,
  0.00204489192497914, 0.00204489192497914, 0.00204489192497914, 
    0.0020448919249787, 0.00204489192497914, 0.00204489192497914, 
    0.00204489192497892, 0.00204489192497914, 0.00204489192497914, 
    0.00204489192497892, 0.00204489192497914, 0.00204489192497914, 
    0.0020448919249787, 0.00204489192497914, 0.00204489192497914, 
    0.0020448919249787, 0.00204489192497914, 0.00204489192497914, 
    0.00204489192497892, 0.00204489192497914, 0.00204489192497892, 
    0.00204489192497914, 0.00204489192497892, 0.00204489192497914, 
    0.00204489192497914, 0.00204489192497914, 0.00204489192497914, 
    0.00204489192497914, 0.00204489192497892, 0.00204489192497914, 
    0.00204489192497914, 0.00204489192497914, 0.00204489192497892, 
    0.00204489192497914, 0.00204489192497892, 0.00204489192497914, 
    0.00204489192497914, 0.00204489192497892, 0.00204489192497914, 
    0.00204489192497914, 0.00204489192497914, 0.00204489192497892, 
    0.00204489192497914, 0.00204489192497914, 0.00204489192497892, 
    0.00204489192497914, 0.00204489192497914, 0.00204489192497892, 
    0.00204489192497914, 0.00204489192497892, 0.00204489192497914, 
    0.00204489192497914, 0.00204489192497914, 0.00204489192497914, 
    0.00204489192497914, 0.00204489192497914,
  0.00205689315234014, 0.00205689315234014, 0.00205689315234014, 
    0.0020568931523397, 0.00205689315234014, 0.00205689315233992, 
    0.0020568931523397, 0.00205689315234014, 0.00205689315233992, 
    0.0020568931523397, 0.00205689315233992, 0.00205689315234014, 
    0.0020568931523397, 0.00205689315233992, 0.00205689315234014, 
    0.0020568931523397, 0.00205689315234014, 0.00205689315234014, 
    0.0020568931523397, 0.00205689315233992, 0.0020568931523397, 
    0.00205689315234014, 0.0020568931523397, 0.00205689315233992, 
    0.00205689315233992, 0.00205689315233992, 0.00205689315233992, 
    0.00205689315233992, 0.0020568931523397, 0.00205689315233992, 
    0.00205689315233992, 0.00205689315233992, 0.0020568931523397, 
    0.00205689315234014, 0.0020568931523397, 0.00205689315233992, 
    0.00205689315234014, 0.0020568931523397, 0.00205689315233992, 
    0.00205689315233992, 0.00205689315233992, 0.0020568931523397, 
    0.00205689315233992, 0.00205689315233992, 0.0020568931523397, 
    0.00205689315234014, 0.00205689315233992, 0.0020568931523397, 
    0.00205689315234014, 0.0020568931523397, 0.00205689315233992, 
    0.00205689315233992, 0.00205689315233992, 0.00205689315233992, 
    0.00205689315233992, 0.00205689315233992,
  0.00206882476106718, 0.00206882476106718, 0.00206882476106718, 
    0.00206882476106673, 0.00206882476106718, 0.00206882476106696, 
    0.00206882476106696, 0.00206882476106718, 0.00206882476106696, 
    0.00206882476106696, 0.00206882476106696, 0.00206882476106718, 
    0.00206882476106673, 0.00206882476106696, 0.00206882476106718, 
    0.00206882476106673, 0.00206882476106718, 0.00206882476106718, 
    0.00206882476106696, 0.00206882476106696, 0.00206882476106696, 
    0.00206882476106718, 0.00206882476106696, 0.00206882476106696, 
    0.00206882476106696, 0.00206882476106696, 0.00206882476106696, 
    0.00206882476106696, 0.00206882476106696, 0.00206882476106696, 
    0.00206882476106696, 0.00206882476106696, 0.00206882476106696, 
    0.00206882476106718, 0.00206882476106696, 0.00206882476106696, 
    0.00206882476106718, 0.00206882476106696, 0.00206882476106696, 
    0.00206882476106696, 0.00206882476106696, 0.00206882476106696, 
    0.00206882476106696, 0.00206882476106696, 0.00206882476106696, 
    0.00206882476106718, 0.00206882476106696, 0.00206882476106696, 
    0.00206882476106718, 0.00206882476106696, 0.00206882476106696, 
    0.00206882476106696, 0.00206882476106696, 0.00206882476106696, 
    0.00206882476106696, 0.00206882476106696,
  0.00208068634738279, 0.00208068634738279, 0.00208068634738279, 
    0.00208068634738234, 0.00208068634738279, 0.00208068634738279, 
    0.00208068634738257, 0.00208068634738279, 0.00208068634738279, 
    0.00208068634738257, 0.00208068634738279, 0.00208068634738279, 
    0.00208068634738234, 0.00208068634738279, 0.00208068634738279, 
    0.00208068634738234, 0.00208068634738279, 0.00208068634738279, 
    0.00208068634738257, 0.00208068634738279, 0.00208068634738257, 
    0.00208068634738279, 0.00208068634738257, 0.00208068634738279, 
    0.00208068634738279, 0.00208068634738279, 0.00208068634738279, 
    0.00208068634738279, 0.00208068634738257, 0.00208068634738279, 
    0.00208068634738279, 0.00208068634738279, 0.00208068634738257, 
    0.00208068634738279, 0.00208068634738257, 0.00208068634738279, 
    0.00208068634738279, 0.00208068634738257, 0.00208068634738279, 
    0.00208068634738279, 0.00208068634738279, 0.00208068634738257, 
    0.00208068634738279, 0.00208068634738279, 0.00208068634738257, 
    0.00208068634738279, 0.00208068634738279, 0.00208068634738257, 
    0.00208068634738279, 0.00208068634738257, 0.00208068634738279, 
    0.00208068634738279, 0.00208068634738279, 0.00208068634738279, 
    0.00208068634738279, 0.00208068634738279,
  0.00209247750985675, 0.00209247750985675, 0.00209247750985675, 
    0.00209247750985608, 0.00209247750985675, 0.00209247750985653, 
    0.00209247750985631, 0.00209247750985675, 0.00209247750985653, 
    0.00209247750985631, 0.00209247750985653, 0.00209247750985675, 
    0.00209247750985608, 0.00209247750985653, 0.00209247750985675, 
    0.00209247750985608, 0.00209247750985675, 0.00209247750985675, 
    0.00209247750985631, 0.00209247750985653, 0.00209247750985631, 
    0.00209247750985675, 0.00209247750985631, 0.00209247750985653, 
    0.00209247750985653, 0.00209247750985653, 0.00209247750985653, 
    0.00209247750985653, 0.00209247750985631, 0.00209247750985653, 
    0.00209247750985653, 0.00209247750985653, 0.00209247750985631, 
    0.00209247750985675, 0.00209247750985631, 0.00209247750985653, 
    0.00209247750985675, 0.00209247750985631, 0.00209247750985653, 
    0.00209247750985653, 0.00209247750985653, 0.00209247750985631, 
    0.00209247750985653, 0.00209247750985653, 0.00209247750985631, 
    0.00209247750985675, 0.00209247750985653, 0.00209247750985631, 
    0.00209247750985675, 0.00209247750985631, 0.00209247750985653, 
    0.00209247750985653, 0.00209247750985653, 0.00209247750985653, 
    0.00209247750985653, 0.00209247750985653,
  0.00210419784931015, 0.00210419784931015, 0.00210419784931015, 
    0.00210419784930971, 0.00210419784931015, 0.00210419784930993, 
    0.00210419784930993, 0.00210419784931015, 0.00210419784930993, 
    0.00210419784930993, 0.00210419784930993, 0.00210419784931015, 
    0.00210419784930971, 0.00210419784930993, 0.00210419784931015, 
    0.00210419784930971, 0.00210419784931015, 0.00210419784931015, 
    0.00210419784930993, 0.00210419784930993, 0.00210419784930993, 
    0.00210419784931015, 0.00210419784930993, 0.00210419784930993, 
    0.00210419784930993, 0.00210419784930993, 0.00210419784930993, 
    0.00210419784930993, 0.00210419784930993, 0.00210419784930993, 
    0.00210419784930993, 0.00210419784930993, 0.00210419784930993, 
    0.00210419784931015, 0.00210419784930993, 0.00210419784930993, 
    0.00210419784931015, 0.00210419784930993, 0.00210419784930993, 
    0.00210419784930993, 0.00210419784930993, 0.00210419784930993, 
    0.00210419784930993, 0.00210419784930993, 0.00210419784930993, 
    0.00210419784931015, 0.00210419784930993, 0.00210419784930993, 
    0.00210419784931015, 0.00210419784930993, 0.00210419784930993, 
    0.00210419784930993, 0.00210419784930993, 0.00210419784930993, 
    0.00210419784930993, 0.00210419784930993,
  0.00211584696916045, 0.00211584696916045, 0.00211584696916045, 
    0.00211584696915978, 0.00211584696916045, 0.00211584696916023, 
    0.00211584696916001, 0.00211584696916045, 0.00211584696916023, 
    0.00211584696916001, 0.00211584696916023, 0.00211584696916045, 
    0.00211584696915978, 0.00211584696916023, 0.00211584696916045, 
    0.00211584696915978, 0.00211584696916045, 0.00211584696916045, 
    0.00211584696916001, 0.00211584696916023, 0.00211584696916001, 
    0.00211584696916045, 0.00211584696916001, 0.00211584696916023, 
    0.00211584696916023, 0.00211584696916023, 0.00211584696916023, 
    0.00211584696916023, 0.00211584696916001, 0.00211584696916023, 
    0.00211584696916023, 0.00211584696916023, 0.00211584696916001, 
    0.00211584696916045, 0.00211584696916001, 0.00211584696916023, 
    0.00211584696916045, 0.00211584696916001, 0.00211584696916023, 
    0.00211584696916023, 0.00211584696916023, 0.00211584696916001, 
    0.00211584696916023, 0.00211584696916023, 0.00211584696916001, 
    0.00211584696916045, 0.00211584696916023, 0.00211584696916001, 
    0.00211584696916045, 0.00211584696916001, 0.00211584696916023, 
    0.00211584696916023, 0.00211584696916023, 0.00211584696916023, 
    0.00211584696916023, 0.00211584696916023,
  0.0021274244751337, 0.0021274244751337, 0.0021274244751337, 
    0.00212742447513303, 0.0021274244751337, 0.00212742447513348, 
    0.00212742447513325, 0.0021274244751337, 0.00212742447513348, 
    0.00212742447513325, 0.00212742447513348, 0.0021274244751337, 
    0.00212742447513303, 0.00212742447513348, 0.0021274244751337, 
    0.00212742447513303, 0.0021274244751337, 0.0021274244751337, 
    0.00212742447513325, 0.00212742447513348, 0.00212742447513325, 
    0.0021274244751337, 0.00212742447513325, 0.00212742447513348, 
    0.00212742447513348, 0.00212742447513348, 0.00212742447513348, 
    0.00212742447513348, 0.00212742447513325, 0.00212742447513348, 
    0.00212742447513348, 0.00212742447513348, 0.00212742447513325, 
    0.0021274244751337, 0.00212742447513325, 0.00212742447513348, 
    0.0021274244751337, 0.00212742447513325, 0.00212742447513348, 
    0.00212742447513348, 0.00212742447513348, 0.00212742447513325, 
    0.00212742447513348, 0.00212742447513348, 0.00212742447513325, 
    0.0021274244751337, 0.00212742447513348, 0.00212742447513325, 
    0.0021274244751337, 0.00212742447513325, 0.00212742447513348, 
    0.00212742447513348, 0.00212742447513348, 0.00212742447513348, 
    0.00212742447513348, 0.00212742447513348,
  0.00213892997530341, 0.00213892997530341, 0.00213892997530341, 
    0.00213892997530296, 0.00213892997530341, 0.00213892997530318, 
    0.00213892997530318, 0.00213892997530341, 0.00213892997530318, 
    0.00213892997530318, 0.00213892997530318, 0.00213892997530341, 
    0.00213892997530296, 0.00213892997530318, 0.00213892997530341, 
    0.00213892997530296, 0.00213892997530341, 0.00213892997530341, 
    0.00213892997530318, 0.00213892997530318, 0.00213892997530318, 
    0.00213892997530341, 0.00213892997530318, 0.00213892997530318, 
    0.00213892997530318, 0.00213892997530318, 0.00213892997530318, 
    0.00213892997530318, 0.00213892997530318, 0.00213892997530318, 
    0.00213892997530318, 0.00213892997530318, 0.00213892997530318, 
    0.00213892997530341, 0.00213892997530318, 0.00213892997530318, 
    0.00213892997530341, 0.00213892997530318, 0.00213892997530318, 
    0.00213892997530318, 0.00213892997530318, 0.00213892997530318, 
    0.00213892997530318, 0.00213892997530318, 0.00213892997530318, 
    0.00213892997530341, 0.00213892997530318, 0.00213892997530318, 
    0.00213892997530341, 0.00213892997530318, 0.00213892997530318, 
    0.00213892997530318, 0.00213892997530318, 0.00213892997530318, 
    0.00213892997530318, 0.00213892997530318,
  0.00215036308026262, 0.00215036308026262, 0.00215036308026262, 
    0.00215036308026217, 0.00215036308026262, 0.00215036308026262, 
    0.0021503630802624, 0.00215036308026262, 0.00215036308026262, 
    0.0021503630802624, 0.00215036308026262, 0.00215036308026262, 
    0.00215036308026217, 0.00215036308026262, 0.00215036308026262, 
    0.00215036308026217, 0.00215036308026262, 0.00215036308026262, 
    0.0021503630802624, 0.00215036308026262, 0.0021503630802624, 
    0.00215036308026262, 0.0021503630802624, 0.00215036308026262, 
    0.00215036308026262, 0.00215036308026262, 0.00215036308026262, 
    0.00215036308026262, 0.0021503630802624, 0.00215036308026262, 
    0.00215036308026262, 0.00215036308026262, 0.0021503630802624, 
    0.00215036308026262, 0.0021503630802624, 0.00215036308026262, 
    0.00215036308026262, 0.0021503630802624, 0.00215036308026262, 
    0.00215036308026262, 0.00215036308026262, 0.0021503630802624, 
    0.00215036308026262, 0.00215036308026262, 0.0021503630802624, 
    0.00215036308026262, 0.00215036308026262, 0.0021503630802624, 
    0.00215036308026262, 0.0021503630802624, 0.00215036308026262, 
    0.00215036308026262, 0.00215036308026262, 0.00215036308026262, 
    0.00215036308026262, 0.00215036308026262,
  0.00216172340308507, 0.00216172340308507, 0.00216172340308507, 
    0.00216172340308463, 0.00216172340308507, 0.00216172340308507, 
    0.00216172340308485, 0.00216172340308507, 0.00216172340308507, 
    0.00216172340308485, 0.00216172340308507, 0.00216172340308507, 
    0.00216172340308463, 0.00216172340308507, 0.00216172340308507, 
    0.00216172340308463, 0.00216172340308507, 0.00216172340308507, 
    0.00216172340308485, 0.00216172340308507, 0.00216172340308485, 
    0.00216172340308507, 0.00216172340308485, 0.00216172340308507, 
    0.00216172340308507, 0.00216172340308507, 0.00216172340308507, 
    0.00216172340308507, 0.00216172340308485, 0.00216172340308507, 
    0.00216172340308507, 0.00216172340308507, 0.00216172340308485, 
    0.00216172340308507, 0.00216172340308485, 0.00216172340308507, 
    0.00216172340308507, 0.00216172340308485, 0.00216172340308507, 
    0.00216172340308507, 0.00216172340308507, 0.00216172340308485, 
    0.00216172340308507, 0.00216172340308507, 0.00216172340308485, 
    0.00216172340308507, 0.00216172340308507, 0.00216172340308485, 
    0.00216172340308507, 0.00216172340308485, 0.00216172340308507, 
    0.00216172340308507, 0.00216172340308507, 0.00216172340308507, 
    0.00216172340308507, 0.00216172340308507 ;

 h =
  4544.23173916444, 4544.23173916444, 4544.79426389874, 4575.27187875418, 
    4627.88387506815, 4656.53924392246, 4631.08347903984, 4577.49706734492, 
    4552.47814461172, 4565.54221912462, 4586.18364719751, 4594.30447609547, 
    4574.39206650845, 4527.69684711849, 4495.83801948936, 4492.14709328146, 
    4467.64380074904, 4399.44136055673, 4327.49472148068, 4302.29688279779, 
    4320.35897876608, 4343.08814634039, 4358.20738541416, 4349.46475029001, 
    4289.75441283314, 4215.81804710384, 4185.22222271129, 4187.05275653615, 
    4189.38818301993, 4186.4490169725, 4175.66341773197, 4142.07739985843, 
    4075.70044918496, 3997.00312800151, 3944.25371901054, 3935.16549206096, 
    3951.2558047985, 3958.64548793587, 3943.45989706591, 3911.34708277734, 
    3862.1715666883, 3780.79737664238, 3678.11557646457, 3595.67176022016, 
    3501.49492621635, 3289.25979329267, 2896.58205795875, 2352.40586806033, 
    1772.09928153261, 1302.56677967285, 960.976870860982, 711.196259578647, 
    522.555355162128, 395.323088498131, 323.662451586529, 323.662451586529,
  4544.23173916444, 4544.23173916444, 4544.79426389874, 4575.27187875418, 
    4627.88387506815, 4656.53924392246, 4631.08347903984, 4577.49706734492, 
    4552.47814461172, 4565.54221912462, 4586.18364719751, 4594.30447609547, 
    4574.39206650845, 4527.69684711849, 4495.83801948936, 4492.14709328146, 
    4467.64380074904, 4399.44136055673, 4327.49472148068, 4302.29688279779, 
    4320.35897876608, 4343.08814634039, 4358.20738541416, 4349.46475029001, 
    4289.75441283314, 4215.81804710384, 4185.22222271129, 4187.05275653615, 
    4189.38818301993, 4186.4490169725, 4175.66341773197, 4142.07739985843, 
    4075.70044918496, 3997.00312800151, 3944.25371901054, 3935.16549206096, 
    3951.2558047985, 3958.64548793587, 3943.45989706591, 3911.34708277734, 
    3862.1715666883, 3780.79737664238, 3678.11557646457, 3595.67176022016, 
    3501.49492621635, 3289.25979329267, 2896.58205795875, 2352.40586806033, 
    1772.09928153261, 1302.56677967285, 960.976870860982, 711.196259578647, 
    522.555355162128, 395.323088498131, 323.662451586529, 323.662451586529,
  4581.20306850219, 4581.20306850219, 4581.05443610493, 4604.71946120312, 
    4646.54670934288, 4668.91718302023, 4642.97795096356, 4589.43046853591, 
    4562.31846514785, 4574.72143430655, 4598.07616632174, 4608.02692384179, 
    4587.5322195804, 4538.40625260849, 4498.02567931232, 4481.39651749719, 
    4448.80703087107, 4375.58943533342, 4294.01949303288, 4259.57370812034, 
    4280.9909609781, 4321.60253935474, 4357.0287159001, 4362.45089786222, 
    4311.35787693119, 4235.03204846224, 4189.87261251325, 4180.88537292758, 
    4180.97041782351, 4171.26804870582, 4146.13681235275, 4103.17921234677, 
    4046.36081877392, 3997.51670687154, 3978.95990758941, 3987.28481777666, 
    3999.29846022342, 3992.84820420204, 3963.40744799293, 3922.91335533047, 
    3878.55474333038, 3809.91438417508, 3702.02941591236, 3569.16450006744, 
    3373.21026382655, 3037.25614865833, 2559.08504641728, 2018.77701672062, 
    1508.65439707269, 1101.85843894156, 804.857064242746, 589.420523815565, 
    432.405454431678, 327.867105788503, 270.561290302579, 270.561290302579,
  4623.48833534044, 4623.48833534044, 4625.14308297671, 4638.80853527542, 
    4659.10093049708, 4664.876579305, 4636.29923315107, 4586.95346909775, 
    4559.88098009503, 4569.42963393316, 4592.64138892843, 4602.2119480859, 
    4578.84784914869, 4525.46862983985, 4475.64605906825, 4446.28825789006, 
    4409.6961336633, 4343.22514035204, 4268.75493274308, 4235.30178810939, 
    4256.20727567624, 4300.30483051158, 4341.06981543873, 4355.63545056018, 
    4320.84189534038, 4250.86150468709, 4189.93962693495, 4165.34013134978, 
    4163.87865036288, 4153.10365452407, 4121.53069379165, 4078.59485956991, 
    4038.31985303755, 4014.94129633134, 4013.96482627076, 4024.25773046066, 
    4026.96701675567, 4008.19534275141, 3968.61092777677, 3925.89555819141, 
    3889.10678853173, 3815.03229319934, 3652.32423194131, 3403.83859850201, 
    3048.63099772166, 2567.14694332822, 2033.12121939942, 1549.58325861452, 
    1149.410358201, 833.849817994801, 605.111913755601, 441.745291281403, 
    325.709794087748, 248.1380027957, 206.709043091792, 206.709043091792,
  4652.49641856838, 4652.49641856838, 4658.5461386928, 4662.93531597116, 
    4657.56341975582, 4640.42860451954, 4608.81642327584, 4571.97481931722, 
    4553.27888378034, 4559.03073255249, 4572.42395869682, 4572.33661759364, 
    4543.54532272951, 4489.45676601025, 4436.98801095366, 4401.77185089924, 
    4368.26614983131, 4322.03878856609, 4275.39563775351, 4255.77206939713, 
    4262.12073770524, 4270.89520606311, 4282.30934941684, 4297.82260378007, 
    4292.73002600475, 4249.92511298711, 4190.16411093688, 4155.80925090521, 
    4152.98117612948, 4148.64273940564, 4127.72165322691, 4101.17960632973, 
    4079.27211849663, 4060.8538276248, 4043.02344561869, 4027.71648229933, 
    4011.3481185846, 3983.18480503743, 3942.4715340666, 3901.76154164396, 
    3843.27458580368, 3685.46003687713, 3384.03405107853, 2990.73822956482, 
    2524.82272759487, 2005.92978069869, 1524.47099468206, 1144.66824908798, 
    846.049317940853, 610.484254076365, 442.456197990811, 323.9578135515, 
    239.886940147896, 183.087521960577, 152.880194252125, 152.880194252125,
  4659.13365936528, 4659.13365936528, 4675.43398069902, 4680.91745536224, 
    4657.66545888755, 4616.97801431754, 4579.62166961895, 4558.72163052341, 
    4554.67947359429, 4557.09097731079, 4553.84507677578, 4538.80438734522, 
    4508.69910722481, 4464.94124411728, 4419.78874711566, 4383.70059947938, 
    4352.531597622, 4315.71217121884, 4279.26319547345, 4264.80249812204, 
    4255.28910969561, 4220.77925907525, 4195.4200373486, 4215.46374165356, 
    4250.20252577742, 4251.82402282647, 4217.24173710575, 4186.55755234997, 
    4179.09714390133, 4176.52566650864, 4167.57510472287, 4157.86750123282, 
    4149.69353671237, 4132.89991472317, 4099.23465982375, 4054.36492033476, 
    4005.39597026007, 3953.25007095246, 3898.19546619301, 3821.44278441447, 
    3651.28505169201, 3311.16691219192, 2843.15538265381, 2362.62555133848, 
    1901.79030526253, 1465.89892099186, 1101.2866479768, 824.843822806377, 
    606.941334723719, 439.458989396382, 321.98879850632, 237.517464793998, 
    175.947038438146, 133.294688359389, 109.884937990091, 109.884937990091,
  4647.63529134803, 4647.63529134803, 4681.35148584362, 4700.55364451643, 
    4670.25970768922, 4607.61855649259, 4555.94730699649, 4536.8265102513, 
    4534.06571154281, 4527.24178105183, 4512.46491043904, 4493.88426033577, 
    4472.97585543645, 4447.24280229628, 4417.65876141512, 4390.84235993417, 
    4361.44573105093, 4301.58012341757, 4221.80030742787, 4191.51282768478, 
    4205.43577850412, 4193.82916410683, 4175.47459867039, 4202.14147844874, 
    4254.5132421351, 4285.25796122482, 4279.75955338952, 4259.27367699597, 
    4243.37739999847, 4232.64894977857, 4222.03372015607, 4211.33917252256, 
    4202.71346119134, 4190.03262671499, 4159.8625352122, 4102.99413920884, 
    4023.22836404036, 3932.55425236281, 3817.39975844179, 3612.52282600939, 
    3244.67739026829, 2734.00318511326, 2202.4614281815, 1747.57433009297, 
    1370.64878144944, 1048.11980560431, 787.951232380888, 587.759925055099, 
    429.667825556643, 313.14237482486, 231.94229675481, 171.8256163584, 
    126.946473875121, 94.7817862435477, 76.6650168625554, 76.6650168625554,
  4637.68969497669, 4637.68969497669, 4677.52803120923, 4692.73412900199, 
    4651.63967498131, 4588.19028259844, 4539.38068468956, 4510.11573477237, 
    4485.20928962466, 4459.68061337293, 4441.86485429655, 4433.39421457502, 
    4428.37308665449, 4421.83206469579, 4413.81411909414, 4407.98611895634, 
    4385.720936857, 4296.76810484593, 4163.08967015618, 4112.91227510697, 
    4170.96318975353, 4229.84071062217, 4255.28755154373, 4284.0517524371, 
    4322.53333122122, 4353.06468929402, 4361.85029231426, 4346.32875071427, 
    4319.39222334353, 4295.89375871934, 4272.12995894136, 4243.75772320817, 
    4220.99251678725, 4205.55370015074, 4180.28050399216, 4124.31391812456, 
    4029.62070005339, 3884.35765879391, 3627.65277117482, 3210.64769654756, 
    2666.51653057594, 2111.10050803224, 1636.34089602099, 1268.69199028966, 
    984.177998675156, 750.852294306836, 564.164699106238, 418.910247037904, 
    305.411496577657, 223.314271548412, 165.078777990805, 121.594604096877, 
    89.4592573763288, 66.1016868210483, 52.9644744472566, 52.9644744472566,
  4655.11660036142, 4655.11660036142, 4670.71017112609, 4640.2033972255, 
    4578.48435599508, 4555.73206062764, 4556.74475142744, 4528.66197025972, 
    4476.18024170199, 4431.52143962979, 4410.04166580416, 4406.15450279078, 
    4410.44737587045, 4419.12953263844, 4430.91037105882, 4442.69928865785, 
    4433.08713903214, 4359.98417850935, 4243.02753461369, 4191.54003458094, 
    4238.09651438767, 4302.58231814134, 4341.70731665728, 4368.51072827602, 
    4394.65775758866, 4421.48649514877, 4436.78299307274, 4420.79392651344, 
    4382.48971757325, 4347.61675794033, 4311.86659266128, 4267.78157218745, 
    4230.98244048305, 4203.45544599825, 4165.04368089032, 4095.17624398876, 
    3969.78509514393, 3721.36659555542, 3260.14276258651, 2660.39777091905, 
    2062.90760035477, 1572.30440162224, 1194.1278121366, 912.869622010108, 
    700.487004202836, 529.815402810136, 394.779509869509, 291.559155614352, 
    213.270111252041, 156.945280733921, 115.840190262992, 84.9505239394382, 
    62.5787481068954, 46.5053157320914, 37.6536739418347, 37.6536739418347,
  4722.17499895874, 4722.17499895874, 4711.72505206442, 4648.95236897551, 
    4589.95841975627, 4618.0849854606, 4665.92878030228, 4640.80534759011, 
    4573.59132227387, 4521.43144949398, 4494.05507496239, 4481.67958954755, 
    4478.87686643682, 4483.87423316343, 4493.58353364064, 4502.37703498201, 
    4499.81523266211, 4469.49207647492, 4413.90362619637, 4370.18203777397, 
    4358.29582978939, 4364.60689649414, 4379.85412032965, 4401.33306252238, 
    4426.24355326677, 4456.31380503157, 4479.31480120011, 4466.27910799341, 
    4421.69480901602, 4377.66805770294, 4336.62967611443, 4290.87854499481, 
    4249.24786919094, 4205.62996030446, 4129.87435582875, 3989.11344011646, 
    3749.44565231115, 3333.71377326732, 2707.39215845518, 2066.84332325927, 
    1533.4063370843, 1137.51387586013, 846.518820470319, 638.219763078127, 
    484.524898946922, 364.86949581633, 271.047325791245, 200.655914745441, 
    148.528742712036, 110.450993728711, 81.8217421229109, 60.0664150976212, 
    44.39150007444, 33.2283846328971, 27.1455914382647, 27.1455914382647,
  4839.197637147, 4839.197637147, 4833.20613518488, 4801.29393291243, 
    4785.08356147458, 4828.43249278775, 4863.26510967357, 4826.50193817306, 
    4762.91104655535, 4717.54642191982, 4686.17511130547, 4659.47704694789, 
    4634.40152762302, 4609.6371402811, 4590.58506774037, 4580.92455758778, 
    4574.48352202061, 4561.09053613555, 4531.59048054844, 4486.21162143848, 
    4439.53578308103, 4411.6966868979, 4410.32633597315, 4425.42114582258, 
    4445.71469973072, 4472.81246759508, 4498.17248118439, 4490.88682500138, 
    4445.49244773682, 4391.73051521803, 4348.32178645424, 4312.30383890512, 
    4271.68361300608, 4199.60689726054, 4039.12679141241, 3734.62510038382, 
    3291.31385317629, 2719.9800418162, 2076.29148568086, 1541.85372600583, 
    1130.96582493334, 822.176542462913, 596.974285161318, 442.382119308157, 
    331.452595963358, 249.050390407283, 185.464703758093, 138.466926437112, 
    104.011387437909, 78.0292501844521, 57.9614899389249, 42.6572007825565, 
    31.6454058609897, 23.8642346370132, 19.6604871852787, 19.6604871852787,
  4970.66419408737, 4970.66419408737, 4975.1587636182, 4982.44464757379, 
    5001.46833408445, 5030.23970843441, 5031.67364608269, 4992.92680239878, 
    4950.01298633855, 4916.42676778564, 4878.37902257174, 4834.80398179935, 
    4785.1867957837, 4728.50368077253, 4684.44128994845, 4666.14613894863, 
    4657.02876733997, 4638.94145816627, 4606.57786254995, 4561.77123589576, 
    4515.78390701885, 4486.13536541385, 4482.40245163123, 4496.40249647202, 
    4511.83478368329, 4526.04849492881, 4536.66631291294, 4522.4078719028, 
    4471.49269377475, 4405.39131088651, 4358.63802729304, 4333.11171033397, 
    4282.7337667682, 4139.38324482518, 3822.40794773347, 3297.5027851464, 
    2669.50595564834, 2052.3693377238, 1518.54720504216, 1127.47844918619, 
    828.075997332773, 594.219763613423, 421.987403819266, 307.341369845669, 
    227.067799567441, 169.488750048895, 126.464245699632, 95.4213355999122, 
    72.5806101206411, 54.8664994530235, 41.0314297053813, 30.5919710750778, 
    22.9923757922265, 17.5226730036082, 14.563966661654, 14.563966661654,
  5071.78968633837, 5071.78968633837, 5071.26768457787, 5078.95756132154, 
    5095.01037700239, 5107.42625091151, 5101.81445138946, 5081.97710501549, 
    5062.2563244778, 5032.71694318789, 4981.12649542033, 4922.90080226929, 
    4863.73787752757, 4799.57683135895, 4755.19735635622, 4744.04211661822, 
    4738.10320181809, 4719.04868696445, 4693.05417092001, 4663.40329183095, 
    4629.08626498677, 4598.70044222693, 4589.27088805911, 4601.03343159064, 
    4611.5360000834, 4607.68492192521, 4590.25656654651, 4553.51533591393, 
    4489.10246928203, 4411.32751206983, 4358.95876454559, 4328.21443151194, 
    4230.21445944968, 3955.78039263282, 3449.26310649583, 2755.11619613271, 
    2062.23614660648, 1501.13286080552, 1092.34349880951, 802.92410049247, 
    583.348716844789, 416.747059981793, 293.335353246967, 210.128482888655, 
    153.07836771147, 114.019792684054, 85.7988988319871, 65.5563766715868, 
    50.425537292467, 38.585086499834, 29.2690563082526, 22.250764294712, 
    17.1184670858479, 13.5187279623415, 11.6699447476716, 11.6699447476716,
  5123.6037491913, 5123.6037491913, 5114.98082386404, 5108.13546112219, 
    5107.43143459747, 5111.18561269296, 5113.94560251188, 5113.12016054178, 
    5103.95373683565, 5066.9858340723, 4999.25517723011, 4934.34500773128, 
    4884.41875751488, 4836.32584331279, 4805.14664663132, 4800.43567708298, 
    4796.05471248216, 4781.55536295418, 4769.2285492328, 4758.08073197528, 
    4736.05652541613, 4704.18424551834, 4682.35257080251, 4678.71262119273, 
    4674.20509152265, 4651.44770526897, 4609.10376095326, 4549.97174305126, 
    4472.46334737095, 4387.23521323761, 4323.09654640801, 4252.33889775095, 
    4044.2089370089, 3591.15778156123, 2934.65519077142, 2200.04145574465, 
    1568.09496054666, 1107.79128336172, 790.433250015548, 566.679079229781, 
    404.088477087324, 289.051310596887, 204.766845173323, 145.25349312548, 
    104.341975527756, 77.452359634942, 58.7784672768897, 45.5126595684195, 
    35.4903783850075, 27.5711601191515, 21.2350821651204, 16.4750942128851, 
    13.1996423965538, 11.2415790576685, 10.409478761505, 10.409478761505,
  5146.21917865266, 5146.21917865266, 5130.5142314379, 5111.45367395597, 
    5098.66022087426, 5099.38474696456, 5111.07325669628, 5122.69199744876, 
    5116.84029818707, 5071.59309554911, 4992.31657389434, 4922.65026436163, 
    4880.75897154188, 4849.25680825932, 4829.06982285497, 4824.11821546715, 
    4817.9895359485, 4807.30427498796, 4802.63851679231, 4800.47860369378, 
    4786.56429461038, 4756.71252659308, 4725.94913540466, 4705.57636932373, 
    4685.38639863575, 4649.34244850199, 4591.86038780602, 4517.82591387005, 
    4430.41260237482, 4336.33917868715, 4243.39811826083, 4086.08625529088, 
    3712.99188964242, 3082.46617377548, 2363.74045082882, 1700.02083959312, 
    1181.05917326087, 816.179419198417, 566.530139165009, 396.590716460574, 
    279.266599916123, 199.152883508988, 141.004320834194, 99.1288898794317, 
    70.6338321356094, 52.3837883832172, 40.1896894301902, 31.5995748748693, 
    25.0565945490081, 19.8574133551127, 15.7259832375162, 12.7859964397438, 
    11.0518349948811, 10.2800747563701, 10.0549181389887, 10.0549181389887,
  5162.88918317251, 5162.88918317251, 5137.45214422988, 5105.24156387863, 
    5083.20388945779, 5083.30833025408, 5101.94116544786, 5121.80875134795, 
    5120.09511952797, 5076.64032326632, 4997.86645060181, 4922.27382395131, 
    4871.77628850713, 4838.61491421393, 4819.90348010959, 4813.12007411494, 
    4805.75069982894, 4796.8403012922, 4794.03612663521, 4793.12417743015, 
    4781.43080943953, 4754.17220459011, 4723.49046337874, 4700.60039593835, 
    4677.97598602367, 4637.64098156932, 4570.63339318825, 4484.20027901151, 
    4383.61300523262, 4266.82282893864, 4114.89468148605, 3832.23348024767, 
    3294.11742427269, 2552.28931008592, 1849.48421544287, 1290.50808114165, 
    875.981588372673, 590.375783525561, 399.93392619858, 275.312605870548, 
    192.0469031884, 135.790008706509, 95.1757032073565, 66.2786027706133, 
    47.0576688794302, 35.0387804028303, 27.4226014978858, 22.0640038541592, 
    17.9562040835183, 14.7674378660872, 12.3789868551569, 10.8949028043696, 
    10.2223264155853, 10.0310955856371, 10.0029839377891, 10.0029839377891,
  5176.15916541235, 5176.15916541235, 5143.10547454374, 5099.77308200526, 
    5069.28913238004, 5065.84832059337, 5082.19850684781, 5098.68134721257, 
    5097.4598669813, 5065.19578460196, 5002.89617090307, 4930.95147344904, 
    4866.81387930512, 4817.38321972187, 4790.13190073947, 4781.45742887454, 
    4774.65741142494, 4767.27899810242, 4767.12367988064, 4768.96490446636, 
    4759.27665670042, 4733.92776066712, 4706.08030959187, 4687.70558738151, 
    4670.3384629767, 4631.41761354207, 4557.75671859636, 4456.37143674168, 
    4330.48344391035, 4163.63318405878, 3909.41132926724, 3467.10107177856, 
    2794.92068100642, 2026.83916048148, 1396.59999751819, 952.981885836902, 
    640.426000845145, 427.458484169389, 286.950241446432, 194.490278002865, 
    133.095631723312, 92.7924469017267, 64.475721731366, 44.8174204035951, 
    31.917084413833, 23.9754864126556, 19.3027225302532, 16.1003788893387, 
    13.6551729265486, 11.880080649277, 10.7359352604221, 10.1860477045788, 
    10.0224076750767, 10.0005131170989, 10.0001248664912, 10.0001248664912,
  5190.49000271153, 5190.49000271153, 5154.04106075283, 5101.66983316406, 
    5059.89609810296, 5045.48383366365, 5047.98922608201, 5049.38722622769, 
    5043.56773764359, 5025.41741844366, 4988.74703613935, 4934.83347015575, 
    4869.76620993803, 4807.15467022898, 4769.04117307282, 4757.46417456461, 
    4750.35513134789, 4743.95695448364, 4748.79768189956, 4756.51604654305, 
    4749.23608844465, 4722.91705974371, 4692.9392359658, 4673.6785440653, 
    4658.15870992903, 4622.16393645736, 4546.21137357283, 4428.11076013958, 
    4258.81831383792, 4000.66583884069, 3595.59658158535, 2981.33218784106, 
    2238.65068576824, 1543.1353088323, 1036.88391925549, 703.1331436664, 
    471.554918465099, 311.204526462214, 206.176962460931, 137.666248330503, 
    92.9415810233869, 64.2791451281258, 44.657596877656, 31.3521396018396, 
    22.6673925198056, 17.2855829930371, 14.3301018868186, 12.5535014641448, 
    11.3240329459503, 10.540456048312, 10.1447411855493, 10.0181871666948, 
    10, 10.000019806029, 10, 10,
  5199.52300481727, 5199.52300481727, 5163.56116209495, 5104.42198191636, 
    5049.46722240014, 5020.21690163272, 5006.65335648548, 4993.47638321382, 
    4983.42893008031, 4976.68810447706, 4962.96201999946, 4932.19502389073, 
    4879.78324856891, 4817.32271840589, 4774.50265584544, 4759.51480393845, 
    4749.45383624614, 4741.91772240244, 4749.52713660876, 4759.54742330249, 
    4749.60826114169, 4716.50008334076, 4678.02411533748, 4649.55459298059, 
    4625.78018022577, 4586.6159596643, 4510.50943325523, 4375.61146176183, 
    4135.48775609206, 3732.78859107865, 3161.29302314604, 2442.96767456191, 
    1733.64569739517, 1170.40157220408, 784.529739221816, 526.873764273077, 
    348.036801595876, 224.862756509542, 146.501563078794, 97.5599921298659, 
    66.3908246073321, 45.923354479416, 31.9393025583426, 22.698991026034, 
    16.8322121265398, 13.3322223580698, 11.5983456481262, 10.7812121114461, 
    10.3295129060452, 10.0954833024034, 10.0130965956596, 10, 10, 10, 10, 10,
  5172.77885125431, 5172.77885125431, 5146.95971893599, 5094.40749613154, 
    5036.40458001211, 4998.44596839565, 4976.11602561955, 4957.40656247379, 
    4947.28311547567, 4948.42766996238, 4949.89363590525, 4935.12888535496, 
    4894.03057068821, 4837.25897468012, 4794.75005608659, 4776.64399203855, 
    4763.45455115915, 4753.26239410765, 4756.71723175367, 4760.32042929743, 
    4741.7520204705, 4698.43287393831, 4649.11120138805, 4606.46587495899, 
    4562.79351333728, 4506.87073710926, 4422.31677705593, 4252.63889255741, 
    3895.44488278705, 3318.42290261877, 2633.86384511762, 1927.73197336663, 
    1328.05421995354, 890.66084410437, 589.23412466988, 384.645701229384, 
    248.658245023644, 158.66733086782, 102.942452550315, 68.9917714809962, 
    47.5674038312381, 32.9722252501071, 23.1307091696819, 16.8766766793574, 
    13.1580387477077, 11.2182888505073, 10.4255437263116, 10.155987335909, 
    10.0483464689256, 10.0075820262996, 10, 10, 10, 10, 10, 10,
  5111.14634555927, 5111.14634555927, 5106.26684250578, 5076.24515755, 
    5027.88540409757, 4987.39338863837, 4959.8107474887, 4940.52219438317, 
    4935.88819921325, 4947.27902198854, 4959.27361352726, 4949.05825277259, 
    4908.21957176732, 4853.43283294704, 4811.93323156036, 4791.46126498583, 
    4776.68428685794, 4763.34789424196, 4757.06393648163, 4748.41402147964, 
    4719.91122597929, 4668.12686599268, 4609.93657049945, 4554.56446228579, 
    4491.31270741627, 4411.97153202787, 4286.89088754598, 4014.06849099919, 
    3491.77267499983, 2789.38780962284, 2099.26261300059, 1487.40770222521, 
    1012.06684866134, 675.234849259198, 437.281121230085, 277.144768883424, 
    176.620238729104, 112.895663801299, 73.6599108387008, 49.3232344050752, 
    34.0271065418672, 23.7321368206641, 17.1527504144492, 13.2571637164537, 
    11.2016697522007, 10.3392195191824, 10.0756837160021, 10.0176576270894, 
    10.0031038825953, 10, 10, 10, 10, 10, 10, 10,
  5049.67138595013, 5049.67138595013, 5067.60542406193, 5063.89751079851, 
    5027.89791006065, 4983.53545629374, 4946.16700208192, 4923.72299755764, 
    4927.27133349758, 4951.89349447876, 4970.83309546978, 4956.52677131828, 
    4908.95898213139, 4854.58766776207, 4816.06694550385, 4794.74130811645, 
    4777.76876993947, 4760.60980808219, 4746.04567094837, 4727.83896141457, 
    4692.66132560991, 4636.28879526445, 4572.80886105318, 4511.3712003401, 
    4439.94461384366, 4329.14045770584, 4102.02256111553, 3649.22205601242, 
    2977.10289873391, 2255.68701552403, 1639.63288075758, 1137.09911118288, 
    761.641712868952, 498.854936350624, 315.368254462607, 197.198806933474, 
    126.258718727844, 82.0493841141155, 54.1239438784196, 36.1478147737722, 
    24.9594624553114, 17.7929160663186, 13.5674415653257, 11.3434302398691, 
    10.3733786617825, 10.0688613757661, 10.0074899455388, 10.0007299190201, 
    10, 10, 10, 10, 10, 10, 10, 10,
  4999.03556930938, 4999.03556930938, 5032.14086251412, 5048.28484582927, 
    5023.73569218206, 4978.24449098455, 4934.20304861928, 4908.61071313013, 
    4914.21514607438, 4940.79083122903, 4955.49329669772, 4931.13782760769, 
    4877.5424232746, 4828.98293610024, 4799.90633385549, 4780.44608713745, 
    4758.79576844505, 4737.09632226665, 4720.53233062683, 4700.08086456384, 
    4661.60660176137, 4602.69040983417, 4536.59002524094, 4471.45651343746, 
    4385.51001397637, 4210.34160397227, 3836.85759572864, 3216.67430934666, 
    2482.76587414399, 1812.79939294674, 1275.45036422527, 862.196272294677, 
    568.017740600984, 364.966557312296, 227.183842455158, 142.025400143616, 
    91.7879620845661, 60.5475569673054, 40.2515336648567, 26.9127192972148, 
    18.7547685381955, 13.964586045641, 11.5041184744298, 10.4367013737252, 
    10.0824245746129, 10.0075873411873, 10.0000621687022, 10, 10, 10, 10, 10, 
    10, 10, 10, 10,
  4960.7524801354, 4960.7524801354, 4994.57084579647, 5015.13350185835, 
    4997.99025716321, 4961.20480882811, 4925.8566001965, 4904.17746400561, 
    4902.9481481801, 4914.51958764567, 4913.98546717604, 4878.82474845302, 
    4824.26765752253, 4787.30532704934, 4772.03206176317, 4756.36639128958, 
    4729.57470277127, 4703.70081063454, 4688.20473373084, 4668.13877617017, 
    4626.96933598358, 4566.77400091861, 4499.44130537502, 4422.43737009986, 
    4290.39912446114, 4005.9601969358, 3486.12931013106, 2770.44371614665, 
    2051.15653682688, 1455.25519795456, 988.931305351921, 647.01502956072, 
    418.469072263054, 265.673439604375, 165.100743160168, 103.717307122545, 
    67.1538768619968, 44.4043874423909, 29.6576088912538, 20.1279260834423, 
    14.550396109898, 11.6859547903259, 10.4875128482173, 10.0957659248058, 
    10.0091708644146, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  4936.11912035897, 4936.11912035897, 4955.26915695677, 4960.5002022062, 
    4940.47641760816, 4916.1464097819, 4899.13078528273, 4885.16938159534, 
    4872.31578361781, 4865.37498957917, 4856.38731906834, 4822.71797097881, 
    4774.88373098531, 4748.59270822205, 4742.77001795915, 4730.41738926457, 
    4702.28637805698, 4674.10539449487, 4656.23361632123, 4632.98593479284, 
    4590.44720348649, 4533.11814210648, 4464.8656257746, 4362.05977661571, 
    4145.05030563499, 3710.00894683796, 3062.62802228546, 2318.68245452405, 
    1652.64714112384, 1139.06739681325, 754.005083347575, 480.980258901242, 
    305.566020361594, 191.768871485782, 118.573747201614, 74.5667938930242, 
    48.6774959836614, 32.4361987813435, 21.9168141024988, 15.4326363392078, 
    12.0063423297871, 10.5616434608605, 10.1079274632098, 10.0105873126637, 
    10.0000186791801, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  4887.2560406231, 4887.2560406231, 4886.85201609211, 4872.30271956829, 
    4845.41117668184, 4824.62265897612, 4813.35993617845, 4794.51654393397, 
    4760.33559603793, 4737.99048339646, 4741.34995380856, 4733.1603489658, 
    4702.60013007058, 4682.99510572864, 4679.02690860183, 4668.76873511235, 
    4644.41727821069, 4616.97270816365, 4594.8122023315, 4570.48653589544, 
    4535.84551212804, 4488.70785586877, 4416.70936019091, 4267.84999953574, 
    3928.05440160251, 3326.93224784872, 2602.3534324532, 1903.86770962884, 
    1318.65799925866, 878.724020912957, 567.370566240149, 356.420286038599, 
    224.384368864872, 140.388440220965, 86.6043816278155, 54.4864586683328, 
    36.0163989181802, 24.3523960305856, 16.9100698003414, 12.6953358416383, 
    10.7854145450795, 10.1538714924126, 10.016322574306, 10.0003510627118, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  4801.79829678032, 4801.79829678032, 4785.51058290586, 4760.27810161887, 
    4731.89302069667, 4704.12957670381, 4677.87149238163, 4637.64797039214, 
    4576.49610753292, 4543.10628480412, 4569.3320150847, 4597.44133554402, 
    4588.37273592226, 4570.95688228334, 4560.99418593481, 4547.75532645776, 
    4526.48514915931, 4501.56227442719, 4479.63115942357, 4464.47190245198, 
    4449.58271634254, 4415.25625921267, 4323.48379599903, 4093.9535581332, 
    3613.50625994771, 2891.45755600271, 2159.08970711296, 1544.57184634539, 
    1049.44547308013, 677.205531527741, 427.456807627975, 266.603101496854, 
    166.82201155934, 103.777496806263, 63.8559358322598, 40.4197198224133, 
    27.2239126381836, 18.9252187079723, 13.8459601936894, 11.2712268461851, 
    10.2901542475205, 10.0386291354675, 10.0019966973595, 10, 10, 10, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 10,
  4727.02285991146, 4727.02285991146, 4700.09419700867, 4669.80933413962, 
    4644.47163112952, 4613.04518300323, 4573.79041006497, 4521.68505216492, 
    4456.60375689636, 4426.78738177263, 4462.52369024686, 4505.23214129452, 
    4507.25153800635, 4486.0186349032, 4460.61721341729, 4433.37625374002, 
    4406.76041372769, 4382.44744662599, 4364.97764915308, 4362.49232863653, 
    4363.75760168316, 4326.65549809419, 4181.76299396045, 3837.92591288345, 
    3236.56927857968, 2478.44917265539, 1788.36256914993, 1244.14215094085, 
    824.585568336075, 518.778090443587, 322.10498843693, 199.737512531272, 
    124.077253582492, 76.9107029059059, 47.7679686550082, 30.8773733078067, 
    21.3615529599495, 15.4812555338298, 12.0779116061839, 10.5547135738679, 
    10.089561163426, 10.0063246827668, 10, 10, 10, 10, 10, 10, 10, 10, 10, 
    10, 10, 10, 10, 10,
  4616.05449450345, 4616.05449450345, 4601.03653710479, 4586.22050354798, 
    4574.76344804034, 4552.14367188861, 4519.22691564942, 4482.91941923461, 
    4447.09309708272, 4437.32644167042, 4468.88797284249, 4506.15544018085, 
    4513.58556342406, 4490.63935297604, 4451.72445858854, 4410.87017159726, 
    4376.48254456304, 4350.4134254351, 4335.19351656813, 4334.74092718997, 
    4330.1295967234, 4259.6738474441, 4023.73375463756, 3540.83502032133, 
    2835.44619178622, 2091.26124286338, 1471.35991090596, 993.821038231705, 
    642.080148015422, 399.589818434971, 246.931965177376, 152.587296351689, 
    94.4736174182958, 58.9581120114086, 37.3573099043511, 24.6803019014494, 
    17.4346756049812, 13.2064277319777, 11.0139187523135, 10.2001808377869, 
    10.0194124334715, 10.0004873000753, 10.0000163860455, 10, 10, 10, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 10,
  4388.45499413225, 4388.45499413225, 4412.69757254262, 4440.76188122343, 
    4454.32642340893, 4443.77695655915, 4424.46768529927, 4413.32664300872, 
    4409.57122898848, 4418.14821171211, 4447.08789598383, 4482.15217749897, 
    4495.30518449382, 4473.64010733752, 4437.19847774213, 4407.34070341218, 
    4380.62483518681, 4353.02347285656, 4330.59419387152, 4315.90856727412, 
    4285.70621593811, 4160.74555217737, 3814.28253741995, 3200.28907781825, 
    2431.78566404984, 1734.79638011504, 1200.67737018551, 799.319378354336, 
    509.612915096757, 315.219875520945, 193.706380174743, 119.702740590367, 
    74.2576921658226, 46.669016521812, 30.1132972141873, 20.2981912957317, 
    14.6621559315857, 11.6881776614399, 10.4203373138598, 10.0609453682501, 
    10.0045036418369, 10.0002203215302, 10, 10, 10, 10, 10, 10, 10, 10, 10, 
    10, 10, 10, 10, 10,
  4149.01571339975, 4149.01571339975, 4191.11783336121, 4234.2288353717, 
    4250.47238350395, 4237.75698057301, 4218.22134864859, 4208.4366488055, 
    4204.09362988181, 4205.28522337295, 4219.46656473449, 4237.1296682332, 
    4229.27669817631, 4189.14028064601, 4161.62444589177, 4169.09854893174, 
    4170.94919985913, 4141.98212772406, 4098.96990739928, 4060.95489038577, 
    4010.76472146909, 3852.84221657056, 3442.31324699904, 2784.20820042765, 
    2049.46686233756, 1435.57960024816, 981.344750877847, 647.782117235577, 
    409.57694668889, 251.592217689998, 154.366489527467, 96.4991507057383, 
    60.3806643385852, 37.9789708407552, 24.7196635371172, 17.0299890653755, 
    12.7863374491214, 10.826809723809, 10.162936549461, 10.0191001679898, 
    10.0011720352377, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  4011.82008535928, 4011.82008535928, 4022.77013449021, 4024.52799336808, 
    4010.78749904848, 3985.41248286322, 3953.91220086486, 3919.22495296686, 
    3881.89234099429, 3844.30611396935, 3810.79752490424, 3777.46961865125, 
    3724.85186977377, 3658.5723129732, 3638.39722250391, 3680.9218484277, 
    3712.13401644999, 3678.15102469608, 3601.67619379714, 3537.70342723393, 
    3494.63771680641, 3369.43022728182, 2998.76586075633, 2402.19150986505, 
    1760.48797606723, 1222.70201868364, 823.400597087819, 537.986253902339, 
    337.879047583519, 206.748290785476, 127.237959422347, 80.7134230333706, 
    51.1939192039835, 32.3088767537537, 21.1801595174696, 14.8887054020675, 
    11.6544994903164, 10.3885464101792, 10.0561648541273, 10.0039138060888, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3923.12609855637, 3923.12609855637, 3897.27893508507, 3857.74517083855, 
    3822.88815990133, 3796.59583501158, 3760.55006921451, 3702.87291545834, 
    3631.02544026278, 3546.51799708542, 3452.41398045105, 3368.12896878141, 
    3299.58195181178, 3247.90923595321, 3243.95261704729, 3292.21983622061, 
    3326.61324852029, 3279.24864302443, 3163.02321652507, 3070.35644726451, 
    3046.01107933634, 2983.92055337905, 2694.8276608548, 2175.56065571925, 
    1608.58668972091, 1114.74849759263, 742.356287198545, 480.891512511174, 
    302.19965160457, 185.384163831752, 113.77572585922, 72.3094678372059, 
    46.42866874255, 29.5464977727653, 19.4295727901744, 13.7534319267703, 
    11.0665614626471, 10.190052993248, 10.0181144689625, 10.000671067418, 
    10.0000219641831, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3830.14602593956, 3830.14602593956, 3796.77393253335, 3753.43012995293, 
    3722.95904793933, 3704.97085505299, 3667.14149475081, 3593.38049263348, 
    3502.37885758472, 3397.16478963598, 3278.20865563353, 3180.62448664423, 
    3131.50456221156, 3122.42693791535, 3139.40436342407, 3171.80441522109, 
    3185.25358566856, 3118.93934036762, 2971.38382772115, 2850.60827525239, 
    2827.24903922201, 2803.84146300579, 2573.32233960731, 2094.26522599658, 
    1558.12500290486, 1083.06340921438, 718.22429956445, 459.655875840931, 
    287.326002896674, 176.654020009561, 108.330064043346, 68.4542851635969, 
    44.1676615910654, 28.5025092075394, 18.8260300336639, 13.294449866969, 
    10.8350610039873, 10.1280246815522, 10.010377638874, 10.0003480749477, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3756.17000237666, 3756.17000237666, 3731.59775036371, 3697.89985381481, 
    3673.44729274386, 3659.06736079483, 3616.522612787, 3530.44847371164, 
    3436.42169729927, 3347.12230889334, 3253.16641624978, 3175.35734826599, 
    3142.18137237787, 3151.82462844282, 3176.83620189116, 3194.83473797697, 
    3185.66539703096, 3105.60199465358, 2951.16214430058, 2815.29884462757, 
    2765.79002043676, 2721.5564003064, 2484.97052859275, 2005.30229549282, 
    1483.8020090508, 1034.9483369041, 685.534354371935, 432.531750335323, 
    267.720081221938, 164.848639243923, 101.399602204598, 63.7789489994822, 
    41.1964088088524, 27.1192355027574, 18.2721508752003, 13.0352800675696, 
    10.7484588459055, 10.1163292253955, 10.0108887368136, 10.0005269121419, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3720.24622881651, 3720.24622881651, 3695.54889929353, 3655.3178991069, 
    3624.11154851884, 3615.2774174082, 3587.00269735964, 3514.62787944754, 
    3436.57113291195, 3372.37081772538, 3307.85480079123, 3247.79033189277, 
    3213.85813625765, 3214.52395771136, 3232.01116241345, 3240.22188594625, 
    3216.59664886538, 3134.97923687234, 2997.61521045526, 2862.94380882712, 
    2774.33067701416, 2667.35003963622, 2378.71191870917, 1884.97711330584, 
    1376.95492747365, 954.356378739467, 627.758077957933, 392.102709787848, 
    241.472409867714, 148.547981560455, 91.3425243066205, 57.5082062153008, 
    37.285122085822, 24.9647786970087, 17.2894918025721, 12.6383929758253, 
    10.6177444727306, 10.0842063575763, 10.0052652755136, 10, 10, 10, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3716.99767974781, 3716.99767974781, 3678.25832845059, 3619.3481973661, 
    3578.98294620222, 3580.66382591329, 3582.46677093211, 3546.74692074078, 
    3494.89193962983, 3442.79013746363, 3383.50459174402, 3324.26536892205, 
    3283.71319416693, 3270.7649196346, 3274.62306323157, 3272.03484565554, 
    3239.09967630765, 3159.91708456433, 3040.53870222754, 2914.42136531486, 
    2799.83284512515, 2629.85572292145, 2272.60277944449, 1759.53226880811, 
    1264.68362608744, 864.450358355574, 564.588416286183, 352.71030742076, 
    217.840121577415, 134.238343526031, 82.6648845486766, 52.2208072088846, 
    33.8973636624134, 22.8031994445339, 16.1051298486417, 12.1401899689354, 
    10.4797250943687, 10.0645052237544, 10.0052237701732, 10.0002766630273, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3736.28565796575, 3736.28565796575, 3683.85251007521, 3615.95814850175, 
    3576.4561970644, 3581.73833716013, 3595.63839706645, 3582.16942632036, 
    3546.37228134537, 3497.84373656117, 3438.04372236093, 3377.12961270603, 
    3330.73820049205, 3307.07070025587, 3299.09884507364, 3287.33571702546, 
    3247.77171976569, 3164.9535493562, 3046.99423822845, 2923.57069301325, 
    2798.1523242531, 2586.94181610343, 2178.71239155108, 1662.17362922171, 
    1187.79618214915, 803.992203700001, 522.539859712086, 327.775364220996, 
    202.705972496952, 124.106734267115, 76.1232537808751, 48.4713930723974, 
    31.8959471079217, 21.6209966503862, 15.3594947519482, 11.7901869316948, 
    10.3819289178249, 10.0480937502139, 10.0029210821302, 10, 10, 10, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3766.43139210862, 3766.43139210862, 3711.06324913093, 3647.06758155152, 
    3612.36560926698, 3610.32555351616, 3613.48694024747, 3597.28754875667, 
    3561.59773327584, 3514.83617485023, 3461.32958366229, 3403.86920943719, 
    3352.35273834959, 3319.09448395071, 3302.33672306021, 3284.63474608588, 
    3242.33810390076, 3159.85853279641, 3046.21335938782, 2931.27604315517, 
    2809.19845032487, 2576.97316288632, 2132.5644272541, 1613.04675549634, 
    1153.82176914793, 779.560088771833, 504.299154919435, 316.075452833303, 
    195.567909773856, 119.593407756097, 73.3284296905944, 46.8801858944773, 
    31.0865143622674, 21.0405844248915, 14.814413826028, 11.4585970066919, 
    10.2696036699213, 10.0277665914582, 10.0015117598835, 10.0000644610775, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3785.97291950549, 3785.97291950549, 3735.47128349476, 3677.72400805657, 
    3643.28818126647, 3631.10779813846, 3620.56070608258, 3593.7420938922, 
    3550.20151471266, 3501.57446042461, 3454.21813534855, 3403.29615594604, 
    3351.71756966819, 3312.05053561855, 3285.11726821828, 3256.89411721658, 
    3210.83734364855, 3138.32030975494, 3047.37269968776, 2957.42172230504, 
    2848.48203807726, 2605.29489710413, 2134.95632716296, 1607.2927402674, 
    1152.63687469323, 779.831588123358, 499.787673613171, 310.108315876548, 
    191.719631113694, 118.150306165818, 72.7527866488589, 46.319504692059, 
    30.6444410651756, 20.6318629126344, 14.486368689276, 11.3010873725727, 
    10.2267215032046, 10.0210294100446, 10.0008019045596, 10, 10, 10, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3779.09992050158, 3779.09992050158, 3733.31021054086, 3679.86662343366, 
    3644.63435538579, 3626.01537761518, 3608.18520875199, 3575.0867819061, 
    3522.37510243825, 3462.27413769126, 3408.30167413314, 3361.13412303453, 
    3316.9444779573, 3273.87790446115, 3228.74522142682, 3178.93079666831, 
    3125.16525359895, 3066.06640326213, 3004.88653409442, 2950.78708672352, 
    2869.83867834626, 2637.11394303528, 2162.20937799443, 1623.67061799859, 
    1164.25694904175, 790.624043431336, 505.030056301288, 310.513012869916, 
    190.248297208593, 117.49229935716, 72.8915574395726, 46.2716199110048, 
    30.4900634115824, 20.5213283760692, 14.5349065320772, 11.397090433298, 
    10.2733049609116, 10.0311343506842, 10.0016709838558, 10, 10, 10, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3770.37106395758, 3770.37106395758, 3727.66262426148, 3677.79487182195, 
    3641.82973694807, 3616.61817776818, 3593.8714076632, 3559.62947989686, 
    3496.21506893784, 3405.93796086025, 3315.24705610092, 3250.74421773149, 
    3207.06345318788, 3154.64134846657, 3083.4690277705, 3013.87613723076, 
    2969.4752968327, 2944.60187941578, 2924.74619928355, 2910.88413079755, 
    2864.04190116884, 2655.15334139847, 2186.00261124401, 1626.13337927985, 
    1155.21826990411, 788.021990387383, 508.847757219354, 315.307610754392, 
    191.852692729502, 117.55591976617, 73.1582144671892, 46.3645595194407, 
    30.4747314208694, 20.5937897053354, 14.7030713228801, 11.5157501208775, 
    10.3139902368163, 10.0395225961707, 10.0030038841453, 10.0001466653355, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3787.00453013841, 3787.00453013841, 3748.18155478593, 3701.74353082747, 
    3662.60429189536, 3627.60236257049, 3598.03407212345, 3559.8422170101, 
    3475.08027485218, 3331.75251145273, 3174.85727707907, 3069.22497822846, 
    3014.70174070946, 2953.66596259823, 2869.81141533781, 2804.87034301405, 
    2797.29527579928, 2828.80917568083, 2859.89167364941, 2880.73457821072, 
    2860.08164813801, 2677.31779950809, 2214.53284012439, 1620.66902439342, 
    1126.22091088626, 764.405815633645, 498.435624770413, 313.877451018635, 
    192.040428231099, 116.943125070791, 72.4457974204533, 45.8601525100039, 
    30.2627637243165, 20.6150265827902, 14.7619088353863, 11.534693347568, 
    10.3132324214944, 10.0375027418047, 10.0022000483977, 10, 10, 10, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3810.90452121907, 3810.90452121907, 3774.04564659813, 3728.77663965445, 
    3687.14784112389, 3646.33529705733, 3608.20328049974, 3551.12354545534, 
    3424.74582532088, 3219.52203722426, 3003.67622809467, 2867.81591998379, 
    2816.06137915023, 2776.80662871119, 2723.7470652982, 2693.3691659231, 
    2718.04750395417, 2777.98846288656, 2832.95102779353, 2868.50567497877, 
    2857.79125886445, 2691.70776270657, 2244.98255873436, 1647.72272806123, 
    1144.11751237036, 776.883691224685, 506.803288714702, 319.834764285614, 
    196.799145528879, 120.39241749602, 74.7232356686049, 47.2925849000243, 
    31.1673149998432, 21.2292384939373, 15.0484224300297, 11.6057301119406, 
    10.3130137126761, 10.033150608172, 10.0017039022688, 10.0000784029565, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3826.24917714508, 3826.24917714508, 3785.20530745337, 3734.48102224701, 
    3690.21602185763, 3648.20898339941, 3596.96854340373, 3503.36913372661, 
    3325.41562825746, 3078.19039210233, 2844.60241076616, 2708.46733948161, 
    2675.11539980514, 2684.3773088691, 2696.39135222079, 2712.79359651867, 
    2745.47165199874, 2789.85047035293, 2832.26740029155, 2862.61839969347, 
    2848.78836997392, 2687.39212418284, 2262.7314139474, 1695.0171320809, 
    1202.51645685028, 823.584910375753, 538.120248992009, 341.23550597022, 
    212.448270831842, 130.67927067047, 81.0151634184398, 51.0240930345213, 
    33.4061189932241, 22.722988316686, 15.9439132355225, 12.0313295356759, 
    10.4500524224869, 10.0588453255851, 10.0036634033917, 10, 10, 10, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3836.67970979765, 3836.67970979765, 3788.82657344893, 3726.89409667394, 
    3671.66182768311, 3618.13599571289, 3542.76337736069, 3409.14858692464, 
    3196.47440012559, 2945.08151768468, 2730.53022747171, 2603.16004228534, 
    2575.30557134341, 2624.1802720423, 2697.54571719374, 2752.69194474371, 
    2785.69800274958, 2811.73165315974, 2840.31268238535, 2863.42456006567, 
    2844.82887796461, 2686.41494420883, 2279.6090590975, 1736.08155520326, 
    1253.10555290749, 866.173066508666, 569.752058839368, 364.088643152935, 
    229.115634933454, 141.390835052224, 87.6105056749991, 55.0660960151001, 
    35.9739055743272, 24.5105924984576, 17.1136321767876, 12.645879402195, 
    10.6633023964596, 10.1042280834232, 10.0097735490412, 10.000499057799, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3830.06558168122, 3830.06558168122, 3783.0639687308, 3713.90435324358, 
    3636.77288851886, 3550.36493408301, 3440.58824222145, 3281.70588278163, 
    3063.28772790563, 2829.55400187284, 2637.11158882882, 2507.46407039906, 
    2470.37265893751, 2544.92525306347, 2665.56066518311, 2750.32071640152, 
    2789.55245219945, 2814.00585764589, 2840.90777973695, 2858.00485841671, 
    2829.3642668483, 2667.57576174616, 2270.55191960345, 1739.65932049677, 
    1263.34925892018, 881.678577116521, 586.007485622678, 375.083865648626, 
    236.320602510571, 146.191076122639, 90.9251041023366, 57.3284031190375, 
    37.3524302418679, 25.3441585345462, 17.7189592063586, 13.0430857551887, 
    10.8180111709486, 10.134317589676, 10.0116261986514, 10.0003634929987, 
    10.0000077554596, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3802.15204034138, 3802.15204034138, 3765.37841647344, 3695.28613457666, 
    3591.98235145781, 3465.6869152746, 3325.52728755556, 3158.99436835873, 
    2950.15257112809, 2728.00079121552, 2538.10336899804, 2403.79224667504, 
    2369.80785373108, 2466.29852420229, 2616.84642755758, 2723.12301422135, 
    2772.9972479066, 2801.39109430931, 2826.50783475358, 2836.21006000407, 
    2799.3461496401, 2635.38896832646, 2242.69427422312, 1712.73200389932, 
    1234.05471749743, 863.135349584512, 580.14021345108, 372.145411064465, 
    234.088969871937, 145.360034676313, 91.1085020748485, 57.8197958120538, 
    37.5484813533953, 25.2773242726104, 17.6758885870166, 13.068173079907, 
    10.8459652836869, 10.146477390609, 10.0148185461538, 10.000754886756, 10, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3778.79804664165, 3778.79804664165, 3749.51731090375, 3673.54179673781, 
    3547.95752239168, 3401.30301800498, 3250.04604783059, 3080.35133726789, 
    2874.73340300715, 2652.60001972522, 2461.80935754064, 2346.00433934281, 
    2340.74775561861, 2444.8267981641, 2588.28823886034, 2696.59827242508, 
    2754.96417188183, 2784.71065685748, 2801.44717945349, 2799.86693885243, 
    2755.25156495193, 2591.69398952333, 2210.95913516617, 1694.50290515394, 
    1218.42463872552, 851.521640458071, 574.90267282433, 368.662331793596, 
    231.39046020866, 144.588940642391, 91.3151914610899, 58.0951746126923, 
    37.5617429706909, 25.0859508418192, 17.4454620269941, 12.8870792776797, 
    10.7646489808304, 10.1252404242766, 10.0111946193702, 10.0004077381162, 
    10.00001021067, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3775.75040791738, 3775.75040791738, 3741.07336528078, 3647.74614660853, 
    3505.19457721095, 3358.7677354454, 3211.53441498699, 3035.32872085853, 
    2825.02480738228, 2612.29454028369, 2450.48882910879, 2382.20482743985, 
    2408.07134722317, 2491.28885594068, 2591.2435670627, 2678.71649033686, 
    2736.43831046074, 2764.15425642932, 2771.70247040671, 2761.04008684235, 
    2709.92135043171, 2539.29237224339, 2157.99471976666, 1650.47990524466, 
    1181.65780962268, 821.827098054605, 555.031993283505, 356.811640410843, 
    224.248164734375, 140.816453305406, 89.1263373423167, 56.6274641078605, 
    36.575325548786, 24.3992077521229, 16.9555841202019, 12.5605295559016, 
    10.6256451085232, 10.0939515003336, 10.0082518048884, 10.0004013520705, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3774.30511713892, 3774.30511713892, 3722.02640881132, 3605.41496372113, 
    3451.58898334925, 3312.19679722677, 3172.67559623672, 2994.80101367257, 
    2793.77998452109, 2620.47657089486, 2519.20931071974, 2499.44239741186, 
    2528.98933732804, 2568.85861413317, 2614.02226648085, 2667.6995882277, 
    2713.38178167589, 2737.22233270413, 2740.15343597967, 2721.52909247901, 
    2652.04718110552, 2449.09415721091, 2047.70891556169, 1548.70978045019, 
    1096.34821832724, 748.902504035678, 498.954798698815, 321.117181967121, 
    202.889334595096, 127.623465685258, 80.536246372159, 51.2392610399217, 
    33.4764074806315, 22.7593612192297, 16.1248213438673, 12.1854695927934, 
    10.4943208558286, 10.0639125527817, 10.003890674263, 10, 10, 10, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3742.40937917281, 3742.40937917281, 3667.69075306153, 3528.27410023643, 
    3371.07941690616, 3247.55436341361, 3125.9853104461, 2967.26750473498, 
    2807.34210342743, 2695.15554399751, 2644.18742684887, 2638.16198709892, 
    2643.98038120119, 2639.72551657288, 2638.55931407973, 2657.15506296265, 
    2686.67163136688, 2708.45186909086, 2710.59432879473, 2682.28908123772, 
    2581.24081035262, 2321.76704424462, 1883.59757088458, 1394.30263904459, 
    974.27632570438, 653.548843780523, 427.569942456387, 274.236644860368, 
    174.074694317573, 109.879597521087, 69.3922829327741, 44.5589996490174, 
    29.5673381041828, 20.5462905163687, 14.9761426442559, 11.8200462381412, 
    10.4197005037409, 10.0514105035682, 10.0030731138246, 10.0001515995651, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3678.16706666471, 3678.16706666471, 3583.1160127628, 3419.68120110938, 
    3258.44143191066, 3160.59244636033, 3077.50086962804, 2962.86082775365, 
    2862.54632466184, 2803.70451593646, 2765.93473287466, 2738.68239844681, 
    2713.2354872079, 2677.48856314253, 2644.37821930449, 2636.89874970066, 
    2656.5345246997, 2681.2150274215, 2685.42970320551, 2647.17720795862, 
    2509.10193124951, 2186.15419201617, 1712.04226026979, 1234.8336194334, 
    854.655321566952, 567.513976303326, 364.695214906096, 231.157001123888, 
    146.532970017859, 93.006650417408, 59.1388770168702, 38.6344737926224, 
    25.9440851325094, 18.3545612424267, 13.9577118579068, 11.8229992606818, 
    10.5904440576501, 10.1023153257052, 10.0072103617416, 10, 10, 10, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3622.09305312564, 3622.09305312564, 3513.76371953439, 3328.96359973774, 
    3158.13340086309, 3080.8872902217, 3037.9168517577, 2966.38732203885, 
    2908.49674186499, 2875.07392406226, 2830.70040541757, 2780.20857818542, 
    2733.93431995471, 2680.96660286269, 2631.30069423572, 2612.02933430543, 
    2630.16699876587, 2660.16377423538, 2668.13889771827, 2625.35782064925, 
    2464.39136222717, 2102.99587955717, 1609.87547148693, 1137.52055598363, 
    779.499670452809, 512.842704047382, 323.574143185544, 201.987686189467, 
    127.708746679929, 81.6421785162741, 52.3561318136806, 34.754320370818, 
    23.5644375662486, 17.0099337252208, 13.5588512666172, 12.2295888913736, 
    10.9841414746609, 10.2366097670953, 10.0288442602251, 10.0014422130113, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3622.09305312564, 3622.09305312564, 3513.76371953439, 3328.96359973774, 
    3158.13340086309, 3080.8872902217, 3037.9168517577, 2966.38732203885, 
    2908.49674186499, 2875.07392406226, 2830.70040541757, 2780.20857818542, 
    2733.93431995471, 2680.96660286269, 2631.30069423572, 2612.02933430543, 
    2630.16699876587, 2660.16377423538, 2668.13889771827, 2625.35782064925, 
    2464.39136222717, 2102.99587955717, 1609.87547148693, 1137.52055598363, 
    779.499670452809, 512.842704047382, 323.574143185544, 201.987686189467, 
    127.708746679929, 81.6421785162741, 52.3561318136806, 34.754320370818, 
    23.5644375662486, 17.0099337252208, 13.5588512666172, 12.2295888913736, 
    10.9841414746609, 10.2366097670953, 10.0288442602251, 10.0014422130113, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10 ;

 hraw =
  -4366.50239121825, -4335.35746684726, -4427.10886388705, -4526.04944739549, 
    -4561.55841726347, -4552.84754933129, -4521.64290903755, 
    -4486.80463318586, -4464.49464088212, -4483.71168453245, 
    -4552.44244640719, -4578.94571895624, -4546.7186531714, 
    -4536.14896572379, -4544.47560195782, -4535.4838439057, 
    -4480.66701451313, -4418.1575551887, -4408.64247350954, 
    -4436.35678205475, -4445.2174709372, -4375.46456956896, 
    -4313.50418059949, -4314.37994570519, -4273.14286289598, 
    -4224.20583816325, -4256.05756154934, -4278.82294639798, 
    -4260.34571799248, -4265.32011133082, -4276.62081977215, 
    -4256.74164327314, -4197.09390592453, -4118.43541971945, 
    -4055.09516491712, -4026.39350295586, -4016.74084156003, 
    -3983.26678210761, -3937.8244551023, -3902.06393621947, 
    -3870.56713605585, -3795.20454404039, -3645.50859435813, 
    -3540.21140816848, -3513.81774775605, -3482.9369029039, 
    -3455.70488521883, -3409.21487861364, -3198.6737222268, 
    -2829.20614028059, -2433.42612223143, -2192.29627210657, 
    -2049.3736272387, -1693.31932390848, -982.029244419679, -30.9726630718608,
  -4579.44552316509, -4525.06495953447, -4490.72949669587, -4533.82468773951, 
    -4634.06536160069, -4681.16531935869, -4634.55193948512, 
    -4535.63276572091, -4515.64050020128, -4557.76448925327, 
    -4573.07743338784, -4590.92361823576, -4589.17518891246, 
    -4492.58030849461, -4444.78380432004, -4521.2355047258, 
    -4513.52103888952, -4405.5471780174, -4319.06056174139, 
    -4322.66738886586, -4377.16072243321, -4364.14594128675, 
    -4352.25533085363, -4375.84275228597, -4278.32041963193, 
    -4149.96573352752, -4170.33616635177, -4204.25204656451, 
    -4185.26991509333, -4189.97018757125, -4212.37882189876, 
    -4208.16908925865, -4132.10027233307, -3997.98583121168, 
    -3870.94436873964, -3850.63205320052, -3920.26953147719, 
    -3944.72399356659, -3930.05874474286, -3913.98754840979, 
    -3880.95588434728, -3782.36911923863, -3608.68379594551, 
    -3540.3565006592, -3586.55675921707, -3539.58329447307, 
    -3347.37035479163, -3045.36757683287, -2712.00728159871, 
    -2434.5720140773, -2284.71627064922, -2262.25195334782, 
    -2092.74782999649, -1334.83051173427, -350.165433207007, 378.674442266643,
  -4684.36976556611, -4600.43310887537, -4556.09670864705, -4582.56854250453, 
    -4662.88278034068, -4727.6111525565, -4694.76078347702, 
    -4574.23460329554, -4545.44250434354, -4599.59235313104, 
    -4625.11796216073, -4638.93534939028, -4631.60571347757, 
    -4553.74063105915, -4494.93542129289, -4512.70646124958, 
    -4499.97761318622, -4400.59169207036, -4244.576423828, -4190.28171287391, 
    -4258.35457195882, -4308.11307632999, -4365.68731668937, 
    -4431.56886092963, -4344.22339540602, -4193.00072609595, 
    -4170.16823689938, -4196.17043555786, -4198.11899618081, 
    -4179.13299358085, -4148.74943814046, -4102.31159042893, 
    -4013.32931668609, -3945.42465634125, -3976.91930190784, 
    -4023.08907142524, -4032.08325703663, -4024.21437910627, 
    -3985.69895451177, -3921.01146697551, -3889.42855859101, 
    -3836.46442784673, -3696.62604264662, -3638.15162345249, -3635.246775474, 
    -3426.22209640716, -3017.59838083546, -2537.34562122975, 
    -2133.6822697198, -1935.38479708542, -1976.17847459815, 
    -2012.68181838544, -1729.98465978197, -889.987545787393, 
    175.363684326935, 985.362291490994,
  -4697.07760506537, -4631.27935257165, -4619.18204801187, -4640.91582211168, 
    -4673.76973397041, -4706.13374296005, -4676.56537698174, 
    -4577.00318024001, -4532.23975006885, -4563.92675197045, 
    -4616.49132771834, -4645.04442476618, -4622.62233299876, 
    -4548.8158368865, -4480.57512808514, -4457.38063688033, 
    -4440.52747202658, -4364.60643429504, -4207.9102006218, 
    -4135.46258263311, -4202.97098918329, -4305.08160799523, 
    -4393.75017421053, -4434.56631029983, -4376.57254642024, 
    -4256.79095093232, -4163.7895752116, -4151.38858318232, 
    -4187.91546048842, -4170.72656381081, -4107.64944174067, 
    -4037.49960758477, -3975.01169194897, -3967.01078796765, 
    -4043.50520134332, -4098.36350591422, -4086.88470282358, 
    -4057.86843663306, -3998.43172843815, -3917.36075476411, 
    -3903.71336998782, -3897.39811455298, -3796.26355703871, 
    -3713.06771107856, -3526.8263666899, -2912.23024237937, 
    -2265.52812966751, -1960.2505109295, -1785.10990359731, 
    -1693.48564108172, -1708.94300593584, -1561.86724466993, 
    -1093.88402009536, -358.413452377677, 509.937779922028, 1235.81229947403,
  -4677.46937751464, -4662.86814530245, -4671.88327201197, -4677.3180717393, 
    -4665.18921071001, -4648.21507850126, -4612.48143600927, 
    -4554.99522126549, -4514.13477515911, -4516.44303537464, 
    -4561.28858485285, -4593.71006182329, -4563.9482392989, -4459.1447062053, 
    -4377.65099620752, -4378.01004729042, -4364.67450453815, 
    -4308.44154565127, -4242.85176177432, -4220.12097626979, 
    -4255.40321003604, -4314.83013056875, -4348.80873627713, 
    -4339.06565161058, -4330.43082424691, -4278.36079428623, 
    -4137.69167384301, -4080.05383766484, -4136.31711197953, 
    -4147.85009849959, -4107.70678754262, -4067.36226671777, 
    -4062.39593796999, -4052.82664729724, -3990.95301775912, 
    -3970.59164376705, -4004.65313748558, -3994.9178624802, 
    -3942.95625730744, -3896.74293168826, -3905.61459757192, 
    -3918.24857840296, -3837.33689061697, -3636.73506491096, 
    -3143.85804576959, -2154.74564012013, -1425.78625891939, 
    -1479.5842917936, -1685.63629428205, -1734.73007730144, 
    -1596.48867067138, -1149.40505143171, -454.691025231615, 217.41980209503, 
    739.164379449586, 1009.50003723066,
  -4675.23591034929, -4660.76719980676, -4698.87293901464, -4690.33563419036, 
    -4622.15355164196, -4590.4445813158, -4576.31407772702, 
    -4553.41809639109, -4566.92817788096, -4592.74001648359, 
    -4577.62213652382, -4547.67081459646, -4514.03062298142, 
    -4458.18806637821, -4405.66938019169, -4371.11729570766, 
    -4319.84054298073, -4293.91683213257, -4348.55226566095, 
    -4393.13145125178, -4341.39026613857, -4177.80700891814, 
    -4074.05302628625, -4143.92802783362, -4252.03104987838, 
    -4278.01098000549, -4186.64322988282, -4129.13773922511, 
    -4154.51512218341, -4164.93714270327, -4156.69507303138, 
    -4158.92081771673, -4181.98994586535, -4175.80227213178, 
    -4090.93621769649, -4013.63194431035, -3981.4790725253, 
    -3948.09949941763, -3897.49373871877, -3849.82267828369, -3860.825077465, 
    -3890.02111161884, -3789.83856047361, -3289.64863832156, 
    -2440.33351068484, -1668.90602238586, -1277.61205075809, 
    -1329.92425919282, -1541.66951938715, -1670.67460165795, 
    -1531.67379526407, -954.072783296094, -54.6676442253714, 
    735.109407779365, 1042.99385226616, 771.823030973157,
  -4646.56980695799, -4619.83883619775, -4693.9945710564, -4745.27614795819, 
    -4700.50241784248, -4594.50801814633, -4521.00580550014, 
    -4536.07509449432, -4582.65031449476, -4598.71075226559, 
    -4553.03107855264, -4500.43626710931, -4477.71515843073, 
    -4474.62033773427, -4446.75750104947, -4383.78337155118, 
    -4356.04919849528, -4323.52704951768, -4230.60107056314, 
    -4238.07590813282, -4292.10722237194, -4123.7769421265, -3982.9970001151, 
    -4093.32458099988, -4234.7761772999, -4294.82029618548, 
    -4282.15754288692, -4252.29914290707, -4235.51211596231, 
    -4224.28653888935, -4223.10767989185, -4232.48906874745, 
    -4236.00867285396, -4234.05689676583, -4224.06726475882, 
    -4151.98698821809, -4024.26800743711, -3917.98304737835, 
    -3841.76612078418, -3810.2712950516, -3876.19926405888, 
    -3868.80029597632, -3547.2, -1832.29783217343, -1704.5000799936, -1142.7, 
    -1157.39790416767, -1104.99849612031, -1888.9, -1684.69999200064, 
    -1201.99972002239, -640.6, 308.999440044799, 670.998960083151, 1410, 
    594.55757228372,
  -4569.35660879148, -4572.26153302757, -4676.07088086218, -4810.43710581778, 
    -4834.56933914604, -4624.41177983909, -4447.98370434141, 
    -4487.87962387644, -4485.06060587598, -4417.67666720715, 
    -4411.34891249721, -4429.20900688653, -4432.4915586333, 
    -4420.46428148617, -4389.6649015632, -4374.4132491022, -4457.33976273422, 
    -4371.98400190084, -3896.843212729, -3765.05781219527, -4117.61934872834, 
    -4292.01260114888, -4288.22986689244, -4293.56416103121, 
    -4320.4556475083, -4354.99934586895, -4377.58134411512, 
    -4364.52405801834, -4325.71984761522, -4301.87702019208, 
    -4281.07762113736, -4244.71968026313, -4204.28095574644, 
    -4194.72205992437, -4228.78919174642, -4199.21481577515, 
    -4066.32800819692, -3899.32861884896, -3783.06958176682, 
    -3784.48033500774, -3830.49947204736, -3804.30028797696, 
    -2077.49429645629, -416.299983974404, -1582.49803223998, 
    -698.598784097274, -1704.20026396544, -1129.18251414188, 
    -1441.59951203904, -1599.59876012863, -1275.29993601922, 
    96.0025597952117, 613.997040332763, 1031.98432159313, 1479.9996800256, 
    391.551539942577,
  -4531.7077476706, -4591.5595076082, -4700.50487105803, -4656.08759154873, 
    -4487.5344415001, -4476.67962837448, -4530.32432034073, 
    -4495.31812359929, -4400.71556374405, -4322.67006672181, 
    -4321.78570867929, -4345.58574959135, -4358.36902064848, 
    -4370.86510598444, -4391.17581608243, -4429.83348951071, 
    -4492.07410467317, -4411.54699797769, -4080.02845596448, 
    -3971.60163656104, -4198.8001678607, -4371.17040137357, -4423.219685554, 
    -4421.62108339466, -4419.5080846355, -4443.79725525816, 
    -4483.33883597829, -4457.10391407918, -4380.39311499204, 
    -4365.80152862349, -4341.47376360088, -4251.42445950768, 
    -4204.94225617744, -4201.25364238017, -4173.2393573662, 
    -4125.55967306367, -4114.50042396608, -3928.19920806848, 
    -3883.50024798016, -3806.39989600832, -3806.1001919872, -3512.4014880595, 
    -786.700327973762, -922.198312178545, -345.000599896972, 
    -516.201503879687, -1090.90473521161, -1001.39781588612, 
    -236.502375809931, -1154.80025598016, -104.801903774819, 
    53.0013598912062, 547.008639513592, 1086.99864012154, 310.000959923204, 
    114.496697178,
  -4597.47408561671, -4686.44271368907, -4768.29603385921, -4528.12632171439, 
    -4187.95904257824, -4440.21951483234, -4754.78274669201, 
    -4618.09557306969, -4468.14791555821, -4437.657910619, -4411.51914589114, 
    -4388.14473233919, -4389.07174725903, -4427.78406465831, 
    -4484.37896609526, -4519.10099908748, -4488.33888477424, 
    -4466.36401840606, -4534.0504102332, -4525.44553943285, -4407.8095471153, 
    -4340.36179759552, -4353.36797559432, -4408.22288088122, 
    -4445.03015798222, -4480.45224472708, -4541.18580319599, 
    -4509.95584329504, -4404.65077507231, -4390.87480338709, 
    -4372.89972303596, -4274.32736533121, -4244.26487214649, 
    -4239.13940999584, -4135.23325381178, -4039.0766726301, 
    -4003.40721497062, -3963.94250789329, -3890.2000799936, -3287, 
    -3936.00005599552, -753.199224062076, -1071.6, -994.39559235262, 
    -557.499224062076, -1744.7, -452.794032477413, -1060.89857611391, -924.7, 
    -886.899832013439, -294.102791776772, 336, 889.013118950423, 
    662.998080153509, 264, -27.9029451307429,
  -4776.54361468421, -4823.40232196601, -4853.71185202721, -4788.12376498642, 
    -4720.60767991032, -4871.06486297969, -4979.95137266095, 
    -4847.16336826131, -4738.70611347093, -4716.3297034326, 
    -4692.50664466428, -4666.53818439386, -4646.34549116207, 
    -4626.96383053115, -4599.53358714861, -4566.61497460971, 
    -4553.79644148199, -4568.96659523486, -4588.2522713016, 
    -4529.72136034465, -4412.80401864816, -4364.40767442624, 
    -4372.67511363755, -4386.04820886771, -4389.88409296695, 
    -4420.8019558191, -4503.21582980065, -4514.45321633916, 
    -4434.03625541779, -4376.22773857534, -4343.7198958179, 
    -4308.12222498173, -4270.42593815447, -4224.58337707847, 
    -4157.64274741506, -4057.8262058819, -4130.5007599392, -3893.699632032, 
    -3748.49974403136, -2781.49783217343, -2190.39345649853, 
    -878.000959917445, -987.3, -82.999952008959, -838.400175849623, 
    -473.295448364139, -1308.7991760544, 39.0059197119974, -748.999640028798, 
    -357.596328371171, 31.0011998400532, 234.001839852808, 1048.99600042876, 
    563.012959282884, -64.0000799936004, 188.738658516994,
  -4980.10083072032, -4984.40397697066, -4973.55583217645, -5045.70557250165, 
    -5171.49544565367, -5182.36236973378, -5106.36448243076, 
    -5030.29196449797, -4994.9569175697, -4980.96703304494, 
    -4948.03028996884, -4910.71661403001, -4860.72800135447, 
    -4764.16152411512, -4675.28106011768, -4648.50225724861, 
    -4666.62190752203, -4661.06915460481, -4575.00987002428, 
    -4490.45817100292, -4456.07361055948, -4449.88933092588, 
    -4459.07080291351, -4471.64469158149, -4470.78317597354, 
    -4480.41770276834, -4526.26181414498, -4545.11697283621, 
    -4492.92060388422, -4384.23766848133, -4327.13586619898, 
    -4358.98941423011, -4326.21156522334, -4246.06382766295, 
    -4201.66099309592, -4060.02475287311, -3831.60003199744, 
    -3646.69992800512, -3547.20003999616, -3274.10037596992, 
    -1181.60021593089, -1055.60101593088, -123.89995200384, 
    -1841.40027196992, -1151.20124784769, -851.698120150391, 
    -761.299544074232, -587.80155985601, 11.0000799936004, 215.001759878405, 
    387.998400191948, 691.996240300783, 1300.0004799488, 312.018878637381, 
    449.001599872007, 460.113519120767,
  -5128.34003175684, -5115.8624416599, -5093.50822348363, -5097.53089233748, 
    -5128.06063902122, -5142.37401250871, -5126.84677078492, 
    -5099.79116861202, -5109.84134953142, -5112.35663059892, 
    -5039.90222438892, -4968.81033069893, -4907.9598070985, 
    -4784.43086880086, -4716.39866142545, -4769.74155997112, 
    -4774.51115016396, -4722.13181943344, -4699.42548055088, 
    -4682.81246889618, -4641.93663953415, -4578.15646902801, 
    -4566.73267955896, -4635.82953222611, -4674.98489314166, 
    -4658.87891524762, -4625.94709001198, -4596.92302117517, 
    -4542.49097748476, -4410.95370422642, -4338.23912377606, 
    -4392.14813186563, -4380.58939491802, -4290.41385664181, 
    -4199.54569176974, -4018.16851426325, -3803.8, -3564.99964802816, 
    -3231.80039196864, -1955.7, -1420.99977601792, -55.3009279257642, -21.9, 
    357.996160307182, -349.985833133375, -151.6, -60.4999680025599, 
    50.0018398528084, 270, 210.0000799936, 292.99936005117, 993, 
    704.999600031999, 1212.00335973136, 1330, 556.250412026343,
  -5189.50514430238, -5143.92900500714, -5130.67612486894, -5115.08267239583, 
    -5093.26053427595, -5104.44931000762, -5119.93890658796, 
    -5117.01219661838, -5130.64731829572, -5108.65682046215, 
    -4993.27737080247, -4920.83921744479, -4909.87361074754, 
    -4832.59277091863, -4784.44354119426, -4833.153300163, -4830.75945122308, 
    -4786.52263086127, -4793.73086853798, -4811.37465302495, 
    -4792.47529416052, -4729.06726361912, -4690.67938108406, 
    -4715.3964911671, -4727.33250071056, -4696.91716667864, 
    -4638.12773129207, -4575.15052754337, -4498.73491287484, 
    -4379.20474475387, -4311.84475250453, -4340.14656587848, 
    -4320.98407138902, -4219.20677489046, -4096.60434451181, 
    -4010.9001919776, -3895.70029597632, -3731.10002399232, 
    -2246.20223982337, -1142.2003599712, -534.498880115191, 
    -330.599208069755, -533.499864010879, -65.7998160153591, 342.9896811583, 
    438.991440684761, 615.001920006383, 622.005919200079, 1689.00647948163, 
    2011.01775840011, 991.003919654498, 2204.99744020479, 1234.00031933449, 
    772.998800070354, 1054.99296056317, 506.14969096021,
  -5218.23548232241, -5146.81969778041, -5129.25035479205, -5120.91850189264, 
    -5101.19937350955, -5097.91329375989, -5111.21417173946, 
    -5129.8875231159, -5140.4091337492, -5088.61674583438, -4947.50896961866, 
    -4872.14536133537, -4891.41057574562, -4871.5953966931, 
    -4840.61144651247, -4844.60191327178, -4839.36355497734, 
    -4822.99177064874, -4821.48568570808, -4833.56815322278, 
    -4837.58847707343, -4803.79248256332, -4754.28533480959, 
    -4716.80243284688, -4689.19231315199, -4654.61815284438, 
    -4595.65130746923, -4518.77146092993, -4427.3935017401, 
    -4323.24323842346, -4256.10805433425, -4241.74884424264, 
    -4198.48799115927, -4102.40487900108, -4070.79984800512, 
    -3928.09880807424, -4022.8992400608, -1379.20064825851, 
    -690.100231991679, -517.201711863048, -37.4999439942414, 
    157.999439974409, 436.9999200064, 1520.98016255335, 1297.02079781138, 
    1642.99360051197, 803.004320147141, 886.004879852783, 720.000239980801, 
    866.0001599936, 789.99896010874, 1074.99800015999, 1359.99704039676, 
    546.999520057581, 469.999040076796, 614.787781444798,
  -5257.92746929758, -5189.17360444471, -5141.18846893544, -5098.69723236327, 
    -5063.74745688536, -5066.02010555314, -5102.17767817442, 
    -5149.13815320237, -5171.03472250527, -5122.27007336487, 
    -4989.39924590899, -4885.72130335625, -4855.93044302087, 
    -4842.78617335241, -4834.31762506324, -4830.49215610864, 
    -4817.61517787664, -4803.44573186696, -4803.50879494335, 
    -4806.39793364284, -4795.61691312189, -4760.51107961529, 
    -4721.66874680983, -4698.63365975773, -4683.86822922828, 
    -4649.21115550992, -4571.42442476248, -4483.78395674228, 
    -4394.3745196515, -4279.52322880309, -4203.8, -4132.12486952714, 
    -4071.01321928463, -4134.9, -4060.29999200064, -4047.39999200064, 
    -3433.8, -1582.6960163187, -485.499728021759, -416.2, -23.7996960243186, 
    151.9999200064, 1336, 740.002479801611, 433.00215982721, 448, 
    1176.01023918085, 1084.00199984001, 752, 715.0000799936, 
    614.000399968019, 813, 514.0001599872, 527.001439884868, 644, 
    960.650179162879,
  -5270.32190978305, -5201.07247411982, -5139.60857447681, -5083.5437940692, 
    -5044.18053925594, -5050.98998705976, -5090.50028391725, 
    -5131.33792552272, -5142.07815144534, -5106.98644648581, 
    -5028.04617011141, -4931.55857485433, -4845.67016103384, 
    -4791.97655587831, -4774.64543806077, -4779.42536910547, 
    -4772.4968160884, -4757.99943125799, -4758.32633922763, 
    -4764.82642936777, -4757.69076035184, -4720.22185270476, 
    -4686.50816399612, -4684.23299235216, -4688.87353441646, 
    -4656.76993318635, -4560.38497092242, -4456.13883196489, 
    -4354.01704080386, -4206.00113580577, -4061.07897198855, 
    -3965.53336436977, -3889.74486243002, -3891.39922406208, 
    -3634.29997599872, -3814.79964003456, -2385.3956963443, 
    -1010.20091187329, -633.29988800832, -126.80003199744, 232.005119353661, 
    560.000480550308, 602.000159987201, 304.998560166385, 90, 
    83.0001599872007, 884.991760819137, 1148.99512037118, 749.999840012799, 
    1201.00119987841, 1134.99832013433, 968.000959923204, 858.998800102396, 
    565.0007199872, 468.001119910405, 1041.71006169519,
  -5259.54563902543, -5205.59734039812, -5150.88137372113, -5091.57123252246, 
    -5043.73277612732, -5044.36584549525, -5061.82452270086, 
    -5060.51240216043, -5049.77729126298, -5036.19556321196, 
    -5014.6788469492, -4959.40660942402, -4867.12249686117, 
    -4769.26670290901, -4721.89994643358, -4738.1643129303, 
    -4737.60232168173, -4719.41208038624, -4727.64891529398, 
    -4749.84924081959, -4756.22332914848, -4721.21018275178, 
    -4681.05468841259, -4672.22666426486, -4682.1918886592, 
    -4663.14849636339, -4571.45411040029, -4445.51475181354, 
    -4300.97809409139, -4116.99583198237, -3932.98905869673, 
    -3791.71510137917, -3784.70001599936, -3777.19997600192, 
    -3317.40083989569, -3553.20016798144, -1200.79934405248, 
    -819.099927995521, -55.9003279788807, 514.996080313582, 219.001599705634, 
    483.004159020922, 197.000159987201, 70.0001599680038, 92.0000799872014, 
    252.001359891206, 1250.99808046714, 767.999760038396, 1530.00527957762, 
    651.000080012797, 468.999840000001, 1162.99856011519, 901.996000255995, 
    86.9996000447859, 621.999440044797, 1033.32354845915,
  -5244.42074558127, -5250.14198554283, -5203.36129103571, -5112.34526203775, 
    -5025.90922894146, -5012.73141003437, -5008.41604261056, 
    -4963.74584211676, -4953.60242267676, -4970.16199070085, -4960.354303045, 
    -4940.00539305783, -4898.35372276999, -4798.42548012106, 
    -4736.26723571651, -4761.81193016918, -4746.36966278926, 
    -4710.82798573406, -4745.09259767166, -4781.8699961812, -4772.5425905041, 
    -4730.61387053505, -4681.27268992805, -4649.70365949922, 
    -4650.79216218509, -4649.90546510866, -4589.96928769698, 
    -4450.54944574807, -4254.72986695676, -4058.71856978326, -3926.1, 
    -3731.59955203584, -3482.09989600832, -3545.1, -3434.3998400128, 
    -2742.60039196864, -1265.8, -607.898408127353, 505.006879449631, 359, 
    635.996320294383, 594.001599872007, 188, 58, 78, 127, 1336.01167906565, 
    2381.00183985281, 1785, 1277.00191984641, 558.00063994883, 1204, 
    1355.00407967361, 644.001919846491, 752, 1337.81750695663,
  -5175.97526823593, -5217.71872613481, -5191.42621736705, -5104.18031180319, 
    -5009.15674944726, -4980.93311334648, -4970.99671169752, 
    -4933.72482373274, -4919.17152319191, -4929.14442388627, 
    -4934.50045891758, -4936.66753030482, -4914.33720139337, 
    -4831.96328464279, -4775.08290936861, -4790.3065873416, 
    -4767.74626850801, -4731.36497453988, -4763.14425959699, 
    -4792.60647394454, -4769.57989495479, -4708.69277054663, 
    -4648.95869385346, -4612.41299050555, -4574.12047300218, 
    -4528.72843250537, -4474.16742456449, -4363.39918344637, 
    -4197.64059834775, -4034.32215287528, -3860.20007199424, 
    -3692.09993600448, -3476.80016797568, -3433.0038236941, 
    -3121.99982401984, -1031.10575162241, -119.500167986561, 
    656.002960447904, 160.002479680031, 522.001039916805, 1200.00039980803, 
    220.997440230384, 38.0001599872007, 37.0001599808018, 66.9997600319969, 
    375.001919846409, 2612.99800034556, 2786.0015992769, 1060.9999200064, 
    1598.00191976962, 804.984401983429, 757.013438924861, 834.997680044811, 
    621.99952004478, 906.001599872007, 1426.71969081735,
  -5058.98330001019, -5097.77563457779, -5113.29619651632, -5077.79250081684, 
    -5009.6890476954, -4970.17776174315, -4959.93843737087, 
    -4954.81021216995, -4934.26091326958, -4927.68265119279, 
    -4966.1960585828, -4973.75560395208, -4919.16217657374, 
    -4848.12185483434, -4802.85636230467, -4794.42540921246, 
    -4782.57571265354, -4764.60957393303, -4759.84636312449, 
    -4761.5239101654, -4740.10089083077, -4662.3089239718, -4593.18638566696, 
    -4565.06305773007, -4481.80674669962, -4360.99833266533, 
    -4279.6050506404, -4219.57850745904, -4144.37688799436, 
    -4025.81175130768, -3920.09997600192, -3725.39917606784, 
    -3448.60067992897, -3118.09992800576, -2674.00354375105, 
    -1510.1079193274, -111.199880009599, 14.9999200063996, 748.999359859228, 
    684.001119910405, 159.999040083195, 13.9999200255966, 32.0000799936004, 
    64.9999999552072, 110.000719833621, 1112.99376049917, 2892.00607957762, 
    3783.99712053114, 1405.00415966722, 408.00143986561, 767.0128784709, 
    227.998960083195, 757.999760019199, 1086.99216035193, 1130.99880009599, 
    1236.58840786041,
  -4966.31381865562, -5018.11397698977, -5089.72476615988, -5093.3918208702, 
    -5025.97805130694, -4979.63379523513, -4943.75693222971, 
    -4903.78018253175, -4914.27320970406, -4969.67488097459, 
    -5017.76861934149, -5006.22631738866, -4935.59011506599, 
    -4862.20327511546, -4815.94457813916, -4801.03824836825, 
    -4794.97683134682, -4781.09414571848, -4755.44732618623, 
    -4735.95329307379, -4710.52897272395, -4640.35193203634, 
    -4566.51003087851, -4518.29782854946, -4444.81097311569, 
    -4346.07243489192, -4258.21971015625, -4199.88511412593, 
    -4138.4602753269, -4002.72567584316, -3557.9, -3515.09954403648, 
    -2425.99325653949, -1962.6, -517.599216062716, -91.8003359731215, 72, 
    154.999280057597, 426.998400127993, 181, 34, 50.9999200063996, 62, 
    204.997280217588, 713.011999040055, 2157, 2881.98272138232, 
    1785.00759939203, 2336, 1419.00375969922, 929.994160466924, 
    1168.17850987678, 1332.57874831176, 1433.08983516932, 1421.8837804624, 
    1347.44431586253,
  -4909.03986766662, -4959.75193408826, -5061.61207078935, -5099.88388128755, 
    -5046.88052148926, -4986.85650146632, -4919.94164065214, 
    -4856.39927435363, -4884.39666750492, -4969.67622278552, 
    -5009.68721360435, -4974.493292978, -4891.97694419282, -4829.26481904966, 
    -4800.64800168806, -4790.7013697995, -4770.78622793022, 
    -4743.92231471044, -4727.58261102457, -4711.61415273218, 
    -4678.43425739687, -4613.98319624045, -4536.39689138447, 
    -4469.78521206926, -4422.90345789998, -4371.46152561186, 
    -4288.41552457244, -4208.05197437424, -4115.62268008986, 
    -3940.3852326789, -3700.29992800576, -3403.89908008191, 
    -2173.50558365889, -618.998752099834, -92.7998880127989, 
    115.002399308891, 44.9996800255985, 768.004639596826, 491.985441529475, 
    22, 39.0000799936004, 89.9984801535879, 351.001679865608, 
    669.003279686423, 1069.99952009599, 2118.00111991041, 3657.99576161898, 
    1209.0000800064, 1517.0001599872, 2058.99176097271, 1885.989601126, 
    1610.20923956792, 1683.13516906763, 1718.23971293621, 1692.88949908363, 
    1609.41288314617,
  -4893.94830553226, -4903.67187122005, -4987.78618072258, -5053.28894168147, 
    -5041.78562266846, -4972.76562509351, -4908.73120232008, 
    -4890.78597975025, -4891.32075487885, -4906.56386368252, 
    -4930.74650570422, -4881.27308257274, -4777.87375738251, 
    -4750.20547326133, -4767.75215126293, -4760.48985573821, 
    -4712.69761335856, -4668.7913629943, -4677.94453976346, 
    -4681.48188471994, -4639.07488757066, -4561.61439386452, 
    -4483.61834731306, -4426.14026507163, -4368.86412695966, 
    -4296.27090581968, -4205.66824221042, -4115.24823224032, 
    -4017.88307029561, -3865.31578654396, -3514.00008799296, -3088.199400064, 
    -2200.89032204135, -65.6008399328038, -33.8001039904007, 
    -7.80001599744028, 229.004639628821, 286.998400191982, 27.0001599935997, 
    27.9999200063996, 64, 293.999520435134, 855.994400447974, 
    2137.01311825297, 2862.99456040318, 2811.99832013439, 2285.99936015358, 
    2271.96880266223, 1534.99880009599, 1304.9996800384, 1929.9968003264, 
    1679.25637863742, 1781.25486238606, 1814.05598487794, 1787.79209080556, 
    1736.62688617378,
  -4954.63996932092, -4931.67896998666, -4985.16296253671, -5002.68109414676, 
    -4956.20020870832, -4936.97150657785, -4938.29342146753, 
    -4931.72075475811, -4925.44332573766, -4922.63556166847, 
    -4910.16465222912, -4843.12479704755, -4753.38382063635, 
    -4744.57960120022, -4773.30971947033, -4766.18165292741, 
    -4711.4666645756, -4663.67617221086, -4676.93721753444, 
    -4668.75904805667, -4604.08706221522, -4531.34228854022, 
    -4472.68479032611, -4414.92373685846, -4305.88281531881, 
    -4166.92462332802, -4052.01353933698, -3947.46222828288, 
    -3883.2981139358, -3838.00035197184, -3602.1, -2470.79854411647, 
    -117.79994400448, 92, 375.000399968002, 4.00015998720073, 32, 0, 
    1.99992000639963, 48, 386.996320294383, 751.003039756814, 1668, 
    2427.0009599232, 3146.9998400128, 1918, 2181.00455963522, 2087.999200064, 
    1880.9260647839, 1710.38864938962, 1667.58003802793, 1765.2205911297, 
    1873.1789881401, 1800.53112908911, 1713.8586920359, 1764.21807499338,
  -4945.98153183344, -4929.75452508672, -4952.85203648337, -4911.60323860642, 
    -4824.01863422835, -4838.954065941, -4884.28972603562, -4867.97019830976, 
    -4831.83682130525, -4815.49580682346, -4825.2303290347, 
    -4796.57787293005, -4734.38343545632, -4722.65458195021, 
    -4738.48633611127, -4733.43556529127, -4697.15503648822, 
    -4659.48973205965, -4650.37588239205, -4618.6238701106, 
    -4555.78879501205, -4511.40738819265, -4467.9798050974, 
    -4384.78139681574, -4233.47781348472, -4036.65559869137, 
    -3854.10217875228, -3756.52493271871, -3764.34936814333, 
    -3733.90070393344, -3330.49854411651, -1038.88680896448, 
    -116.099896015361, 99.0035197183361, 55.0003999744026, 28.0005599487981, 
    181.991600672153, 2, 10.9998400191982, 65.0003999679927, 
    266.020478079759, 1163.01839834867, 1931.00703943667, 2945.00423952646, 
    2370.00368019183, 2256.99360051212, 2248.99720013434, 1864.00975896317, 
    1714.60952194052, 1754.33022473759, 1841.19251971097, 1982.80425206223, 
    2060.59171329643, 1872.29973276646, 1702.3882789144, 1787.14199170774,
  -4753.92116965098, -4771.74865936474, -4754.66082372193, -4737.23615105834, 
    -4720.23433951428, -4664.53049353575, -4641.34896940601, 
    -4651.92555896186, -4506.54114214485, -4377.1753587048, 
    -4523.93190934385, -4626.75233303395, -4562.81415642523, 
    -4542.72805789257, -4561.43769244952, -4558.88445008376, 
    -4544.97675797874, -4520.46776903807, -4483.7549890534, 
    -4464.16806173956, -4465.31067968519, -4453.21226533125, 
    -4389.91031979259, -4268.47179314205, -4135.01419687297, 
    -3932.84680308575, -3639.86072084416, -3762.50028797696, 
    -3675.80020798272, -3398.60113590656, -2087.70013598912, 
    -138.799808032636, 149.000480697491, 100.005359571209, 573.997519808065, 
    133.004000083151, 57, 6, 31.0000000000005, 370.997760179196, 
    740.99967974405, 1892.99863963527, 2906.00719942401, 2181.00255962244, 
    1712.00303976961, 1564.00399968001, 1193.00215993599, 1869.00183992319, 
    1720.1705388299, 1940.31399192604, 2068.32199729932, 2186.91979916685, 
    2268.93726469066, 2142.24173057394, 1954.08286241233, 1878.21571912234,
  -4772.5715835379, -4756.73685681121, -4670.024484999, -4632.95736808845, 
    -4648.8274295557, -4582.00984392544, -4515.63223559958, 
    -4492.17448425359, -4332.65137024364, -4206.65296543475, 
    -4366.64222379103, -4488.86736372153, -4436.88283637317, 
    -4400.6067064223, -4387.24345012308, -4359.33193555949, 
    -4341.77897198708, -4321.53130260117, -4280.94032442968, 
    -4288.71662689592, -4341.57032541401, -4343.57997381327, 
    -4265.80736332804, -4134.18016836401, -4014.46758544214, 
    -3829.33787128792, -3524.57351830121, -3409, -3456.39988800896, 
    -2834.60192784577, -699.8, 157.001999840009, 257.997680185589, 827, 
    441.9999200064, 505.996720262385, 17, 11, 51.999120070396, 671, 
    1104.00503959682, 1990.00231981441, 2003.92744140311, 1808.61275542019, 
    1596.41470827813, 1456.74121619008, 1417.12109379165, 1509.27318988953, 
    1792.83592717904, 2084.33837293641, 2156.98873074153, 2201.80244262974, 
    2282.48735933356, 2243.58191390146, 2110.96089297348, 1981.32995462759,
  -4835.10106786167, -4786.25272517268, -4683.95086143519, -4609.61685677962, 
    -4597.02517094631, -4599.33109743332, -4563.24419201157, 
    -4482.54387298154, -4438.23157460178, -4447.07926679468, 
    -4477.32147011198, -4503.28728485834, -4504.06937123297, -4466.095681615, 
    -4398.80617062444, -4326.89871653114, -4284.01603073756, 
    -4261.77871415713, -4240.58980402963, -4260.28088579784, 
    -4305.49303614766, -4294.64068597519, -4217.19062703603, 
    -4093.71148273569, -3943.17500267207, -3720.85450320949, 
    -3398.06487194677, -3017.89986401088, -3066.59984001024, 
    -1526.90189583297, -459.4, 226.003599257702, 651.003520044753, 
    924.992960563188, 629.988321452684, 60.0018399807888, 19.90001599872, 
    27.000000006399, 433.594104263687, 873.996400287994, 1407.018478848, 
    2280.99240077436, 1937.5314166931, 1704.23077127553, 1511.25833746911, 
    1332.6112373401, 1280.6193193397, 1446.06996907239, 1753.84509644373, 
    2004.76309524412, 2035.75262236624, 2045.97275251606, 2108.10101530704, 
    2090.28085555594, 2039.44269792474, 2031.76149635031,
  -4240.53907603643, -4360.70194996259, -4435.57592196041, -4493.08022952507, 
    -4534.57392515708, -4517.95258047111, -4490.4482656144, 
    -4501.90946234804, -4536.79218176887, -4566.35218461263, 
    -4577.86732645478, -4624.31481749101, -4692.9980243462, 
    -4695.37163539905, -4637.43920688086, -4564.15483016658, 
    -4517.66094905117, -4498.71891192815, -4487.05035506676, 
    -4484.98533803679, -4480.70863362774, -4442.51291414756, 
    -4350.54731927436, -4199.3946235267, -3991.77983294845, 
    -3607.71822071454, -2964.57181080759, -2565.79956003521, 
    -2347.00241574526, -1746.59900831808, -263.800135989118, 
    587.005519929572, 591.001599385596, 1430.00783937268, 827.999199699256, 
    91.000319987201, 36.6000559955191, 143.896160327036, 982.799488035216, 
    1569.00079993599, 1946.01711845741, 1590.0005608062, 1756.13543251202, 
    1604.97693309305, 1506.75128950385, 1327.01056624092, 1226.09918987132, 
    1336.05425381138, 1507.84228568293, 1667.51695049594, 1811.46710850144, 
    1927.49713867987, 1991.1817623675, 1981.07919785788, 1966.6111637006, 
    2004.77997067482,
  -3727.84043013123, -3960.87187162626, -4140.47582988292, -4270.42348332104, 
    -4331.01418405679, -4271.37716745341, -4230.8460199085, 
    -4295.27147810436, -4315.01424987385, -4300.19805996796, 
    -4349.85294812676, -4432.99424793069, -4475.48592026681, 
    -4415.22666221711, -4370.43661882712, -4416.19746606245, 
    -4418.65527230645, -4370.73383166418, -4341.206936093, -4309.51974479263, 
    -4267.92520311642, -4236.00688888962, -4173.01715231479, 
    -4029.69204148995, -3810.7, -3295.83231628877, -2325.70117590592, 
    -1427.9, -1041.49999200064, -996.800223982081, 659, 874.994560435175, 
    530.999280057597, 1791, 940.99336053117, 101, 43.1, 781.304263658899, 
    1954.09957603392, 1182, 2017.00295976321, 2231.00143988481, 
    1520.6136272622, 1474.63426140043, 1487.47125139749, 1403.58000061303, 
    1311.34592769832, 1315.80493921199, 1367.61738322069, 1477.34664543872, 
    1666.43603040867, 1815.90674407166, 1870.93007330722, 1885.15839335751, 
    1917.40119401724, 1989.32928247261,
  -3897.76245864223, -3992.39803555783, -4026.03994765812, -4010.08172193818, 
    -3973.46133937245, -3935.20045991308, -3893.54344024197, 
    -3842.85838909534, -3787.14023343764, -3752.60941776174, 
    -3760.58195701222, -3765.38379293489, -3682.11381301404, 
    -3454.80397609695, -3385.27079766346, -3607.74336829211, 
    -3694.03891564039, -3593.7651902258, -3504.06801624368, -3443.8080003448, 
    -3420.1441415748, -3458.28151076028, -3497.19968603179, 
    -3440.83223064661, -3314.79524838013, -2544.99948804927, 
    -2137.90451958276, -1234.19968802496, -1293.39924806271, 
    256.993600454368, 136.999520038396, 331.001119884811, 1558.99952013437, 
    972.003279737624, 228.010799001695, 135.000239961604, 336.999600031997, 
    1690.9955200896, 1626.99856012798, 1569.0003199744, 1558.99847981444, 
    1196.0000799872, 1400.57241206125, 1394.10987237946, 1437.41785150018, 
    1494.65175972314, 1492.19799561243, 1437.50545666683, 1503.20022256434, 
    1630.3244103404, 1657.76057867861, 1654.92929478521, 1684.55442175339, 
    1747.27942788208, 1860.78036773494, 2006.10582381425,
  -4018.16166320194, -3987.42639058567, -3906.14664344586, -3804.51996030814, 
    -3734.1964198581, -3734.81655113249, -3719.03125109846, 
    -3628.71191059263, -3549.33960728931, -3462.92659154185, 
    -3314.88289863987, -3200.17511477481, -3123.73752158561, 
    -2990.6339136217, -2954.21848833516, -3102.85676586136, 
    -3214.84035827653, -3158.99189799718, -2951.26479831874, 
    -2814.62151687828, -2855.61574549812, -2993.23986631448, 
    -3116.26383664193, -3125.9114211384, -3117.09995200384, 
    -2830.38734741621, -2764.22040335118, -2567.50056795455, 
    -949.910310794794, -21, 383.001759859173, 1102.01039871989, 
    1061.00280016008, 529.015838732557, 684.990640601644, 193.998720166408, 
    457.998080153629, 1779.00151985921, 1623.00111987199, 1661.00159987198, 
    1529.9998399872, 1677.00511973113, 1549.47870620713, 1484.66878196235, 
    1429.96598098507, 1450.60098721108, 1466.13414427272, 1443.40483629168, 
    1532.39218011158, 1634.86054191845, 1574.17983179685, 1526.60244709025, 
    1596.26270587915, 1717.98362796965, 1826.67098575104, 1886.39227640318,
  -3915.43871468778, -3846.07175805324, -3767.86140113457, -3703.59973871701, 
    -3676.85823097273, -3696.71856568686, -3688.14160602412, 
    -3609.31676766956, -3535.25644645524, -3412.91732322195, 
    -3171.66246806789, -3004.9079050542, -3007.62747085445, 
    -3091.04551887743, -3125.43374170679, -3089.37044583677, 
    -3164.76387102391, -3173.22531245562, -2868.39713114611, 
    -2652.90642887167, -2728.63061614849, -2913.88979666605, 
    -3058.72089574524, -3093.89329525704, -3130.6, -3099.39176570957, 
    -3107.40006399488, -3018.2, -715.89999200064, -117.400639948802, 306, 
    458.98904087675, 795.994080473573, 1842, 871.997280217588, 
    765.992240620765, 864, 1181.99632029438, 990, 1610, 1659.00239980801, 
    1855.00423966082, 1766.5641783443, 1667.72560308751, 1526.31525402282, 
    1416.98446902459, 1355.12879732969, 1348.55900477638, 1427.52701148809, 
    1506.72335190681, 1489.44465279557, 1511.21671871775, 1638.96364890697, 
    1796.5903508513, 1860.02213087107, 1791.14442269497,
  -3829.55765943175, -3742.82677126978, -3710.40544115055, -3695.92912262433, 
    -3686.97100160771, -3702.16039206123, -3647.70040378809, 
    -3488.25828235059, -3375.50805747382, -3310.59712757627, 
    -3212.22045322642, -3116.24951715006, -3083.77726201297, 
    -3151.95887209645, -3211.04828183961, -3196.93140844719, 
    -3224.90510947454, -3177.66279605977, -2899.29750023615, 
    -2683.55948738348, -2688.50254934315, -2805.59327610301, 
    -2918.53491365536, -2974.20330711254, -3031.50954469229, 
    -3089.89671140909, -3149.1999760032, -1906.69993600512, 
    -1102.80016799168, -100.899952016638, 83.9975201983957, 1066.98168254696, 
    988.991600959921, 1833.00751939841, 1780.98632096639, 1096.00247973761, 
    1196.0004799616, 1271.99840017919, 1289.00031992321, 1553.99800016, 
    1443.99928010879, 1797.99528035838, 1753.10145887375, 1773.86900744182, 
    1721.45976018152, 1595.13712413176, 1442.73524968263, 1347.92941638405, 
    1412.23489096235, 1543.80816652629, 1587.3534783096, 1622.65374878776, 
    1719.63933539325, 1865.49213516211, 1963.52814144396, 1953.39783680445,
  -3766.94359355576, -3704.62203224099, -3704.73438453279, -3668.60569341394, 
    -3606.56028970732, -3640.76294164376, -3621.93841898409, 
    -3455.08000411361, -3346.01949004033, -3329.13940282662, 
    -3314.0029491714, -3262.52017323787, -3199.57594490173, 
    -3195.23734278873, -3237.38770754254, -3277.45730566245, 
    -3262.74235068373, -3167.71205354074, -3002.28722605533, 
    -2833.80873977702, -2735.161951857, -2754.36270490901, -2831.14876799126, 
    -2900.43864265636, -2963.31810293471, -2953.86520862831, 
    -3135.2001599872, -1057.89989600832, -799.199872019194, 
    -73.2001279897603, 358.010959123032, 1263.0066389247, 608.017837913536, 
    1151.99592032646, 1039.99799989752, 884.999040000025, 1478.99776017923, 
    1684.00112003197, 1262.00039999999, 1483.00095992319, 1475.9997600192, 
    1684.00424019821, 1688.54857273536, 1797.0514665969, 1838.70515734289, 
    1679.8505449915, 1518.49529860047, 1528.78786846664, 1591.14433864756, 
    1648.93253064228, 1697.91257639355, 1692.41742940614, 1686.15960691285, 
    1817.49485555173, 1980.02192371804, 2043.38166866202,
  -3743.48175304186, -3720.38745306067, -3701.52762370135, -3595.65678282446, 
    -3472.94232246047, -3540.58238303391, -3623.06207207718, 
    -3561.50481160139, -3512.34576214588, -3483.98209130574, 
    -3400.09103363029, -3320.61298376102, -3283.84455052068, 
    -3272.12388893916, -3284.00922935536, -3300.84423246799, 
    -3262.13806210862, -3181.16282582323, -3098.64028887612, 
    -2969.8182207248, -2825.54273187035, -2782.00754775109, 
    -2817.68480680932, -2870.54677660302, -2891.4, -2892.79920806336, 
    -3097.3, -1107.8, -561.498752099834, -45.3001999840008, 582, 
    912.001839852808, 1311.00631949443, 1380, 973.99552035838, 
    1049.99752019839, 1375, 1221.0001599872, 1343.99680025599, 1442, 
    1800.99392048637, 1413.9997600192, 1532, 1751, 1899.9993600512, 1725, 
    1879.99376049917, 1808.99712023039, 1548, 1413.0002399808, 
    1902.00079993604, 1664.00732608503, 1593.93976801806, 1701.88299509988, 
    1844.92435850306, 1859.75155253835,
  -3820.29844974522, -3771.02658322909, -3675.19525285401, -3566.09522208066, 
    -3506.15378556203, -3552.12468023244, -3614.94044931638, 
    -3613.18654252001, -3587.14941728862, -3538.10992914719, 
    -3450.46835972791, -3372.8921080243, -3332.85402306346, 
    -3317.74475913867, -3314.51497001958, -3308.30208990497, 
    -3278.49054475614, -3192.89920340146, -3040.01448499315, 
    -2902.68023751249, -2817.92605433433, -2751.81134063934, 
    -2697.64538412754, -2678.69201723235, -2675.29992800576, 
    -2993.99766428477, -3092.59996000448, -1563.40099192064, 
    -234.097968103686, 403.987361427107, 537.003999680007, 1396.98944087036, 
    320.000799833623, 845.002479801604, 644.008319206447, 1490.99672046076, 
    1346.0006399488, 1303.00008, 1812.00064, 1396.000799936, 
    2009.99904008958, 1524.00183980161, 1691.9992800576, 1768, 
    1986.99871997441, 1423.0014398848, 1308.99832014719, 1393.9994400512, 
    1711.99496040319, 1707.00079948167, 1532.00015998721, 1636.9761490511, 
    1674.67608171355, 1681.09918088573, 1623.32014736657, 1501.46868604158,
  -3901.86525670945, -3822.53315558842, -3692.24299375836, -3613.95159848924, 
    -3615.12772993582, -3622.05588236587, -3621.86095497886, 
    -3614.53310242103, -3577.57869086474, -3524.01448606968, 
    -3478.39609566359, -3417.55129494009, -3348.43646398579, -3315.549317126, 
    -3309.51966035452, -3305.39922931763, -3287.18376113628, 
    -3198.30879766104, -3007.26751745221, -2861.37413360205, 
    -2815.15149963728, -2778.28569422057, -2690.61159508164, 
    -2598.92540670824, -2297.00014398848, -2940.4035516416, 
    -3086.20001599744, -1180.10077593791, -140.400088001916, 550.01567804165, 
    362.989040876968, 573.97160329598, 718.015838060873, 1069.99936005121, 
    551.011919174281, 1218.99864005763, 1302.9996800256, 1471.9988001344, 
    1524.00079987201, 1783.00151987838, 2070.00087948806, 1573.00255990397, 
    1426.0001599872, 1355.0002399808, 1463, 1397.0000799936, 
    1950.01239861747, 1272.99984005118, 1227.00159987198, 1194.000399968, 
    1455.00415965437, 1609.70550265688, 1695.54775413248, 1529.88250024605, 
    1288.01675026655, 1163.76886539463,
  -3898.79583920152, -3840.90215539596, -3763.87179846434, -3694.60952681737, 
    -3655.80918222701, -3653.29235386281, -3649.54249240997, 
    -3613.60073575075, -3560.10591579596, -3514.15875075126, 
    -3486.72618770153, -3430.02696540972, -3345.21060651481, 
    -3294.70390417031, -3285.30131653378, -3287.91499725639, 
    -3252.90893843815, -3181.40288406984, -3098.5330752102, 
    -2990.61547667381, -2903.33721054612, -2922.93533187065, 
    -2905.78826644558, -2807.98787950383, -3055, -3066.20002399808, 
    -3078.20004799616, -1173.1, -127.699840012799, 309.999440044798, 36, 
    445.005359571225, 247.006319494429, 492, 689.998720102394, 
    1429.99720022399, 1678, 1387.0001599872, 1877.9991200704, 1741, 1299, 
    1519.0001599872, 1322, 1627.0002399808, 1560.0004799616, 1501, 
    1277.9995200384, 1858.99888008959, 1308, 1156.000799936, 
    1318.00015998721, 1496.76164432912, 1429.51471633, 1145.24670373011, 
    947.082460718646, 1045.43739815693,
  -3854.83976402066, -3808.78247874458, -3742.76138497631, -3674.71619588366, 
    -3630.4645871586, -3628.84596214257, -3627.87394675581, 
    -3586.43354953552, -3513.58804364093, -3452.58710118805, 
    -3437.82294119759, -3409.15531123417, -3351.72314642405, 
    -3315.93858324899, -3292.42873355166, -3251.86697758805, 
    -3177.48143989887, -3091.50753170177, -3028.95509286952, 
    -2981.99037535408, -2955.37507084867, -2967.04389670648, 
    -2961.46680614576, -2947.03697350144, -3050.69996800256, -3064.900008, 
    -2427.69797642235, -857.39980801536, -241.699528024958, 67.0003198208272, 
    293.001279897602, 287.002559808015, 121.999440076793, 272.9999200064, 
    856.010239647958, 1113.01055918081, 1719.001199904, 1737, 
    1882.0023198272, 1320.9997600192, 1371.0000799936, 1345.9995200384, 
    1583.0014398848, 1341.00008008319, 1276.9999200064, 1263.0001599872, 
    1237, 1175.99840014079, 1386.99680025599, 1465.9995200576, 
    873.006079590537, 1161.56552706949, 1029.25840718993, 932.380525706175, 
    1000.78805163782, 1265.00379095443,
  -3824.91130090005, -3779.28128773115, -3690.82130793944, -3627.90973900925, 
    -3612.13035846605, -3597.18132258557, -3582.03012229183, 
    -3561.2457632115, -3489.48664018694, -3390.8765536851, -3324.19352157479, 
    -3294.40872791497, -3281.31760560501, -3250.32454219941, 
    -3172.5411996719, -3060.271207793, -2992.13683435146, -2944.374970152, 
    -2867.21527130968, -2872.32539115706, -2944.59195077262, 
    -2922.79825089787, -2885.19813947186, -2950.01685724464, 
    -3042.30001599872, -3057.00001599872, -2059.2085592134, 
    -927.798240140827, -417.999336048636, -106.80000800128, 71.9993600512098, 
    133.992480550445, 154.999040185635, 697.003519718346, 994.002959596971, 
    727.989840921698, 1683.9998400128, 1339.9998400192, 1585, 
    1809.99616030726, 1472.000399968, 1372.0000799936, 1299.9999200064, 
    1409.00007993602, 1585.00087986561, 1333.99928005761, 1349.9980002112, 
    1158, 1378.00111991038, 1327.0028796608, 1289.00167991044, 
    809.64425873436, 769.620257085015, 977.367867337865, 1305.15504203277, 
    1611.91131075551,
  -3841.98343955139, -3813.40923635719, -3747.03594115087, -3695.63360465808, 
    -3667.37982196032, -3615.990082199, -3581.254387245, -3583.67326476154, 
    -3540.91044540428, -3392.3614660072, -3156.11225875091, -3035.1688532966, 
    -3042.22143595922, -2962.11894925491, -2793.75541137531, 
    -2651.8176252072, -2684.40226032161, -2807.28230994835, 
    -2847.58443681844, -2874.72578235348, -2920.33214429217, 
    -2925.84494129473, -2913.94993648386, -2946.33290537739, -2993.4, 
    -3042.80002399808, -2974.09999200064, -939.3, -136.900247980161, 
    -103.9000799936, 9, 168.994560435175, 217.99784017279, 120, 
    371.009679225644, 760.000479961602, 1456, 1951.00215982721, 
    1189.9998400128, 1057, 1227.000799936, 1547.0009599232, 1416, 
    1513.9998400128, 1373.0008799296, 1510, 1471.0004799616, 
    1466.00335973122, 1534, 941.998880089595, 807.999600031981, 
    756.935164862376, 847.935582813274, 1127.12396050783, 1471.84260756179, 
    1785.28335996358,
  -3874.13083494289, -3842.25559646556, -3790.01905426436, -3750.62003524759, 
    -3716.75345419488, -3644.83235247712, -3604.57408616945, 
    -3618.09420830646, -3534.79283536818, -3282.96835619652, 
    -2926.93187094847, -2758.1299592515, -2793.77906035749, 
    -2734.05478598329, -2596.4562100797, -2517.66375750009, -2597.0526761384, 
    -2757.87378474742, -2852.12440882913, -2887.00677737668, 
    -2902.1373479044, -2925.71854412885, -2924.90011778778, 
    -2913.69130731163, -2943.19990400768, -2946.19995200576, 
    -2950.80009598144, -672.401039916802, -100.500127982082, 
    -79.1998720115196, 216.004079673607, 146.002559385672, 85.0003199744006, 
    214.997600191996, 589.993920710344, 804.004959667201, 791.9997600192, 
    1081.99880010239, 853.000079987201, 971.990480761584, 1016.00439980159, 
    1805.99136078078, 1514.9999200064, 1658.98160209905, 1721.99935996162, 
    1440.0005599552, 1630.00407905931, 2129.00655936643, 1205.0018398528, 
    1131.99704026239, 1083.99600039682, 890.004239660807, 1155.99392062077, 
    1322.996720288, 1492.0003199744, 1912.73780832738,
  -3904.82980127621, -3848.09538712728, -3776.66792906165, -3731.33377077723, 
    -3707.59036751035, -3657.79693044675, -3627.47179425326, 
    -3603.97988434431, -3406.28656493624, -3052.4337267058, 
    -2715.03119988611, -2582.6667693461, -2642.35315110197, 
    -2681.44825472452, -2694.93785796588, -2728.74160952466, 
    -2762.92327319896, -2791.3619078538, -2822.09029949916, 
    -2861.34808051511, -2896.59882256533, -2898.41723796768, 
    -2862.80171122629, -2840.3726817699, -2878.59998400128, -2857.000032, 
    -2622.20552807548, -965.400207983357, -304.999680038408, 
    -85.5001439846406, 161.998320134426, 85.0083993727294, 331.003199833599, 
    78.9999200064012, 359.004559622343, 1201.99080134398, 1110.01607871335, 
    1595.98952094084, 720.999040134413, 853.000159987198, 1088.99368075521, 
    853.002080063946, 1218.0063994879, 801.994000492778, 1466.00415951365, 
    1395.00535957112, 1246.99840017283, 1341, 1276.00391968634, 
    1219.00152007035, 1540.00607873952, 1645.00367970554, 1279.99336069762, 
    1318.98896126681, 1662.00431965433, 2028.50414283154,
  -3942.90074841906, -3884.73598553979, -3796.12794397958, -3709.78479259031, 
    -3659.70187976242, -3659.06794505621, -3629.84980869618, 
    -3488.3599656508, -3216.43676349694, -2898.29221992903, -2659.6851885176, 
    -2547.12767162026, -2555.44151683661, -2638.89902726903, 
    -2742.8318196195, -2817.03122341886, -2830.31965679182, 
    -2817.34786179727, -2835.66025109227, -2873.14191398304, 
    -2899.84666833977, -2886.04053632214, -2822.94629263335, 
    -2763.08855369393, -2783.4, -2777.7999600032, -1947.20362371009, -955.7, 
    -421.200487960962, -182.2000799936, 34, 439.994640428775, 
    56.0001599872007, 42, 170.001839852808, 1018.00975921924, 946, 
    1025.99736021119, 808.000159987201, 1003, 990.000319974401, 
    951.002719782412, 1363, 1249.000399968, 1006.00199984001, 1073, 
    1536.00743940483, 1917.99872010239, 1045, 987.999680025599, 
    1620.9956803454, 1526, 1343.9991200704, 1288.99904007675, 2267, 
    1985.99702953563,
  -3946.65953806891, -3888.37076500739, -3803.79940498409, -3709.2370840794, 
    -3630.64611090869, -3586.45395889249, -3504.84214660942, 
    -3317.9904896191, -3041.38064959675, -2784.64819650039, 
    -2647.76098905549, -2507.16697644115, -2396.39076673986, 
    -2522.72014978005, -2716.19136367258, -2786.45004513725, 
    -2796.5270900615, -2811.83219490977, -2858.37876213389, 
    -2890.29955985506, -2886.64698239609, -2865.33428612295, 
    -2800.53649235762, -2706.82386804774, -2589.39996800256, 
    -2628.19978401408, -1640.6061365125, -1446.6001599872, -484.099488061435, 
    -200.300287963523, -21.887848972139, 240.014158182553, 316.999840083196, 
    76.002319814404, 132.992160927922, 127.999200083195, 779.984001279972, 
    1624.00839946879, 715.996960160011, 757.990160787183, 742.999280038402, 
    785.995680723118, 545.001279897602, 743.999919942413, 1066.99488051197, 
    1033.9972802176, 1493.99904014719, 1120.00615925766, 829, 
    1949.98952032646, 2478.99696033931, 1379.99680025599, 488.01031834895, 
    963.003599481239, 2143.98984081278, 1835.87510920124,
  -3893.70870572228, -3817.88095760051, -3764.89993936897, -3720.81525731692, 
    -3631.8115968691, -3439.56905673127, -3267.73556104612, 
    -3167.09020443843, -2934.05053516628, -2663.45551899385, 
    -2546.87673849276, -2358.12386227074, -2167.04776848897, 
    -2373.15359133687, -2680.70396515743, -2762.48697363676, 
    -2766.12848821548, -2790.51001120397, -2844.033986486, -2866.55332398216, 
    -2842.3925436863, -2814.0009658934, -2767.54657260173, -2680.24132356748, 
    -2501.60013598912, -2243.00125643574, -2081.60026397056, 
    -1627.60011199104, -360.599192108792, -151.100319966719, 
    -47.5997760179234, 351.002878944284, 377.003599462412, 247.997600192037, 
    60.0000799872014, 241.995040511964, 238.003839692741, 891.993120575853, 
    331.001119839973, 261.99024078095, 372.002079878375, 395.994240569642, 
    220.000239980796, 213.002399808011, 243.001519865584, 304.002399807963, 
    406.001279891185, 1036.9774420417, 1195.99624030086, 1097.00000008959, 
    1459.00063975684, 1295.00119990398, 1334.99768000629, 757.016638310663, 
    1636.00487960953, 1642.21450240096,
  -3837.66784162251, -3763.9176683439, -3763.16550593624, -3717.97841658618, 
    -3569.95457102244, -3374.20476185172, -3207.27883819991, 
    -3082.92193001845, -2891.12952989984, -2633.52000903718, 
    -2389.06706124599, -2210.88237626729, -2180.72336756831, 
    -2377.69844424413, -2617.06325440598, -2728.07430070144, -2766.485406165, 
    -2787.64604218512, -2813.75077286143, -2815.69021401148, 
    -2788.47872657961, -2761.84836894617, -2732.55988294796, 
    -2671.82669192259, -2567.5, -2240.09969602432, -1655.70232781377, 
    -1280.4, -201.799704023679, -125.50002399808, -29.6, 238.999440044797, 
    158.999600031998, 311, 260.002559795212, 143.000479961602, 944, 
    1069.00351971842, 548.999760019199, 1070, 1064.99680025599, 
    973.000159987201, 459, 203.000319974401, 246.000159987201, 190, 
    168.9999200064, 295.999760019199, 1048, 1215.99632029438, 
    871.002879769736, 933.42047301691, 963.674807740369, 977.209435771568, 
    1084.12890784594, 1356.01289899134,
  -3826.41792866438, -3768.342718734, -3795.1217152408, -3698.90591512845, 
    -3476.20137357516, -3365.96139051863, -3264.25538147365, 
    -3053.02106014547, -2844.81104919955, -2610.24598618413, 
    -2306.61685116086, -2226.49052534623, -2392.77320344125, 
    -2494.05557068863, -2566.04162299693, -2690.66757824698, 
    -2769.31159350953, -2784.3959486376, -2778.57765994373, 
    -2764.36631793783, -2743.30264747296, -2715.15876784678, 
    -2698.37592965202, -2675.82076401149, -2599.3999200064, 
    -2347.29908015357, -1805.8021118112, -1227.10078393727, -858.30020795836, 
    -90.6004239334482, 8.00111991038284, 7.00000000639898, 559.998720204859, 
    230.002399807963, 188.998480185621, 984.985601299284, 1140.00223982077, 
    725.997920288012, 1401.9989600832, 1123.00223982077, 298.999440038406, 
    228.000239974401, 232.000319974395, 487.000879865597, 122, 
    178.000239980796, 314.004079481602, 466.001359923168, 640.001519878377, 
    670.011998995069, 912.986401407677, 779.787924193791, 935.18699552404, 
    894.762383888846, 883.092435083269, 1146.77921603668,
  -3870.4595796952, -3811.03867200388, -3795.42217939812, -3664.59120645684, 
    -3431.33993924243, -3307.09176990446, -3215.87490476165, 
    -3027.72410909892, -2744.27126003413, -2493.49510866326, 
    -2421.93642281962, -2480.224617617, -2561.54621889681, -2570.08514653333, 
    -2586.3454231712, -2673.60817553179, -2734.90113932244, 
    -2746.54872763774, -2741.42001309565, -2732.62878675971, 
    -2711.37906549028, -2662.6039657676, -2655.63698859529, -2669.422656219, 
    -2601.2998400128, -1951.40208780863, -1908.20073592512, 
    -1028.50186385085, -150.600071990398, -70.9999760019205, 
    -10.3000559955191, 22.9998405055459, 445.992880627258, 53.0000799935988, 
    527.99080116481, 962.997521183758, 1054.00175985917, 1455.97592213128, 
    1561.99599992332, 877.009919206248, 547.999360076793, 646.002319788783, 
    376.003679705544, 153.999999993599, 240.999920006401, 301.000479961593, 
    372.002159795178, 267.009599097634, 307.001119910383, 440.002879827202, 
    762.000479993588, 820.923050347278, 931.293064935669, 957.53689710617, 
    1017.18171290567, 1216.20701434571,
  -3887.49776896738, -3809.82283249989, -3723.05957319541, -3565.70470762992, 
    -3369.92071175813, -3260.41395773558, -3156.66469957893, 
    -2964.10393366077, -2727.51287910173, -2583.12487470001, 
    -2634.31188879417, -2700.3011405924, -2683.46586690855, 
    -2647.41471690981, -2635.57048984682, -2659.55178626743, 
    -2692.14619560327, -2714.23602420757, -2717.9430904386, -2704.4996993397, 
    -2667.51085401341, -2601.87431236363, -2578.07695569112, 
    -2556.38948121007, -2530.5, -1833.80015198784, -1854.40029597632, -415.6, 
    -103.19998400128, -40.8003199744012, 10, 20.9999200063996, 
    78.0027997760128, 70, 85.9997600191989, 229.998960083195, 463, 
    1607.01111911045, 1533.00311975041, 1703, 599.998800095995, 
    607.999600031998, 170, 354.9999200064, 320, 369, 549.000719942403, 
    543.000559955203, 496, 600.9999200064, 741.999040076755, 
    869.764520649618, 926.717598359729, 1031.65184825422, 1186.00212695138, 
    1342.24602322975,
  -3839.47376390341, -3736.45774828774, -3608.93772227138, -3410.93872088301, 
    -3218.26075360314, -3195.68433556816, -3131.03738901321, 
    -2903.17440533884, -2827.15423089608, -2867.74991409888, 
    -2811.64852284031, -2761.58062095102, -2758.94299224915, 
    -2714.58917214364, -2651.98173972255, -2625.40804384504, 
    -2653.5204950213, -2698.46875572708, -2704.29735065293, 
    -2674.75929043075, -2622.83888613203, -2557.02145971339, 
    -2483.84341289434, -2344.02479543712, -1929.89730421572, 
    -1579.28032189693, -1537.30003199296, -1232.20035997119, -97.79996000384, 
    -15.3001599737646, 79.9986401088208, 227.997760313579, 435.987760505909, 
    116.000879929587, -0.39999199935985, 112.99728001286, 226.998480121623, 
    776.002719398488, 917.99936007669, 1500.98528117783, 1041.01215884782, 
    712.991520691256, 300.998480121623, 678.001919852762, 424.000159987198, 
    499.000559955191, 487.000000031995, 608.0001599808, 637.000479961593, 
    639.00303964802, 731, 842.02784786653, 916.091492142188, 1050.5963405874, 
    1221.5325516491, 1367.77630871181,
  -3763.86345138056, -3640.39772426845, -3534.32039606405, -3271.09012173541, 
    -2962.04845284716, -2985.79530381883, -3066.7374540159, -2953.5353179653, 
    -2923.28098988581, -2952.75264338969, -2863.35452417633, 
    -2778.63033551535, -2746.85656954581, -2674.91982517127, 
    -2591.6564570073, -2559.42339071227, -2601.09683265301, 
    -2664.06225275186, -2675.34229994753, -2656.42684256247, 
    -2624.63509263441, -2563.78395128044, -2423.57617834088, 
    -2143.41982104701, -1499.79956803457, -1277.40198380927, 
    -1006.99984001792, -155.100047996159, -54.4000959807994, 
    217.001279699198, 633.001039916784, 977.990961075007, 1624.98808062121, 
    314.020318374089, 102.996480371176, 90.9978402559832, 182.000479961593, 
    791.971282892978, 1274.00735911041, 1273.98912087057, 609.004719692622, 
    821.011918912003, 819.998880089617, 700.0000799936, 705.000719923241, 
    627, 669.999520064002, 701, 765.000399967994, 733.000159974398, 
    590.000000006394, 808.467952036669, 890.279884578051, 1043.54815267953, 
    1209.78128897582, 1318.7555653446,
  -3714.0826057299, -3579.37901576364, -3421.48458083715, -3113.96297487135, 
    -2792.14447567085, -2828.0084786086, -3012.80113756122, 
    -3059.05617033024, -2983.00704334985, -2881.94101101085, 
    -2839.78392639135, -2789.02437065516, -2690.89702956553, 
    -2579.2120673481, -2504.30791520002, -2498.98421342107, 
    -2549.89015159972, -2609.356639828, -2631.77411332326, -2644.59868261642, 
    -2641.48694838309, -2556.87594358591, -2308.11799839496, 
    -1863.47122549394, -1545.1, -585.792928565733, -326.906551475865, -110.4, 
    32.0039996800183, 377.996560275187, 559, 1076.99248060157, 
    765.00655947523, 262, -59.5006319494429, -158.90004799616, 147, 
    1287.00439964802, 1681.99280057597, 1559, 1629.99176065916, 
    1316.98976081915, 1177, 287.999120070396, 702.999840012799, 622, 
    515.000239980801, 662.000639948803, 936, 938.003519718416, 
    617.999440044774, 816.371797062067, 888.949620919657, 1044.58038477611, 
    1191.95155911212, 1251.03033823289 ;

 alpha =
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, _, 
    _, _, _, _, _, _, _ ;

 f =
  7.27220521664304e-05, 7.27220521664304e-05, 7.27220521664304e-05, 
    7.27220521664304e-05, 7.27220521664304e-05, 7.27220521664304e-05, 
    7.27220521664304e-05, 7.27220521664304e-05, 7.27220521664304e-05, 
    7.27220521664304e-05, 7.27220521664304e-05, 7.27220521664304e-05, 
    7.27220521664304e-05, 7.27220521664304e-05, 7.27220521664304e-05, 
    7.27220521664304e-05, 7.27220521664304e-05, 7.27220521664304e-05, 
    7.27220521664304e-05, 7.27220521664304e-05, 7.27220521664304e-05, 
    7.27220521664304e-05, 7.27220521664304e-05, 7.27220521664304e-05, 
    7.27220521664304e-05, 7.27220521664304e-05, 7.27220521664304e-05, 
    7.27220521664304e-05, 7.27220521664304e-05, 7.27220521664304e-05, 
    7.27220521664304e-05, 7.27220521664304e-05, 7.27220521664304e-05, 
    7.27220521664304e-05, 7.27220521664304e-05, 7.27220521664304e-05, 
    7.27220521664304e-05, 7.27220521664304e-05, 7.27220521664304e-05, 
    7.27220521664304e-05, 7.27220521664304e-05, 7.27220521664304e-05, 
    7.27220521664304e-05, 7.27220521664304e-05, 7.27220521664304e-05, 
    7.27220521664304e-05, 7.27220521664304e-05, 7.27220521664304e-05, 
    7.27220521664304e-05, 7.27220521664304e-05, 7.27220521664304e-05, 
    7.27220521664304e-05, 7.27220521664304e-05, 7.27220521664304e-05, 
    7.27220521664304e-05, 7.27220521664304e-05,
  7.34536129691974e-05, 7.34536129691974e-05, 7.34536129691974e-05, 
    7.34536129691974e-05, 7.34536129691974e-05, 7.34536129691974e-05, 
    7.34536129691974e-05, 7.34536129691974e-05, 7.34536129691974e-05, 
    7.34536129691974e-05, 7.34536129691974e-05, 7.34536129691974e-05, 
    7.34536129691974e-05, 7.34536129691974e-05, 7.34536129691974e-05, 
    7.34536129691974e-05, 7.34536129691974e-05, 7.34536129691974e-05, 
    7.34536129691974e-05, 7.34536129691974e-05, 7.34536129691974e-05, 
    7.34536129691974e-05, 7.34536129691974e-05, 7.34536129691974e-05, 
    7.34536129691974e-05, 7.34536129691974e-05, 7.34536129691974e-05, 
    7.34536129691974e-05, 7.34536129691974e-05, 7.34536129691974e-05, 
    7.34536129691974e-05, 7.34536129691974e-05, 7.34536129691974e-05, 
    7.34536129691974e-05, 7.34536129691974e-05, 7.34536129691974e-05, 
    7.34536129691974e-05, 7.34536129691974e-05, 7.34536129691974e-05, 
    7.34536129691974e-05, 7.34536129691974e-05, 7.34536129691974e-05, 
    7.34536129691974e-05, 7.34536129691974e-05, 7.34536129691974e-05, 
    7.34536129691974e-05, 7.34536129691974e-05, 7.34536129691974e-05, 
    7.34536129691974e-05, 7.34536129691974e-05, 7.34536129691974e-05, 
    7.34536129691974e-05, 7.34536129691974e-05, 7.34536129691974e-05, 
    7.34536129691974e-05, 7.34536129691974e-05,
  7.41826876400814e-05, 7.41826876400814e-05, 7.41826876400814e-05, 
    7.41826876400814e-05, 7.41826876400814e-05, 7.41826876400814e-05, 
    7.41826876400814e-05, 7.41826876400814e-05, 7.41826876400814e-05, 
    7.41826876400814e-05, 7.41826876400814e-05, 7.41826876400814e-05, 
    7.41826876400814e-05, 7.41826876400814e-05, 7.41826876400814e-05, 
    7.41826876400814e-05, 7.41826876400814e-05, 7.41826876400814e-05, 
    7.41826876400814e-05, 7.41826876400814e-05, 7.41826876400814e-05, 
    7.41826876400814e-05, 7.41826876400814e-05, 7.41826876400814e-05, 
    7.41826876400814e-05, 7.41826876400814e-05, 7.41826876400814e-05, 
    7.41826876400814e-05, 7.41826876400814e-05, 7.41826876400814e-05, 
    7.41826876400814e-05, 7.41826876400814e-05, 7.41826876400814e-05, 
    7.41826876400814e-05, 7.41826876400814e-05, 7.41826876400814e-05, 
    7.41826876400814e-05, 7.41826876400814e-05, 7.41826876400814e-05, 
    7.41826876400814e-05, 7.41826876400814e-05, 7.41826876400814e-05, 
    7.41826876400814e-05, 7.41826876400814e-05, 7.41826876400814e-05, 
    7.41826876400814e-05, 7.41826876400814e-05, 7.41826876400814e-05, 
    7.41826876400814e-05, 7.41826876400814e-05, 7.41826876400814e-05, 
    7.41826876400814e-05, 7.41826876400814e-05, 7.41826876400814e-05, 
    7.41826876400814e-05, 7.41826876400814e-05,
  7.49092515026137e-05, 7.49092515026137e-05, 7.49092515026137e-05, 
    7.49092515026137e-05, 7.49092515026137e-05, 7.49092515026137e-05, 
    7.49092515026137e-05, 7.49092515026137e-05, 7.49092515026137e-05, 
    7.49092515026137e-05, 7.49092515026137e-05, 7.49092515026137e-05, 
    7.49092515026137e-05, 7.49092515026137e-05, 7.49092515026137e-05, 
    7.49092515026137e-05, 7.49092515026137e-05, 7.49092515026137e-05, 
    7.49092515026137e-05, 7.49092515026137e-05, 7.49092515026137e-05, 
    7.49092515026137e-05, 7.49092515026137e-05, 7.49092515026137e-05, 
    7.49092515026137e-05, 7.49092515026137e-05, 7.49092515026137e-05, 
    7.49092515026137e-05, 7.49092515026137e-05, 7.49092515026137e-05, 
    7.49092515026137e-05, 7.49092515026137e-05, 7.49092515026137e-05, 
    7.49092515026137e-05, 7.49092515026137e-05, 7.49092515026137e-05, 
    7.49092515026137e-05, 7.49092515026137e-05, 7.49092515026137e-05, 
    7.49092515026137e-05, 7.49092515026137e-05, 7.49092515026137e-05, 
    7.49092515026137e-05, 7.49092515026137e-05, 7.49092515026137e-05, 
    7.49092515026137e-05, 7.49092515026137e-05, 7.49092515026137e-05, 
    7.49092515026137e-05, 7.49092515026137e-05, 7.49092515026137e-05, 
    7.49092515026137e-05, 7.49092515026137e-05, 7.49092515026137e-05, 
    7.49092515026137e-05, 7.49092515026137e-05,
  7.56332799653071e-05, 7.56332799653071e-05, 7.56332799653071e-05, 
    7.56332799653071e-05, 7.56332799653071e-05, 7.56332799653071e-05, 
    7.56332799653071e-05, 7.56332799653071e-05, 7.56332799653071e-05, 
    7.56332799653071e-05, 7.56332799653071e-05, 7.56332799653071e-05, 
    7.56332799653071e-05, 7.56332799653071e-05, 7.56332799653071e-05, 
    7.56332799653071e-05, 7.56332799653071e-05, 7.56332799653071e-05, 
    7.56332799653071e-05, 7.56332799653071e-05, 7.56332799653071e-05, 
    7.56332799653071e-05, 7.56332799653071e-05, 7.56332799653071e-05, 
    7.56332799653071e-05, 7.56332799653071e-05, 7.56332799653071e-05, 
    7.56332799653071e-05, 7.56332799653071e-05, 7.56332799653071e-05, 
    7.56332799653071e-05, 7.56332799653071e-05, 7.56332799653071e-05, 
    7.56332799653071e-05, 7.56332799653071e-05, 7.56332799653071e-05, 
    7.56332799653071e-05, 7.56332799653071e-05, 7.56332799653071e-05, 
    7.56332799653071e-05, 7.56332799653071e-05, 7.56332799653071e-05, 
    7.56332799653071e-05, 7.56332799653071e-05, 7.56332799653071e-05, 
    7.56332799653071e-05, 7.56332799653071e-05, 7.56332799653071e-05, 
    7.56332799653071e-05, 7.56332799653071e-05, 7.56332799653071e-05, 
    7.56332799653071e-05, 7.56332799653071e-05, 7.56332799653071e-05, 
    7.56332799653071e-05, 7.56332799653071e-05,
  7.63547485224882e-05, 7.63547485224882e-05, 7.63547485224882e-05, 
    7.63547485224882e-05, 7.63547485224882e-05, 7.63547485224882e-05, 
    7.63547485224882e-05, 7.63547485224882e-05, 7.63547485224882e-05, 
    7.63547485224882e-05, 7.63547485224882e-05, 7.63547485224882e-05, 
    7.63547485224882e-05, 7.63547485224882e-05, 7.63547485224882e-05, 
    7.63547485224882e-05, 7.63547485224882e-05, 7.63547485224882e-05, 
    7.63547485224882e-05, 7.63547485224882e-05, 7.63547485224882e-05, 
    7.63547485224882e-05, 7.63547485224882e-05, 7.63547485224882e-05, 
    7.63547485224882e-05, 7.63547485224882e-05, 7.63547485224882e-05, 
    7.63547485224882e-05, 7.63547485224882e-05, 7.63547485224882e-05, 
    7.63547485224882e-05, 7.63547485224882e-05, 7.63547485224882e-05, 
    7.63547485224882e-05, 7.63547485224882e-05, 7.63547485224882e-05, 
    7.63547485224882e-05, 7.63547485224882e-05, 7.63547485224882e-05, 
    7.63547485224882e-05, 7.63547485224882e-05, 7.63547485224882e-05, 
    7.63547485224882e-05, 7.63547485224882e-05, 7.63547485224882e-05, 
    7.63547485224882e-05, 7.63547485224882e-05, 7.63547485224882e-05, 
    7.63547485224882e-05, 7.63547485224882e-05, 7.63547485224882e-05, 
    7.63547485224882e-05, 7.63547485224882e-05, 7.63547485224882e-05, 
    7.63547485224882e-05, 7.63547485224882e-05,
  7.70736327551271e-05, 7.70736327551271e-05, 7.70736327551271e-05, 
    7.70736327551271e-05, 7.70736327551271e-05, 7.70736327551271e-05, 
    7.70736327551271e-05, 7.70736327551271e-05, 7.70736327551271e-05, 
    7.70736327551271e-05, 7.70736327551271e-05, 7.70736327551271e-05, 
    7.70736327551271e-05, 7.70736327551271e-05, 7.70736327551271e-05, 
    7.70736327551271e-05, 7.70736327551271e-05, 7.70736327551271e-05, 
    7.70736327551271e-05, 7.70736327551271e-05, 7.70736327551271e-05, 
    7.70736327551271e-05, 7.70736327551271e-05, 7.70736327551271e-05, 
    7.70736327551271e-05, 7.70736327551271e-05, 7.70736327551271e-05, 
    7.70736327551271e-05, 7.70736327551271e-05, 7.70736327551271e-05, 
    7.70736327551271e-05, 7.70736327551271e-05, 7.70736327551271e-05, 
    7.70736327551271e-05, 7.70736327551271e-05, 7.70736327551271e-05, 
    7.70736327551271e-05, 7.70736327551271e-05, 7.70736327551271e-05, 
    7.70736327551271e-05, 7.70736327551271e-05, 7.70736327551271e-05, 
    7.70736327551271e-05, 7.70736327551271e-05, 7.70736327551271e-05, 
    7.70736327551271e-05, 7.70736327551271e-05, 7.70736327551271e-05, 
    7.70736327551271e-05, 7.70736327551271e-05, 7.70736327551271e-05, 
    7.70736327551271e-05, 7.70736327551271e-05, 7.70736327551271e-05, 
    7.70736327551271e-05, 7.70736327551271e-05,
  7.77899083316634e-05, 7.77899083316634e-05, 7.77899083316634e-05, 
    7.77899083316634e-05, 7.77899083316634e-05, 7.77899083316634e-05, 
    7.77899083316634e-05, 7.77899083316634e-05, 7.77899083316634e-05, 
    7.77899083316634e-05, 7.77899083316634e-05, 7.77899083316634e-05, 
    7.77899083316634e-05, 7.77899083316634e-05, 7.77899083316634e-05, 
    7.77899083316634e-05, 7.77899083316634e-05, 7.77899083316634e-05, 
    7.77899083316634e-05, 7.77899083316634e-05, 7.77899083316634e-05, 
    7.77899083316634e-05, 7.77899083316634e-05, 7.77899083316634e-05, 
    7.77899083316634e-05, 7.77899083316634e-05, 7.77899083316634e-05, 
    7.77899083316634e-05, 7.77899083316634e-05, 7.77899083316634e-05, 
    7.77899083316634e-05, 7.77899083316634e-05, 7.77899083316634e-05, 
    7.77899083316634e-05, 7.77899083316634e-05, 7.77899083316634e-05, 
    7.77899083316634e-05, 7.77899083316634e-05, 7.77899083316634e-05, 
    7.77899083316634e-05, 7.77899083316634e-05, 7.77899083316634e-05, 
    7.77899083316634e-05, 7.77899083316634e-05, 7.77899083316634e-05, 
    7.77899083316634e-05, 7.77899083316634e-05, 7.77899083316634e-05, 
    7.77899083316634e-05, 7.77899083316634e-05, 7.77899083316634e-05, 
    7.77899083316634e-05, 7.77899083316634e-05, 7.77899083316634e-05, 
    7.77899083316634e-05, 7.77899083316634e-05,
  7.85035510088301e-05, 7.85035510088301e-05, 7.85035510088301e-05, 
    7.85035510088301e-05, 7.85035510088301e-05, 7.85035510088301e-05, 
    7.85035510088301e-05, 7.85035510088301e-05, 7.85035510088301e-05, 
    7.85035510088301e-05, 7.85035510088301e-05, 7.85035510088301e-05, 
    7.85035510088301e-05, 7.85035510088301e-05, 7.85035510088301e-05, 
    7.85035510088301e-05, 7.85035510088301e-05, 7.85035510088301e-05, 
    7.85035510088301e-05, 7.85035510088301e-05, 7.85035510088301e-05, 
    7.85035510088301e-05, 7.85035510088301e-05, 7.85035510088301e-05, 
    7.85035510088301e-05, 7.85035510088301e-05, 7.85035510088301e-05, 
    7.85035510088301e-05, 7.85035510088301e-05, 7.85035510088301e-05, 
    7.85035510088301e-05, 7.85035510088301e-05, 7.85035510088301e-05, 
    7.85035510088301e-05, 7.85035510088301e-05, 7.85035510088301e-05, 
    7.85035510088301e-05, 7.85035510088301e-05, 7.85035510088301e-05, 
    7.85035510088301e-05, 7.85035510088301e-05, 7.85035510088301e-05, 
    7.85035510088301e-05, 7.85035510088301e-05, 7.85035510088301e-05, 
    7.85035510088301e-05, 7.85035510088301e-05, 7.85035510088301e-05, 
    7.85035510088301e-05, 7.85035510088301e-05, 7.85035510088301e-05, 
    7.85035510088301e-05, 7.85035510088301e-05, 7.85035510088301e-05, 
    7.85035510088301e-05, 7.85035510088301e-05,
  7.92145366324742e-05, 7.92145366324742e-05, 7.92145366324742e-05, 
    7.92145366324742e-05, 7.92145366324742e-05, 7.92145366324742e-05, 
    7.92145366324742e-05, 7.92145366324742e-05, 7.92145366324742e-05, 
    7.92145366324742e-05, 7.92145366324742e-05, 7.92145366324742e-05, 
    7.92145366324742e-05, 7.92145366324742e-05, 7.92145366324742e-05, 
    7.92145366324742e-05, 7.92145366324742e-05, 7.92145366324742e-05, 
    7.92145366324742e-05, 7.92145366324742e-05, 7.92145366324742e-05, 
    7.92145366324742e-05, 7.92145366324742e-05, 7.92145366324742e-05, 
    7.92145366324742e-05, 7.92145366324742e-05, 7.92145366324742e-05, 
    7.92145366324742e-05, 7.92145366324742e-05, 7.92145366324742e-05, 
    7.92145366324742e-05, 7.92145366324742e-05, 7.92145366324742e-05, 
    7.92145366324742e-05, 7.92145366324742e-05, 7.92145366324742e-05, 
    7.92145366324742e-05, 7.92145366324742e-05, 7.92145366324742e-05, 
    7.92145366324742e-05, 7.92145366324742e-05, 7.92145366324742e-05, 
    7.92145366324742e-05, 7.92145366324742e-05, 7.92145366324742e-05, 
    7.92145366324742e-05, 7.92145366324742e-05, 7.92145366324742e-05, 
    7.92145366324742e-05, 7.92145366324742e-05, 7.92145366324742e-05, 
    7.92145366324742e-05, 7.92145366324742e-05, 7.92145366324742e-05, 
    7.92145366324742e-05, 7.92145366324742e-05,
  7.9922841138374e-05, 7.9922841138374e-05, 7.9922841138374e-05, 
    7.9922841138374e-05, 7.9922841138374e-05, 7.9922841138374e-05, 
    7.9922841138374e-05, 7.9922841138374e-05, 7.9922841138374e-05, 
    7.9922841138374e-05, 7.9922841138374e-05, 7.9922841138374e-05, 
    7.9922841138374e-05, 7.9922841138374e-05, 7.9922841138374e-05, 
    7.9922841138374e-05, 7.9922841138374e-05, 7.9922841138374e-05, 
    7.9922841138374e-05, 7.9922841138374e-05, 7.9922841138374e-05, 
    7.9922841138374e-05, 7.9922841138374e-05, 7.9922841138374e-05, 
    7.9922841138374e-05, 7.9922841138374e-05, 7.9922841138374e-05, 
    7.9922841138374e-05, 7.9922841138374e-05, 7.9922841138374e-05, 
    7.9922841138374e-05, 7.9922841138374e-05, 7.9922841138374e-05, 
    7.9922841138374e-05, 7.9922841138374e-05, 7.9922841138374e-05, 
    7.9922841138374e-05, 7.9922841138374e-05, 7.9922841138374e-05, 
    7.9922841138374e-05, 7.9922841138374e-05, 7.9922841138374e-05, 
    7.9922841138374e-05, 7.9922841138374e-05, 7.9922841138374e-05, 
    7.9922841138374e-05, 7.9922841138374e-05, 7.9922841138374e-05, 
    7.9922841138374e-05, 7.9922841138374e-05, 7.9922841138374e-05, 
    7.9922841138374e-05, 7.9922841138374e-05, 7.9922841138374e-05, 
    7.9922841138374e-05, 7.9922841138374e-05,
  8.06284405530537e-05, 8.06284405530537e-05, 8.06284405530537e-05, 
    8.06284405530537e-05, 8.06284405530537e-05, 8.06284405530537e-05, 
    8.06284405530537e-05, 8.06284405530537e-05, 8.06284405530537e-05, 
    8.06284405530537e-05, 8.06284405530537e-05, 8.06284405530537e-05, 
    8.06284405530537e-05, 8.06284405530537e-05, 8.06284405530537e-05, 
    8.06284405530537e-05, 8.06284405530537e-05, 8.06284405530537e-05, 
    8.06284405530537e-05, 8.06284405530537e-05, 8.06284405530537e-05, 
    8.06284405530537e-05, 8.06284405530537e-05, 8.06284405530537e-05, 
    8.06284405530537e-05, 8.06284405530537e-05, 8.06284405530537e-05, 
    8.06284405530537e-05, 8.06284405530537e-05, 8.06284405530537e-05, 
    8.06284405530537e-05, 8.06284405530537e-05, 8.06284405530537e-05, 
    8.06284405530537e-05, 8.06284405530537e-05, 8.06284405530537e-05, 
    8.06284405530537e-05, 8.06284405530537e-05, 8.06284405530537e-05, 
    8.06284405530537e-05, 8.06284405530537e-05, 8.06284405530537e-05, 
    8.06284405530537e-05, 8.06284405530537e-05, 8.06284405530537e-05, 
    8.06284405530537e-05, 8.06284405530537e-05, 8.06284405530537e-05, 
    8.06284405530537e-05, 8.06284405530537e-05, 8.06284405530537e-05, 
    8.06284405530537e-05, 8.06284405530537e-05, 8.06284405530537e-05, 
    8.06284405530537e-05, 8.06284405530537e-05,
  8.13313109945947e-05, 8.13313109945947e-05, 8.13313109945947e-05, 
    8.13313109945947e-05, 8.13313109945947e-05, 8.13313109945947e-05, 
    8.13313109945947e-05, 8.13313109945947e-05, 8.13313109945947e-05, 
    8.13313109945947e-05, 8.13313109945947e-05, 8.13313109945947e-05, 
    8.13313109945947e-05, 8.13313109945947e-05, 8.13313109945947e-05, 
    8.13313109945947e-05, 8.13313109945947e-05, 8.13313109945947e-05, 
    8.13313109945947e-05, 8.13313109945947e-05, 8.13313109945947e-05, 
    8.13313109945947e-05, 8.13313109945947e-05, 8.13313109945947e-05, 
    8.13313109945947e-05, 8.13313109945947e-05, 8.13313109945947e-05, 
    8.13313109945947e-05, 8.13313109945947e-05, 8.13313109945947e-05, 
    8.13313109945947e-05, 8.13313109945947e-05, 8.13313109945947e-05, 
    8.13313109945947e-05, 8.13313109945947e-05, 8.13313109945947e-05, 
    8.13313109945947e-05, 8.13313109945947e-05, 8.13313109945947e-05, 
    8.13313109945947e-05, 8.13313109945947e-05, 8.13313109945947e-05, 
    8.13313109945947e-05, 8.13313109945947e-05, 8.13313109945947e-05, 
    8.13313109945947e-05, 8.13313109945947e-05, 8.13313109945947e-05, 
    8.13313109945947e-05, 8.13313109945947e-05, 8.13313109945947e-05, 
    8.13313109945947e-05, 8.13313109945947e-05, 8.13313109945947e-05, 
    8.13313109945947e-05, 8.13313109945947e-05,
  8.2031428673444e-05, 8.2031428673444e-05, 8.2031428673444e-05, 
    8.2031428673444e-05, 8.2031428673444e-05, 8.2031428673444e-05, 
    8.2031428673444e-05, 8.2031428673444e-05, 8.2031428673444e-05, 
    8.2031428673444e-05, 8.2031428673444e-05, 8.2031428673444e-05, 
    8.2031428673444e-05, 8.2031428673444e-05, 8.2031428673444e-05, 
    8.2031428673444e-05, 8.2031428673444e-05, 8.2031428673444e-05, 
    8.2031428673444e-05, 8.2031428673444e-05, 8.2031428673444e-05, 
    8.2031428673444e-05, 8.2031428673444e-05, 8.2031428673444e-05, 
    8.2031428673444e-05, 8.2031428673444e-05, 8.2031428673444e-05, 
    8.2031428673444e-05, 8.2031428673444e-05, 8.2031428673444e-05, 
    8.2031428673444e-05, 8.2031428673444e-05, 8.2031428673444e-05, 
    8.2031428673444e-05, 8.2031428673444e-05, 8.2031428673444e-05, 
    8.2031428673444e-05, 8.2031428673444e-05, 8.2031428673444e-05, 
    8.2031428673444e-05, 8.2031428673444e-05, 8.2031428673444e-05, 
    8.2031428673444e-05, 8.2031428673444e-05, 8.2031428673444e-05, 
    8.2031428673444e-05, 8.2031428673444e-05, 8.2031428673444e-05, 
    8.2031428673444e-05, 8.2031428673444e-05, 8.2031428673444e-05, 
    8.2031428673444e-05, 8.2031428673444e-05, 8.2031428673444e-05, 
    8.2031428673444e-05, 8.2031428673444e-05,
  8.27287698932196e-05, 8.27287698932196e-05, 8.27287698932196e-05, 
    8.27287698932196e-05, 8.27287698932196e-05, 8.27287698932196e-05, 
    8.27287698932196e-05, 8.27287698932196e-05, 8.27287698932196e-05, 
    8.27287698932196e-05, 8.27287698932196e-05, 8.27287698932196e-05, 
    8.27287698932196e-05, 8.27287698932196e-05, 8.27287698932196e-05, 
    8.27287698932196e-05, 8.27287698932196e-05, 8.27287698932196e-05, 
    8.27287698932196e-05, 8.27287698932196e-05, 8.27287698932196e-05, 
    8.27287698932196e-05, 8.27287698932196e-05, 8.27287698932196e-05, 
    8.27287698932196e-05, 8.27287698932196e-05, 8.27287698932196e-05, 
    8.27287698932196e-05, 8.27287698932196e-05, 8.27287698932196e-05, 
    8.27287698932196e-05, 8.27287698932196e-05, 8.27287698932196e-05, 
    8.27287698932196e-05, 8.27287698932196e-05, 8.27287698932196e-05, 
    8.27287698932196e-05, 8.27287698932196e-05, 8.27287698932196e-05, 
    8.27287698932196e-05, 8.27287698932196e-05, 8.27287698932196e-05, 
    8.27287698932196e-05, 8.27287698932196e-05, 8.27287698932196e-05, 
    8.27287698932196e-05, 8.27287698932196e-05, 8.27287698932196e-05, 
    8.27287698932196e-05, 8.27287698932196e-05, 8.27287698932196e-05, 
    8.27287698932196e-05, 8.27287698932196e-05, 8.27287698932196e-05, 
    8.27287698932196e-05, 8.27287698932196e-05,
  8.3423311051512e-05, 8.3423311051512e-05, 8.3423311051512e-05, 
    8.3423311051512e-05, 8.3423311051512e-05, 8.3423311051512e-05, 
    8.3423311051512e-05, 8.3423311051512e-05, 8.3423311051512e-05, 
    8.3423311051512e-05, 8.3423311051512e-05, 8.3423311051512e-05, 
    8.3423311051512e-05, 8.3423311051512e-05, 8.3423311051512e-05, 
    8.3423311051512e-05, 8.3423311051512e-05, 8.3423311051512e-05, 
    8.3423311051512e-05, 8.3423311051512e-05, 8.3423311051512e-05, 
    8.3423311051512e-05, 8.3423311051512e-05, 8.3423311051512e-05, 
    8.3423311051512e-05, 8.3423311051512e-05, 8.3423311051512e-05, 
    8.3423311051512e-05, 8.3423311051512e-05, 8.3423311051512e-05, 
    8.3423311051512e-05, 8.3423311051512e-05, 8.3423311051512e-05, 
    8.3423311051512e-05, 8.3423311051512e-05, 8.3423311051512e-05, 
    8.3423311051512e-05, 8.3423311051512e-05, 8.3423311051512e-05, 
    8.3423311051512e-05, 8.3423311051512e-05, 8.3423311051512e-05, 
    8.3423311051512e-05, 8.3423311051512e-05, 8.3423311051512e-05, 
    8.3423311051512e-05, 8.3423311051512e-05, 8.3423311051512e-05, 
    8.3423311051512e-05, 8.3423311051512e-05, 8.3423311051512e-05, 
    8.3423311051512e-05, 8.3423311051512e-05, 8.3423311051512e-05, 
    8.3423311051512e-05, 8.3423311051512e-05,
  8.41150286406838e-05, 8.41150286406838e-05, 8.41150286406838e-05, 
    8.41150286406838e-05, 8.41150286406838e-05, 8.41150286406838e-05, 
    8.41150286406838e-05, 8.41150286406838e-05, 8.41150286406838e-05, 
    8.41150286406838e-05, 8.41150286406838e-05, 8.41150286406838e-05, 
    8.41150286406838e-05, 8.41150286406838e-05, 8.41150286406838e-05, 
    8.41150286406838e-05, 8.41150286406838e-05, 8.41150286406838e-05, 
    8.41150286406838e-05, 8.41150286406838e-05, 8.41150286406838e-05, 
    8.41150286406838e-05, 8.41150286406838e-05, 8.41150286406838e-05, 
    8.41150286406838e-05, 8.41150286406838e-05, 8.41150286406838e-05, 
    8.41150286406838e-05, 8.41150286406838e-05, 8.41150286406838e-05, 
    8.41150286406838e-05, 8.41150286406838e-05, 8.41150286406838e-05, 
    8.41150286406838e-05, 8.41150286406838e-05, 8.41150286406838e-05, 
    8.41150286406838e-05, 8.41150286406838e-05, 8.41150286406838e-05, 
    8.41150286406838e-05, 8.41150286406838e-05, 8.41150286406838e-05, 
    8.41150286406838e-05, 8.41150286406838e-05, 8.41150286406838e-05, 
    8.41150286406838e-05, 8.41150286406838e-05, 8.41150286406838e-05, 
    8.41150286406838e-05, 8.41150286406838e-05, 8.41150286406838e-05, 
    8.41150286406838e-05, 8.41150286406838e-05, 8.41150286406838e-05, 
    8.41150286406838e-05, 8.41150286406838e-05,
  8.48038992486644e-05, 8.48038992486644e-05, 8.48038992486644e-05, 
    8.48038992486644e-05, 8.48038992486644e-05, 8.48038992486644e-05, 
    8.48038992486644e-05, 8.48038992486644e-05, 8.48038992486644e-05, 
    8.48038992486644e-05, 8.48038992486644e-05, 8.48038992486644e-05, 
    8.48038992486644e-05, 8.48038992486644e-05, 8.48038992486644e-05, 
    8.48038992486644e-05, 8.48038992486644e-05, 8.48038992486644e-05, 
    8.48038992486644e-05, 8.48038992486644e-05, 8.48038992486644e-05, 
    8.48038992486644e-05, 8.48038992486644e-05, 8.48038992486644e-05, 
    8.48038992486644e-05, 8.48038992486644e-05, 8.48038992486644e-05, 
    8.48038992486644e-05, 8.48038992486644e-05, 8.48038992486644e-05, 
    8.48038992486644e-05, 8.48038992486644e-05, 8.48038992486644e-05, 
    8.48038992486644e-05, 8.48038992486644e-05, 8.48038992486644e-05, 
    8.48038992486644e-05, 8.48038992486644e-05, 8.48038992486644e-05, 
    8.48038992486644e-05, 8.48038992486644e-05, 8.48038992486644e-05, 
    8.48038992486644e-05, 8.48038992486644e-05, 8.48038992486644e-05, 
    8.48038992486644e-05, 8.48038992486644e-05, 8.48038992486644e-05, 
    8.48038992486644e-05, 8.48038992486644e-05, 8.48038992486644e-05, 
    8.48038992486644e-05, 8.48038992486644e-05, 8.48038992486644e-05, 
    8.48038992486644e-05, 8.48038992486644e-05,
  8.54898995597434e-05, 8.54898995597434e-05, 8.54898995597434e-05, 
    8.54898995597434e-05, 8.54898995597434e-05, 8.54898995597434e-05, 
    8.54898995597434e-05, 8.54898995597434e-05, 8.54898995597434e-05, 
    8.54898995597434e-05, 8.54898995597434e-05, 8.54898995597434e-05, 
    8.54898995597434e-05, 8.54898995597434e-05, 8.54898995597434e-05, 
    8.54898995597434e-05, 8.54898995597434e-05, 8.54898995597434e-05, 
    8.54898995597434e-05, 8.54898995597434e-05, 8.54898995597434e-05, 
    8.54898995597434e-05, 8.54898995597434e-05, 8.54898995597434e-05, 
    8.54898995597434e-05, 8.54898995597434e-05, 8.54898995597434e-05, 
    8.54898995597434e-05, 8.54898995597434e-05, 8.54898995597434e-05, 
    8.54898995597434e-05, 8.54898995597434e-05, 8.54898995597434e-05, 
    8.54898995597434e-05, 8.54898995597434e-05, 8.54898995597434e-05, 
    8.54898995597434e-05, 8.54898995597434e-05, 8.54898995597434e-05, 
    8.54898995597434e-05, 8.54898995597434e-05, 8.54898995597434e-05, 
    8.54898995597434e-05, 8.54898995597434e-05, 8.54898995597434e-05, 
    8.54898995597434e-05, 8.54898995597434e-05, 8.54898995597434e-05, 
    8.54898995597434e-05, 8.54898995597434e-05, 8.54898995597434e-05, 
    8.54898995597434e-05, 8.54898995597434e-05, 8.54898995597434e-05, 
    8.54898995597434e-05, 8.54898995597434e-05,
  8.6173006355359e-05, 8.6173006355359e-05, 8.6173006355359e-05, 
    8.6173006355359e-05, 8.6173006355359e-05, 8.6173006355359e-05, 
    8.6173006355359e-05, 8.6173006355359e-05, 8.6173006355359e-05, 
    8.6173006355359e-05, 8.6173006355359e-05, 8.6173006355359e-05, 
    8.6173006355359e-05, 8.6173006355359e-05, 8.6173006355359e-05, 
    8.6173006355359e-05, 8.6173006355359e-05, 8.6173006355359e-05, 
    8.6173006355359e-05, 8.6173006355359e-05, 8.6173006355359e-05, 
    8.6173006355359e-05, 8.6173006355359e-05, 8.6173006355359e-05, 
    8.6173006355359e-05, 8.6173006355359e-05, 8.6173006355359e-05, 
    8.6173006355359e-05, 8.6173006355359e-05, 8.6173006355359e-05, 
    8.6173006355359e-05, 8.6173006355359e-05, 8.6173006355359e-05, 
    8.6173006355359e-05, 8.6173006355359e-05, 8.6173006355359e-05, 
    8.6173006355359e-05, 8.6173006355359e-05, 8.6173006355359e-05, 
    8.6173006355359e-05, 8.6173006355359e-05, 8.6173006355359e-05, 
    8.6173006355359e-05, 8.6173006355359e-05, 8.6173006355359e-05, 
    8.6173006355359e-05, 8.6173006355359e-05, 8.6173006355359e-05, 
    8.6173006355359e-05, 8.6173006355359e-05, 8.6173006355359e-05, 
    8.6173006355359e-05, 8.6173006355359e-05, 8.6173006355359e-05, 
    8.6173006355359e-05, 8.6173006355359e-05,
  8.68531965148842e-05, 8.68531965148842e-05, 8.68531965148842e-05, 
    8.68531965148842e-05, 8.68531965148842e-05, 8.68531965148842e-05, 
    8.68531965148842e-05, 8.68531965148842e-05, 8.68531965148842e-05, 
    8.68531965148842e-05, 8.68531965148842e-05, 8.68531965148842e-05, 
    8.68531965148842e-05, 8.68531965148842e-05, 8.68531965148842e-05, 
    8.68531965148842e-05, 8.68531965148842e-05, 8.68531965148842e-05, 
    8.68531965148842e-05, 8.68531965148842e-05, 8.68531965148842e-05, 
    8.68531965148842e-05, 8.68531965148842e-05, 8.68531965148842e-05, 
    8.68531965148842e-05, 8.68531965148842e-05, 8.68531965148842e-05, 
    8.68531965148842e-05, 8.68531965148842e-05, 8.68531965148842e-05, 
    8.68531965148842e-05, 8.68531965148842e-05, 8.68531965148842e-05, 
    8.68531965148842e-05, 8.68531965148842e-05, 8.68531965148842e-05, 
    8.68531965148842e-05, 8.68531965148842e-05, 8.68531965148842e-05, 
    8.68531965148842e-05, 8.68531965148842e-05, 8.68531965148842e-05, 
    8.68531965148842e-05, 8.68531965148842e-05, 8.68531965148842e-05, 
    8.68531965148842e-05, 8.68531965148842e-05, 8.68531965148842e-05, 
    8.68531965148842e-05, 8.68531965148842e-05, 8.68531965148842e-05, 
    8.68531965148842e-05, 8.68531965148842e-05, 8.68531965148842e-05, 
    8.68531965148842e-05, 8.68531965148842e-05,
  8.75304470164095e-05, 8.75304470164095e-05, 8.75304470164095e-05, 
    8.75304470164095e-05, 8.75304470164095e-05, 8.75304470164095e-05, 
    8.75304470164095e-05, 8.75304470164095e-05, 8.75304470164095e-05, 
    8.75304470164095e-05, 8.75304470164095e-05, 8.75304470164095e-05, 
    8.75304470164095e-05, 8.75304470164095e-05, 8.75304470164095e-05, 
    8.75304470164095e-05, 8.75304470164095e-05, 8.75304470164095e-05, 
    8.75304470164095e-05, 8.75304470164095e-05, 8.75304470164095e-05, 
    8.75304470164095e-05, 8.75304470164095e-05, 8.75304470164095e-05, 
    8.75304470164095e-05, 8.75304470164095e-05, 8.75304470164095e-05, 
    8.75304470164095e-05, 8.75304470164095e-05, 8.75304470164095e-05, 
    8.75304470164095e-05, 8.75304470164095e-05, 8.75304470164095e-05, 
    8.75304470164095e-05, 8.75304470164095e-05, 8.75304470164095e-05, 
    8.75304470164095e-05, 8.75304470164095e-05, 8.75304470164095e-05, 
    8.75304470164095e-05, 8.75304470164095e-05, 8.75304470164095e-05, 
    8.75304470164095e-05, 8.75304470164095e-05, 8.75304470164095e-05, 
    8.75304470164095e-05, 8.75304470164095e-05, 8.75304470164095e-05, 
    8.75304470164095e-05, 8.75304470164095e-05, 8.75304470164095e-05, 
    8.75304470164095e-05, 8.75304470164095e-05, 8.75304470164095e-05, 
    8.75304470164095e-05, 8.75304470164095e-05,
  8.82047349375217e-05, 8.82047349375217e-05, 8.82047349375217e-05, 
    8.82047349375217e-05, 8.82047349375217e-05, 8.82047349375217e-05, 
    8.82047349375217e-05, 8.82047349375217e-05, 8.82047349375217e-05, 
    8.82047349375217e-05, 8.82047349375217e-05, 8.82047349375217e-05, 
    8.82047349375217e-05, 8.82047349375217e-05, 8.82047349375217e-05, 
    8.82047349375217e-05, 8.82047349375217e-05, 8.82047349375217e-05, 
    8.82047349375217e-05, 8.82047349375217e-05, 8.82047349375217e-05, 
    8.82047349375217e-05, 8.82047349375217e-05, 8.82047349375217e-05, 
    8.82047349375217e-05, 8.82047349375217e-05, 8.82047349375217e-05, 
    8.82047349375217e-05, 8.82047349375217e-05, 8.82047349375217e-05, 
    8.82047349375217e-05, 8.82047349375217e-05, 8.82047349375217e-05, 
    8.82047349375217e-05, 8.82047349375217e-05, 8.82047349375217e-05, 
    8.82047349375217e-05, 8.82047349375217e-05, 8.82047349375217e-05, 
    8.82047349375217e-05, 8.82047349375217e-05, 8.82047349375217e-05, 
    8.82047349375217e-05, 8.82047349375217e-05, 8.82047349375217e-05, 
    8.82047349375217e-05, 8.82047349375217e-05, 8.82047349375217e-05, 
    8.82047349375217e-05, 8.82047349375217e-05, 8.82047349375217e-05, 
    8.82047349375217e-05, 8.82047349375217e-05, 8.82047349375217e-05, 
    8.82047349375217e-05, 8.82047349375217e-05,
  8.88760374560798e-05, 8.88760374560798e-05, 8.88760374560798e-05, 
    8.88760374560798e-05, 8.88760374560798e-05, 8.88760374560798e-05, 
    8.88760374560798e-05, 8.88760374560798e-05, 8.88760374560798e-05, 
    8.88760374560798e-05, 8.88760374560798e-05, 8.88760374560798e-05, 
    8.88760374560798e-05, 8.88760374560798e-05, 8.88760374560798e-05, 
    8.88760374560798e-05, 8.88760374560798e-05, 8.88760374560798e-05, 
    8.88760374560798e-05, 8.88760374560798e-05, 8.88760374560798e-05, 
    8.88760374560798e-05, 8.88760374560798e-05, 8.88760374560798e-05, 
    8.88760374560798e-05, 8.88760374560798e-05, 8.88760374560798e-05, 
    8.88760374560798e-05, 8.88760374560798e-05, 8.88760374560798e-05, 
    8.88760374560798e-05, 8.88760374560798e-05, 8.88760374560798e-05, 
    8.88760374560798e-05, 8.88760374560798e-05, 8.88760374560798e-05, 
    8.88760374560798e-05, 8.88760374560798e-05, 8.88760374560798e-05, 
    8.88760374560798e-05, 8.88760374560798e-05, 8.88760374560798e-05, 
    8.88760374560798e-05, 8.88760374560798e-05, 8.88760374560798e-05, 
    8.88760374560798e-05, 8.88760374560798e-05, 8.88760374560798e-05, 
    8.88760374560798e-05, 8.88760374560798e-05, 8.88760374560798e-05, 
    8.88760374560798e-05, 8.88760374560798e-05, 8.88760374560798e-05, 
    8.88760374560798e-05, 8.88760374560798e-05,
  8.9544331850988e-05, 8.9544331850988e-05, 8.9544331850988e-05, 
    8.9544331850988e-05, 8.9544331850988e-05, 8.9544331850988e-05, 
    8.9544331850988e-05, 8.9544331850988e-05, 8.9544331850988e-05, 
    8.9544331850988e-05, 8.9544331850988e-05, 8.9544331850988e-05, 
    8.9544331850988e-05, 8.9544331850988e-05, 8.9544331850988e-05, 
    8.9544331850988e-05, 8.9544331850988e-05, 8.9544331850988e-05, 
    8.9544331850988e-05, 8.9544331850988e-05, 8.9544331850988e-05, 
    8.9544331850988e-05, 8.9544331850988e-05, 8.9544331850988e-05, 
    8.9544331850988e-05, 8.9544331850988e-05, 8.9544331850988e-05, 
    8.9544331850988e-05, 8.9544331850988e-05, 8.9544331850988e-05, 
    8.9544331850988e-05, 8.9544331850988e-05, 8.9544331850988e-05, 
    8.9544331850988e-05, 8.9544331850988e-05, 8.9544331850988e-05, 
    8.9544331850988e-05, 8.9544331850988e-05, 8.9544331850988e-05, 
    8.9544331850988e-05, 8.9544331850988e-05, 8.9544331850988e-05, 
    8.9544331850988e-05, 8.9544331850988e-05, 8.9544331850988e-05, 
    8.9544331850988e-05, 8.9544331850988e-05, 8.9544331850988e-05, 
    8.9544331850988e-05, 8.9544331850988e-05, 8.9544331850988e-05, 
    8.9544331850988e-05, 8.9544331850988e-05, 8.9544331850988e-05, 
    8.9544331850988e-05, 8.9544331850988e-05,
  9.0209595502964e-05, 9.0209595502964e-05, 9.0209595502964e-05, 
    9.0209595502964e-05, 9.0209595502964e-05, 9.0209595502964e-05, 
    9.0209595502964e-05, 9.0209595502964e-05, 9.0209595502964e-05, 
    9.0209595502964e-05, 9.0209595502964e-05, 9.0209595502964e-05, 
    9.0209595502964e-05, 9.0209595502964e-05, 9.0209595502964e-05, 
    9.0209595502964e-05, 9.0209595502964e-05, 9.0209595502964e-05, 
    9.0209595502964e-05, 9.0209595502964e-05, 9.0209595502964e-05, 
    9.0209595502964e-05, 9.0209595502964e-05, 9.0209595502964e-05, 
    9.0209595502964e-05, 9.0209595502964e-05, 9.0209595502964e-05, 
    9.0209595502964e-05, 9.0209595502964e-05, 9.0209595502964e-05, 
    9.0209595502964e-05, 9.0209595502964e-05, 9.0209595502964e-05, 
    9.0209595502964e-05, 9.0209595502964e-05, 9.0209595502964e-05, 
    9.0209595502964e-05, 9.0209595502964e-05, 9.0209595502964e-05, 
    9.0209595502964e-05, 9.0209595502964e-05, 9.0209595502964e-05, 
    9.0209595502964e-05, 9.0209595502964e-05, 9.0209595502964e-05, 
    9.0209595502964e-05, 9.0209595502964e-05, 9.0209595502964e-05, 
    9.0209595502964e-05, 9.0209595502964e-05, 9.0209595502964e-05, 
    9.0209595502964e-05, 9.0209595502964e-05, 9.0209595502964e-05, 
    9.0209595502964e-05, 9.0209595502964e-05,
  9.08718058953048e-05, 9.08718058953048e-05, 9.08718058953048e-05, 
    9.08718058953048e-05, 9.08718058953048e-05, 9.08718058953048e-05, 
    9.08718058953048e-05, 9.08718058953048e-05, 9.08718058953048e-05, 
    9.08718058953048e-05, 9.08718058953048e-05, 9.08718058953048e-05, 
    9.08718058953048e-05, 9.08718058953048e-05, 9.08718058953048e-05, 
    9.08718058953048e-05, 9.08718058953048e-05, 9.08718058953048e-05, 
    9.08718058953048e-05, 9.08718058953048e-05, 9.08718058953048e-05, 
    9.08718058953048e-05, 9.08718058953048e-05, 9.08718058953048e-05, 
    9.08718058953048e-05, 9.08718058953048e-05, 9.08718058953048e-05, 
    9.08718058953048e-05, 9.08718058953048e-05, 9.08718058953048e-05, 
    9.08718058953048e-05, 9.08718058953048e-05, 9.08718058953048e-05, 
    9.08718058953048e-05, 9.08718058953048e-05, 9.08718058953048e-05, 
    9.08718058953048e-05, 9.08718058953048e-05, 9.08718058953048e-05, 
    9.08718058953048e-05, 9.08718058953048e-05, 9.08718058953048e-05, 
    9.08718058953048e-05, 9.08718058953048e-05, 9.08718058953048e-05, 
    9.08718058953048e-05, 9.08718058953048e-05, 9.08718058953048e-05, 
    9.08718058953048e-05, 9.08718058953048e-05, 9.08718058953048e-05, 
    9.08718058953048e-05, 9.08718058953048e-05, 9.08718058953048e-05, 
    9.08718058953048e-05, 9.08718058953048e-05,
  9.15309406146493e-05, 9.15309406146493e-05, 9.15309406146493e-05, 
    9.15309406146493e-05, 9.15309406146493e-05, 9.15309406146493e-05, 
    9.15309406146493e-05, 9.15309406146493e-05, 9.15309406146493e-05, 
    9.15309406146493e-05, 9.15309406146493e-05, 9.15309406146493e-05, 
    9.15309406146493e-05, 9.15309406146493e-05, 9.15309406146493e-05, 
    9.15309406146493e-05, 9.15309406146493e-05, 9.15309406146493e-05, 
    9.15309406146493e-05, 9.15309406146493e-05, 9.15309406146493e-05, 
    9.15309406146493e-05, 9.15309406146493e-05, 9.15309406146493e-05, 
    9.15309406146493e-05, 9.15309406146493e-05, 9.15309406146493e-05, 
    9.15309406146493e-05, 9.15309406146493e-05, 9.15309406146493e-05, 
    9.15309406146493e-05, 9.15309406146493e-05, 9.15309406146493e-05, 
    9.15309406146493e-05, 9.15309406146493e-05, 9.15309406146493e-05, 
    9.15309406146493e-05, 9.15309406146493e-05, 9.15309406146493e-05, 
    9.15309406146493e-05, 9.15309406146493e-05, 9.15309406146493e-05, 
    9.15309406146493e-05, 9.15309406146493e-05, 9.15309406146493e-05, 
    9.15309406146493e-05, 9.15309406146493e-05, 9.15309406146493e-05, 
    9.15309406146493e-05, 9.15309406146493e-05, 9.15309406146493e-05, 
    9.15309406146493e-05, 9.15309406146493e-05, 9.15309406146493e-05, 
    9.15309406146493e-05, 9.15309406146493e-05,
  9.21869773517361e-05, 9.21869773517361e-05, 9.21869773517361e-05, 
    9.21869773517361e-05, 9.21869773517361e-05, 9.21869773517361e-05, 
    9.21869773517361e-05, 9.21869773517361e-05, 9.21869773517361e-05, 
    9.21869773517361e-05, 9.21869773517361e-05, 9.21869773517361e-05, 
    9.21869773517361e-05, 9.21869773517361e-05, 9.21869773517361e-05, 
    9.21869773517361e-05, 9.21869773517361e-05, 9.21869773517361e-05, 
    9.21869773517361e-05, 9.21869773517361e-05, 9.21869773517361e-05, 
    9.21869773517361e-05, 9.21869773517361e-05, 9.21869773517361e-05, 
    9.21869773517361e-05, 9.21869773517361e-05, 9.21869773517361e-05, 
    9.21869773517361e-05, 9.21869773517361e-05, 9.21869773517361e-05, 
    9.21869773517361e-05, 9.21869773517361e-05, 9.21869773517361e-05, 
    9.21869773517361e-05, 9.21869773517361e-05, 9.21869773517361e-05, 
    9.21869773517361e-05, 9.21869773517361e-05, 9.21869773517361e-05, 
    9.21869773517361e-05, 9.21869773517361e-05, 9.21869773517361e-05, 
    9.21869773517361e-05, 9.21869773517361e-05, 9.21869773517361e-05, 
    9.21869773517361e-05, 9.21869773517361e-05, 9.21869773517361e-05, 
    9.21869773517361e-05, 9.21869773517361e-05, 9.21869773517361e-05, 
    9.21869773517361e-05, 9.21869773517361e-05, 9.21869773517361e-05, 
    9.21869773517361e-05, 9.21869773517361e-05,
  9.28398939021592e-05, 9.28398939021592e-05, 9.28398939021592e-05, 
    9.28398939021592e-05, 9.28398939021592e-05, 9.28398939021592e-05, 
    9.28398939021592e-05, 9.28398939021592e-05, 9.28398939021592e-05, 
    9.28398939021592e-05, 9.28398939021592e-05, 9.28398939021592e-05, 
    9.28398939021592e-05, 9.28398939021592e-05, 9.28398939021592e-05, 
    9.28398939021592e-05, 9.28398939021592e-05, 9.28398939021592e-05, 
    9.28398939021592e-05, 9.28398939021592e-05, 9.28398939021592e-05, 
    9.28398939021592e-05, 9.28398939021592e-05, 9.28398939021592e-05, 
    9.28398939021592e-05, 9.28398939021592e-05, 9.28398939021592e-05, 
    9.28398939021592e-05, 9.28398939021592e-05, 9.28398939021592e-05, 
    9.28398939021592e-05, 9.28398939021592e-05, 9.28398939021592e-05, 
    9.28398939021592e-05, 9.28398939021592e-05, 9.28398939021592e-05, 
    9.28398939021592e-05, 9.28398939021592e-05, 9.28398939021592e-05, 
    9.28398939021592e-05, 9.28398939021592e-05, 9.28398939021592e-05, 
    9.28398939021592e-05, 9.28398939021592e-05, 9.28398939021592e-05, 
    9.28398939021592e-05, 9.28398939021592e-05, 9.28398939021592e-05, 
    9.28398939021592e-05, 9.28398939021592e-05, 9.28398939021592e-05, 
    9.28398939021592e-05, 9.28398939021592e-05, 9.28398939021592e-05, 
    9.28398939021592e-05, 9.28398939021592e-05,
  9.34896681671192e-05, 9.34896681671192e-05, 9.34896681671192e-05, 
    9.34896681671192e-05, 9.34896681671192e-05, 9.34896681671192e-05, 
    9.34896681671192e-05, 9.34896681671192e-05, 9.34896681671192e-05, 
    9.34896681671192e-05, 9.34896681671192e-05, 9.34896681671192e-05, 
    9.34896681671192e-05, 9.34896681671192e-05, 9.34896681671192e-05, 
    9.34896681671192e-05, 9.34896681671192e-05, 9.34896681671192e-05, 
    9.34896681671192e-05, 9.34896681671192e-05, 9.34896681671192e-05, 
    9.34896681671192e-05, 9.34896681671192e-05, 9.34896681671192e-05, 
    9.34896681671192e-05, 9.34896681671192e-05, 9.34896681671192e-05, 
    9.34896681671192e-05, 9.34896681671192e-05, 9.34896681671192e-05, 
    9.34896681671192e-05, 9.34896681671192e-05, 9.34896681671192e-05, 
    9.34896681671192e-05, 9.34896681671192e-05, 9.34896681671192e-05, 
    9.34896681671192e-05, 9.34896681671192e-05, 9.34896681671192e-05, 
    9.34896681671192e-05, 9.34896681671192e-05, 9.34896681671192e-05, 
    9.34896681671192e-05, 9.34896681671192e-05, 9.34896681671192e-05, 
    9.34896681671192e-05, 9.34896681671192e-05, 9.34896681671192e-05, 
    9.34896681671192e-05, 9.34896681671192e-05, 9.34896681671192e-05, 
    9.34896681671192e-05, 9.34896681671192e-05, 9.34896681671192e-05, 
    9.34896681671192e-05, 9.34896681671192e-05,
  9.41362781541716e-05, 9.41362781541716e-05, 9.41362781541716e-05, 
    9.41362781541716e-05, 9.41362781541716e-05, 9.41362781541716e-05, 
    9.41362781541716e-05, 9.41362781541716e-05, 9.41362781541716e-05, 
    9.41362781541716e-05, 9.41362781541716e-05, 9.41362781541716e-05, 
    9.41362781541716e-05, 9.41362781541716e-05, 9.41362781541716e-05, 
    9.41362781541716e-05, 9.41362781541716e-05, 9.41362781541716e-05, 
    9.41362781541716e-05, 9.41362781541716e-05, 9.41362781541716e-05, 
    9.41362781541716e-05, 9.41362781541716e-05, 9.41362781541716e-05, 
    9.41362781541716e-05, 9.41362781541716e-05, 9.41362781541716e-05, 
    9.41362781541716e-05, 9.41362781541716e-05, 9.41362781541716e-05, 
    9.41362781541716e-05, 9.41362781541716e-05, 9.41362781541716e-05, 
    9.41362781541716e-05, 9.41362781541716e-05, 9.41362781541716e-05, 
    9.41362781541716e-05, 9.41362781541716e-05, 9.41362781541716e-05, 
    9.41362781541716e-05, 9.41362781541716e-05, 9.41362781541716e-05, 
    9.41362781541716e-05, 9.41362781541716e-05, 9.41362781541716e-05, 
    9.41362781541716e-05, 9.41362781541716e-05, 9.41362781541716e-05, 
    9.41362781541716e-05, 9.41362781541716e-05, 9.41362781541716e-05, 
    9.41362781541716e-05, 9.41362781541716e-05, 9.41362781541716e-05, 
    9.41362781541716e-05, 9.41362781541716e-05,
  9.47797019779707e-05, 9.47797019779707e-05, 9.47797019779707e-05, 
    9.47797019779707e-05, 9.47797019779707e-05, 9.47797019779707e-05, 
    9.47797019779707e-05, 9.47797019779707e-05, 9.47797019779707e-05, 
    9.47797019779707e-05, 9.47797019779707e-05, 9.47797019779707e-05, 
    9.47797019779707e-05, 9.47797019779707e-05, 9.47797019779707e-05, 
    9.47797019779707e-05, 9.47797019779707e-05, 9.47797019779707e-05, 
    9.47797019779707e-05, 9.47797019779707e-05, 9.47797019779707e-05, 
    9.47797019779707e-05, 9.47797019779707e-05, 9.47797019779707e-05, 
    9.47797019779707e-05, 9.47797019779707e-05, 9.47797019779707e-05, 
    9.47797019779707e-05, 9.47797019779707e-05, 9.47797019779707e-05, 
    9.47797019779707e-05, 9.47797019779707e-05, 9.47797019779707e-05, 
    9.47797019779707e-05, 9.47797019779707e-05, 9.47797019779707e-05, 
    9.47797019779707e-05, 9.47797019779707e-05, 9.47797019779707e-05, 
    9.47797019779707e-05, 9.47797019779707e-05, 9.47797019779707e-05, 
    9.47797019779707e-05, 9.47797019779707e-05, 9.47797019779707e-05, 
    9.47797019779707e-05, 9.47797019779707e-05, 9.47797019779707e-05, 
    9.47797019779707e-05, 9.47797019779707e-05, 9.47797019779707e-05, 
    9.47797019779707e-05, 9.47797019779707e-05, 9.47797019779707e-05, 
    9.47797019779707e-05, 9.47797019779707e-05,
  9.54199178610107e-05, 9.54199178610107e-05, 9.54199178610107e-05, 
    9.54199178610107e-05, 9.54199178610107e-05, 9.54199178610107e-05, 
    9.54199178610107e-05, 9.54199178610107e-05, 9.54199178610107e-05, 
    9.54199178610107e-05, 9.54199178610107e-05, 9.54199178610107e-05, 
    9.54199178610107e-05, 9.54199178610107e-05, 9.54199178610107e-05, 
    9.54199178610107e-05, 9.54199178610107e-05, 9.54199178610107e-05, 
    9.54199178610107e-05, 9.54199178610107e-05, 9.54199178610107e-05, 
    9.54199178610107e-05, 9.54199178610107e-05, 9.54199178610107e-05, 
    9.54199178610107e-05, 9.54199178610107e-05, 9.54199178610107e-05, 
    9.54199178610107e-05, 9.54199178610107e-05, 9.54199178610107e-05, 
    9.54199178610107e-05, 9.54199178610107e-05, 9.54199178610107e-05, 
    9.54199178610107e-05, 9.54199178610107e-05, 9.54199178610107e-05, 
    9.54199178610107e-05, 9.54199178610107e-05, 9.54199178610107e-05, 
    9.54199178610107e-05, 9.54199178610107e-05, 9.54199178610107e-05, 
    9.54199178610107e-05, 9.54199178610107e-05, 9.54199178610107e-05, 
    9.54199178610107e-05, 9.54199178610107e-05, 9.54199178610107e-05, 
    9.54199178610107e-05, 9.54199178610107e-05, 9.54199178610107e-05, 
    9.54199178610107e-05, 9.54199178610107e-05, 9.54199178610107e-05, 
    9.54199178610107e-05, 9.54199178610107e-05,
  9.60569041343627e-05, 9.60569041343627e-05, 9.60569041343627e-05, 
    9.60569041343627e-05, 9.60569041343627e-05, 9.60569041343627e-05, 
    9.60569041343627e-05, 9.60569041343627e-05, 9.60569041343627e-05, 
    9.60569041343627e-05, 9.60569041343627e-05, 9.60569041343627e-05, 
    9.60569041343627e-05, 9.60569041343627e-05, 9.60569041343627e-05, 
    9.60569041343627e-05, 9.60569041343627e-05, 9.60569041343627e-05, 
    9.60569041343627e-05, 9.60569041343627e-05, 9.60569041343627e-05, 
    9.60569041343627e-05, 9.60569041343627e-05, 9.60569041343627e-05, 
    9.60569041343627e-05, 9.60569041343627e-05, 9.60569041343627e-05, 
    9.60569041343627e-05, 9.60569041343627e-05, 9.60569041343627e-05, 
    9.60569041343627e-05, 9.60569041343627e-05, 9.60569041343627e-05, 
    9.60569041343627e-05, 9.60569041343627e-05, 9.60569041343627e-05, 
    9.60569041343627e-05, 9.60569041343627e-05, 9.60569041343627e-05, 
    9.60569041343627e-05, 9.60569041343627e-05, 9.60569041343627e-05, 
    9.60569041343627e-05, 9.60569041343627e-05, 9.60569041343627e-05, 
    9.60569041343627e-05, 9.60569041343627e-05, 9.60569041343627e-05, 
    9.60569041343627e-05, 9.60569041343627e-05, 9.60569041343627e-05, 
    9.60569041343627e-05, 9.60569041343627e-05, 9.60569041343627e-05, 
    9.60569041343627e-05, 9.60569041343627e-05,
  9.66906392384081e-05, 9.66906392384081e-05, 9.66906392384081e-05, 
    9.66906392384081e-05, 9.66906392384081e-05, 9.66906392384081e-05, 
    9.66906392384081e-05, 9.66906392384081e-05, 9.66906392384081e-05, 
    9.66906392384081e-05, 9.66906392384081e-05, 9.66906392384081e-05, 
    9.66906392384081e-05, 9.66906392384081e-05, 9.66906392384081e-05, 
    9.66906392384081e-05, 9.66906392384081e-05, 9.66906392384081e-05, 
    9.66906392384081e-05, 9.66906392384081e-05, 9.66906392384081e-05, 
    9.66906392384081e-05, 9.66906392384081e-05, 9.66906392384081e-05, 
    9.66906392384081e-05, 9.66906392384081e-05, 9.66906392384081e-05, 
    9.66906392384081e-05, 9.66906392384081e-05, 9.66906392384081e-05, 
    9.66906392384081e-05, 9.66906392384081e-05, 9.66906392384081e-05, 
    9.66906392384081e-05, 9.66906392384081e-05, 9.66906392384081e-05, 
    9.66906392384081e-05, 9.66906392384081e-05, 9.66906392384081e-05, 
    9.66906392384081e-05, 9.66906392384081e-05, 9.66906392384081e-05, 
    9.66906392384081e-05, 9.66906392384081e-05, 9.66906392384081e-05, 
    9.66906392384081e-05, 9.66906392384081e-05, 9.66906392384081e-05, 
    9.66906392384081e-05, 9.66906392384081e-05, 9.66906392384081e-05, 
    9.66906392384081e-05, 9.66906392384081e-05, 9.66906392384081e-05, 
    9.66906392384081e-05, 9.66906392384081e-05,
  9.73211017235682e-05, 9.73211017235682e-05, 9.73211017235682e-05, 
    9.73211017235682e-05, 9.73211017235682e-05, 9.73211017235682e-05, 
    9.73211017235682e-05, 9.73211017235682e-05, 9.73211017235682e-05, 
    9.73211017235682e-05, 9.73211017235682e-05, 9.73211017235682e-05, 
    9.73211017235682e-05, 9.73211017235682e-05, 9.73211017235682e-05, 
    9.73211017235682e-05, 9.73211017235682e-05, 9.73211017235682e-05, 
    9.73211017235682e-05, 9.73211017235682e-05, 9.73211017235682e-05, 
    9.73211017235682e-05, 9.73211017235682e-05, 9.73211017235682e-05, 
    9.73211017235682e-05, 9.73211017235682e-05, 9.73211017235682e-05, 
    9.73211017235682e-05, 9.73211017235682e-05, 9.73211017235682e-05, 
    9.73211017235682e-05, 9.73211017235682e-05, 9.73211017235682e-05, 
    9.73211017235682e-05, 9.73211017235682e-05, 9.73211017235682e-05, 
    9.73211017235682e-05, 9.73211017235682e-05, 9.73211017235682e-05, 
    9.73211017235682e-05, 9.73211017235682e-05, 9.73211017235682e-05, 
    9.73211017235682e-05, 9.73211017235682e-05, 9.73211017235682e-05, 
    9.73211017235682e-05, 9.73211017235682e-05, 9.73211017235682e-05, 
    9.73211017235682e-05, 9.73211017235682e-05, 9.73211017235682e-05, 
    9.73211017235682e-05, 9.73211017235682e-05, 9.73211017235682e-05, 
    9.73211017235682e-05, 9.73211017235682e-05,
  9.79482702510304e-05, 9.79482702510304e-05, 9.79482702510304e-05, 
    9.79482702510304e-05, 9.79482702510304e-05, 9.79482702510304e-05, 
    9.79482702510304e-05, 9.79482702510304e-05, 9.79482702510304e-05, 
    9.79482702510304e-05, 9.79482702510304e-05, 9.79482702510304e-05, 
    9.79482702510304e-05, 9.79482702510304e-05, 9.79482702510304e-05, 
    9.79482702510304e-05, 9.79482702510304e-05, 9.79482702510304e-05, 
    9.79482702510304e-05, 9.79482702510304e-05, 9.79482702510304e-05, 
    9.79482702510304e-05, 9.79482702510304e-05, 9.79482702510304e-05, 
    9.79482702510304e-05, 9.79482702510304e-05, 9.79482702510304e-05, 
    9.79482702510304e-05, 9.79482702510304e-05, 9.79482702510304e-05, 
    9.79482702510304e-05, 9.79482702510304e-05, 9.79482702510304e-05, 
    9.79482702510304e-05, 9.79482702510304e-05, 9.79482702510304e-05, 
    9.79482702510304e-05, 9.79482702510304e-05, 9.79482702510304e-05, 
    9.79482702510304e-05, 9.79482702510304e-05, 9.79482702510304e-05, 
    9.79482702510304e-05, 9.79482702510304e-05, 9.79482702510304e-05, 
    9.79482702510304e-05, 9.79482702510304e-05, 9.79482702510304e-05, 
    9.79482702510304e-05, 9.79482702510304e-05, 9.79482702510304e-05, 
    9.79482702510304e-05, 9.79482702510304e-05, 9.79482702510304e-05, 
    9.79482702510304e-05, 9.79482702510304e-05,
  9.85721235934702e-05, 9.85721235934702e-05, 9.85721235934702e-05, 
    9.85721235934702e-05, 9.85721235934702e-05, 9.85721235934702e-05, 
    9.85721235934702e-05, 9.85721235934702e-05, 9.85721235934702e-05, 
    9.85721235934702e-05, 9.85721235934702e-05, 9.85721235934702e-05, 
    9.85721235934702e-05, 9.85721235934702e-05, 9.85721235934702e-05, 
    9.85721235934702e-05, 9.85721235934702e-05, 9.85721235934702e-05, 
    9.85721235934702e-05, 9.85721235934702e-05, 9.85721235934702e-05, 
    9.85721235934702e-05, 9.85721235934702e-05, 9.85721235934702e-05, 
    9.85721235934702e-05, 9.85721235934702e-05, 9.85721235934702e-05, 
    9.85721235934702e-05, 9.85721235934702e-05, 9.85721235934702e-05, 
    9.85721235934702e-05, 9.85721235934702e-05, 9.85721235934702e-05, 
    9.85721235934702e-05, 9.85721235934702e-05, 9.85721235934702e-05, 
    9.85721235934702e-05, 9.85721235934702e-05, 9.85721235934702e-05, 
    9.85721235934702e-05, 9.85721235934702e-05, 9.85721235934702e-05, 
    9.85721235934702e-05, 9.85721235934702e-05, 9.85721235934702e-05, 
    9.85721235934702e-05, 9.85721235934702e-05, 9.85721235934702e-05, 
    9.85721235934702e-05, 9.85721235934702e-05, 9.85721235934702e-05, 
    9.85721235934702e-05, 9.85721235934702e-05, 9.85721235934702e-05, 
    9.85721235934702e-05, 9.85721235934702e-05,
  9.919264063577e-05, 9.919264063577e-05, 9.919264063577e-05, 
    9.919264063577e-05, 9.919264063577e-05, 9.919264063577e-05, 
    9.919264063577e-05, 9.919264063577e-05, 9.919264063577e-05, 
    9.919264063577e-05, 9.919264063577e-05, 9.919264063577e-05, 
    9.919264063577e-05, 9.919264063577e-05, 9.919264063577e-05, 
    9.919264063577e-05, 9.919264063577e-05, 9.919264063577e-05, 
    9.919264063577e-05, 9.919264063577e-05, 9.919264063577e-05, 
    9.919264063577e-05, 9.919264063577e-05, 9.919264063577e-05, 
    9.919264063577e-05, 9.919264063577e-05, 9.919264063577e-05, 
    9.919264063577e-05, 9.919264063577e-05, 9.919264063577e-05, 
    9.919264063577e-05, 9.919264063577e-05, 9.919264063577e-05, 
    9.919264063577e-05, 9.919264063577e-05, 9.919264063577e-05, 
    9.919264063577e-05, 9.919264063577e-05, 9.919264063577e-05, 
    9.919264063577e-05, 9.919264063577e-05, 9.919264063577e-05, 
    9.919264063577e-05, 9.919264063577e-05, 9.919264063577e-05, 
    9.919264063577e-05, 9.919264063577e-05, 9.919264063577e-05, 
    9.919264063577e-05, 9.919264063577e-05, 9.919264063577e-05, 
    9.919264063577e-05, 9.919264063577e-05, 9.919264063577e-05, 
    9.919264063577e-05, 9.919264063577e-05,
  9.98098003757333e-05, 9.98098003757333e-05, 9.98098003757333e-05, 
    9.98098003757333e-05, 9.98098003757333e-05, 9.98098003757333e-05, 
    9.98098003757333e-05, 9.98098003757333e-05, 9.98098003757333e-05, 
    9.98098003757333e-05, 9.98098003757333e-05, 9.98098003757333e-05, 
    9.98098003757333e-05, 9.98098003757333e-05, 9.98098003757333e-05, 
    9.98098003757333e-05, 9.98098003757333e-05, 9.98098003757333e-05, 
    9.98098003757333e-05, 9.98098003757333e-05, 9.98098003757333e-05, 
    9.98098003757333e-05, 9.98098003757333e-05, 9.98098003757333e-05, 
    9.98098003757333e-05, 9.98098003757333e-05, 9.98098003757333e-05, 
    9.98098003757333e-05, 9.98098003757333e-05, 9.98098003757333e-05, 
    9.98098003757333e-05, 9.98098003757333e-05, 9.98098003757333e-05, 
    9.98098003757333e-05, 9.98098003757333e-05, 9.98098003757333e-05, 
    9.98098003757333e-05, 9.98098003757333e-05, 9.98098003757333e-05, 
    9.98098003757333e-05, 9.98098003757333e-05, 9.98098003757333e-05, 
    9.98098003757333e-05, 9.98098003757333e-05, 9.98098003757333e-05, 
    9.98098003757333e-05, 9.98098003757333e-05, 9.98098003757333e-05, 
    9.98098003757333e-05, 9.98098003757333e-05, 9.98098003757333e-05, 
    9.98098003757333e-05, 9.98098003757333e-05, 9.98098003757333e-05, 
    9.98098003757333e-05, 9.98098003757333e-05,
  0.000100423581924796, 0.000100423581924796, 0.000100423581924796, 
    0.000100423581924796, 0.000100423581924796, 0.000100423581924796, 
    0.000100423581924796, 0.000100423581924796, 0.000100423581924796, 
    0.000100423581924796, 0.000100423581924796, 0.000100423581924796, 
    0.000100423581924796, 0.000100423581924796, 0.000100423581924796, 
    0.000100423581924796, 0.000100423581924796, 0.000100423581924796, 
    0.000100423581924796, 0.000100423581924796, 0.000100423581924796, 
    0.000100423581924796, 0.000100423581924796, 0.000100423581924796, 
    0.000100423581924796, 0.000100423581924796, 0.000100423581924796, 
    0.000100423581924796, 0.000100423581924796, 0.000100423581924796, 
    0.000100423581924796, 0.000100423581924796, 0.000100423581924796, 
    0.000100423581924796, 0.000100423581924796, 0.000100423581924796, 
    0.000100423581924796, 0.000100423581924796, 0.000100423581924796, 
    0.000100423581924796, 0.000100423581924796, 0.000100423581924796, 
    0.000100423581924796, 0.000100423581924796, 0.000100423581924796, 
    0.000100423581924796, 0.000100423581924796, 0.000100423581924796, 
    0.000100423581924796, 0.000100423581924796, 0.000100423581924796, 
    0.000100423581924796, 0.000100423581924796, 0.000100423581924796, 
    0.000100423581924796, 0.000100423581924796,
  0.000101033964508733, 0.000101033964508733, 0.000101033964508733, 
    0.000101033964508733, 0.000101033964508733, 0.000101033964508733, 
    0.000101033964508733, 0.000101033964508733, 0.000101033964508733, 
    0.000101033964508733, 0.000101033964508733, 0.000101033964508733, 
    0.000101033964508733, 0.000101033964508733, 0.000101033964508733, 
    0.000101033964508733, 0.000101033964508733, 0.000101033964508733, 
    0.000101033964508733, 0.000101033964508733, 0.000101033964508733, 
    0.000101033964508733, 0.000101033964508733, 0.000101033964508733, 
    0.000101033964508733, 0.000101033964508733, 0.000101033964508733, 
    0.000101033964508733, 0.000101033964508733, 0.000101033964508733, 
    0.000101033964508733, 0.000101033964508733, 0.000101033964508733, 
    0.000101033964508733, 0.000101033964508733, 0.000101033964508733, 
    0.000101033964508733, 0.000101033964508733, 0.000101033964508733, 
    0.000101033964508733, 0.000101033964508733, 0.000101033964508733, 
    0.000101033964508733, 0.000101033964508733, 0.000101033964508733, 
    0.000101033964508733, 0.000101033964508733, 0.000101033964508733, 
    0.000101033964508733, 0.000101033964508733, 0.000101033964508733, 
    0.000101033964508733, 0.000101033964508733, 0.000101033964508733, 
    0.000101033964508733, 0.000101033964508733,
  0.000101640927468363, 0.000101640927468363, 0.000101640927468363, 
    0.000101640927468363, 0.000101640927468363, 0.000101640927468363, 
    0.000101640927468363, 0.000101640927468363, 0.000101640927468363, 
    0.000101640927468363, 0.000101640927468363, 0.000101640927468363, 
    0.000101640927468363, 0.000101640927468363, 0.000101640927468363, 
    0.000101640927468363, 0.000101640927468363, 0.000101640927468363, 
    0.000101640927468363, 0.000101640927468363, 0.000101640927468363, 
    0.000101640927468363, 0.000101640927468363, 0.000101640927468363, 
    0.000101640927468363, 0.000101640927468363, 0.000101640927468363, 
    0.000101640927468363, 0.000101640927468363, 0.000101640927468363, 
    0.000101640927468363, 0.000101640927468363, 0.000101640927468363, 
    0.000101640927468363, 0.000101640927468363, 0.000101640927468363, 
    0.000101640927468363, 0.000101640927468363, 0.000101640927468363, 
    0.000101640927468363, 0.000101640927468363, 0.000101640927468363, 
    0.000101640927468363, 0.000101640927468363, 0.000101640927468363, 
    0.000101640927468363, 0.000101640927468363, 0.000101640927468363, 
    0.000101640927468363, 0.000101640927468363, 0.000101640927468363, 
    0.000101640927468363, 0.000101640927468363, 0.000101640927468363, 
    0.000101640927468363, 0.000101640927468363,
  0.000102244450260243, 0.000102244450260243, 0.000102244450260243, 
    0.000102244450260243, 0.000102244450260243, 0.000102244450260243, 
    0.000102244450260243, 0.000102244450260243, 0.000102244450260243, 
    0.000102244450260243, 0.000102244450260243, 0.000102244450260243, 
    0.000102244450260243, 0.000102244450260243, 0.000102244450260243, 
    0.000102244450260243, 0.000102244450260243, 0.000102244450260243, 
    0.000102244450260243, 0.000102244450260243, 0.000102244450260243, 
    0.000102244450260243, 0.000102244450260243, 0.000102244450260243, 
    0.000102244450260243, 0.000102244450260243, 0.000102244450260243, 
    0.000102244450260243, 0.000102244450260243, 0.000102244450260243, 
    0.000102244450260243, 0.000102244450260243, 0.000102244450260243, 
    0.000102244450260243, 0.000102244450260243, 0.000102244450260243, 
    0.000102244450260243, 0.000102244450260243, 0.000102244450260243, 
    0.000102244450260243, 0.000102244450260243, 0.000102244450260243, 
    0.000102244450260243, 0.000102244450260243, 0.000102244450260243, 
    0.000102244450260243, 0.000102244450260243, 0.000102244450260243, 
    0.000102244450260243, 0.000102244450260243, 0.000102244450260243, 
    0.000102244450260243, 0.000102244450260243, 0.000102244450260243, 
    0.000102244450260243, 0.000102244450260243,
  0.00010284451245737, 0.00010284451245737, 0.00010284451245737, 
    0.00010284451245737, 0.00010284451245737, 0.00010284451245737, 
    0.00010284451245737, 0.00010284451245737, 0.00010284451245737, 
    0.00010284451245737, 0.00010284451245737, 0.00010284451245737, 
    0.00010284451245737, 0.00010284451245737, 0.00010284451245737, 
    0.00010284451245737, 0.00010284451245737, 0.00010284451245737, 
    0.00010284451245737, 0.00010284451245737, 0.00010284451245737, 
    0.00010284451245737, 0.00010284451245737, 0.00010284451245737, 
    0.00010284451245737, 0.00010284451245737, 0.00010284451245737, 
    0.00010284451245737, 0.00010284451245737, 0.00010284451245737, 
    0.00010284451245737, 0.00010284451245737, 0.00010284451245737, 
    0.00010284451245737, 0.00010284451245737, 0.00010284451245737, 
    0.00010284451245737, 0.00010284451245737, 0.00010284451245737, 
    0.00010284451245737, 0.00010284451245737, 0.00010284451245737, 
    0.00010284451245737, 0.00010284451245737, 0.00010284451245737, 
    0.00010284451245737, 0.00010284451245737, 0.00010284451245737, 
    0.00010284451245737, 0.00010284451245737, 0.00010284451245737, 
    0.00010284451245737, 0.00010284451245737, 0.00010284451245737, 
    0.00010284451245737, 0.00010284451245737,
  0.000103441093749867, 0.000103441093749867, 0.000103441093749867, 
    0.000103441093749867, 0.000103441093749867, 0.000103441093749867, 
    0.000103441093749867, 0.000103441093749867, 0.000103441093749867, 
    0.000103441093749867, 0.000103441093749867, 0.000103441093749867, 
    0.000103441093749867, 0.000103441093749867, 0.000103441093749867, 
    0.000103441093749867, 0.000103441093749867, 0.000103441093749867, 
    0.000103441093749867, 0.000103441093749867, 0.000103441093749867, 
    0.000103441093749867, 0.000103441093749867, 0.000103441093749867, 
    0.000103441093749867, 0.000103441093749867, 0.000103441093749867, 
    0.000103441093749867, 0.000103441093749867, 0.000103441093749867, 
    0.000103441093749867, 0.000103441093749867, 0.000103441093749867, 
    0.000103441093749867, 0.000103441093749867, 0.000103441093749867, 
    0.000103441093749867, 0.000103441093749867, 0.000103441093749867, 
    0.000103441093749867, 0.000103441093749867, 0.000103441093749867, 
    0.000103441093749867, 0.000103441093749867, 0.000103441093749867, 
    0.000103441093749867, 0.000103441093749867, 0.000103441093749867, 
    0.000103441093749867, 0.000103441093749867, 0.000103441093749867, 
    0.000103441093749867, 0.000103441093749867, 0.000103441093749867, 
    0.000103441093749867, 0.000103441093749867,
  0.000104034173945676, 0.000104034173945676, 0.000104034173945676, 
    0.000104034173945676, 0.000104034173945676, 0.000104034173945676, 
    0.000104034173945676, 0.000104034173945676, 0.000104034173945676, 
    0.000104034173945676, 0.000104034173945676, 0.000104034173945676, 
    0.000104034173945676, 0.000104034173945676, 0.000104034173945676, 
    0.000104034173945676, 0.000104034173945676, 0.000104034173945676, 
    0.000104034173945676, 0.000104034173945676, 0.000104034173945676, 
    0.000104034173945676, 0.000104034173945676, 0.000104034173945676, 
    0.000104034173945676, 0.000104034173945676, 0.000104034173945676, 
    0.000104034173945676, 0.000104034173945676, 0.000104034173945676, 
    0.000104034173945676, 0.000104034173945676, 0.000104034173945676, 
    0.000104034173945676, 0.000104034173945676, 0.000104034173945676, 
    0.000104034173945676, 0.000104034173945676, 0.000104034173945676, 
    0.000104034173945676, 0.000104034173945676, 0.000104034173945676, 
    0.000104034173945676, 0.000104034173945676, 0.000104034173945676, 
    0.000104034173945676, 0.000104034173945676, 0.000104034173945676, 
    0.000104034173945676, 0.000104034173945676, 0.000104034173945676, 
    0.000104034173945676, 0.000104034173945676, 0.000104034173945676, 
    0.000104034173945676, 0.000104034173945676,
  0.000104623732971234, 0.000104623732971234, 0.000104623732971234, 
    0.000104623732971234, 0.000104623732971234, 0.000104623732971234, 
    0.000104623732971234, 0.000104623732971234, 0.000104623732971234, 
    0.000104623732971234, 0.000104623732971234, 0.000104623732971234, 
    0.000104623732971234, 0.000104623732971234, 0.000104623732971234, 
    0.000104623732971234, 0.000104623732971234, 0.000104623732971234, 
    0.000104623732971234, 0.000104623732971234, 0.000104623732971234, 
    0.000104623732971234, 0.000104623732971234, 0.000104623732971234, 
    0.000104623732971234, 0.000104623732971234, 0.000104623732971234, 
    0.000104623732971234, 0.000104623732971234, 0.000104623732971234, 
    0.000104623732971234, 0.000104623732971234, 0.000104623732971234, 
    0.000104623732971234, 0.000104623732971234, 0.000104623732971234, 
    0.000104623732971234, 0.000104623732971234, 0.000104623732971234, 
    0.000104623732971234, 0.000104623732971234, 0.000104623732971234, 
    0.000104623732971234, 0.000104623732971234, 0.000104623732971234, 
    0.000104623732971234, 0.000104623732971234, 0.000104623732971234, 
    0.000104623732971234, 0.000104623732971234, 0.000104623732971234, 
    0.000104623732971234, 0.000104623732971234, 0.000104623732971234, 
    0.000104623732971234, 0.000104623732971234,
  0.000105209750872159, 0.000105209750872159, 0.000105209750872159, 
    0.000105209750872159, 0.000105209750872159, 0.000105209750872159, 
    0.000105209750872159, 0.000105209750872159, 0.000105209750872159, 
    0.000105209750872159, 0.000105209750872159, 0.000105209750872159, 
    0.000105209750872159, 0.000105209750872159, 0.000105209750872159, 
    0.000105209750872159, 0.000105209750872159, 0.000105209750872159, 
    0.000105209750872159, 0.000105209750872159, 0.000105209750872159, 
    0.000105209750872159, 0.000105209750872159, 0.000105209750872159, 
    0.000105209750872159, 0.000105209750872159, 0.000105209750872159, 
    0.000105209750872159, 0.000105209750872159, 0.000105209750872159, 
    0.000105209750872159, 0.000105209750872159, 0.000105209750872159, 
    0.000105209750872159, 0.000105209750872159, 0.000105209750872159, 
    0.000105209750872159, 0.000105209750872159, 0.000105209750872159, 
    0.000105209750872159, 0.000105209750872159, 0.000105209750872159, 
    0.000105209750872159, 0.000105209750872159, 0.000105209750872159, 
    0.000105209750872159, 0.000105209750872159, 0.000105209750872159, 
    0.000105209750872159, 0.000105209750872159, 0.000105209750872159, 
    0.000105209750872159, 0.000105209750872159, 0.000105209750872159, 
    0.000105209750872159, 0.000105209750872159,
  0.000105792207813923, 0.000105792207813923, 0.000105792207813923, 
    0.000105792207813923, 0.000105792207813923, 0.000105792207813923, 
    0.000105792207813923, 0.000105792207813923, 0.000105792207813923, 
    0.000105792207813923, 0.000105792207813923, 0.000105792207813923, 
    0.000105792207813923, 0.000105792207813923, 0.000105792207813923, 
    0.000105792207813923, 0.000105792207813923, 0.000105792207813923, 
    0.000105792207813923, 0.000105792207813923, 0.000105792207813923, 
    0.000105792207813923, 0.000105792207813923, 0.000105792207813923, 
    0.000105792207813923, 0.000105792207813923, 0.000105792207813923, 
    0.000105792207813923, 0.000105792207813923, 0.000105792207813923, 
    0.000105792207813923, 0.000105792207813923, 0.000105792207813923, 
    0.000105792207813923, 0.000105792207813923, 0.000105792207813923, 
    0.000105792207813923, 0.000105792207813923, 0.000105792207813923, 
    0.000105792207813923, 0.000105792207813923, 0.000105792207813923, 
    0.000105792207813923, 0.000105792207813923, 0.000105792207813923, 
    0.000105792207813923, 0.000105792207813923, 0.000105792207813923, 
    0.000105792207813923, 0.000105792207813923, 0.000105792207813923, 
    0.000105792207813923, 0.000105792207813923, 0.000105792207813923, 
    0.000105792207813923, 0.000105792207813923,
  0.000106371084082523, 0.000106371084082523, 0.000106371084082523, 
    0.000106371084082523, 0.000106371084082523, 0.000106371084082523, 
    0.000106371084082523, 0.000106371084082523, 0.000106371084082523, 
    0.000106371084082523, 0.000106371084082523, 0.000106371084082523, 
    0.000106371084082523, 0.000106371084082523, 0.000106371084082523, 
    0.000106371084082523, 0.000106371084082523, 0.000106371084082523, 
    0.000106371084082523, 0.000106371084082523, 0.000106371084082523, 
    0.000106371084082523, 0.000106371084082523, 0.000106371084082523, 
    0.000106371084082523, 0.000106371084082523, 0.000106371084082523, 
    0.000106371084082523, 0.000106371084082523, 0.000106371084082523, 
    0.000106371084082523, 0.000106371084082523, 0.000106371084082523, 
    0.000106371084082523, 0.000106371084082523, 0.000106371084082523, 
    0.000106371084082523, 0.000106371084082523, 0.000106371084082523, 
    0.000106371084082523, 0.000106371084082523, 0.000106371084082523, 
    0.000106371084082523, 0.000106371084082523, 0.000106371084082523, 
    0.000106371084082523, 0.000106371084082523, 0.000106371084082523, 
    0.000106371084082523, 0.000106371084082523, 0.000106371084082523, 
    0.000106371084082523, 0.000106371084082523, 0.000106371084082523, 
    0.000106371084082523, 0.000106371084082523,
  0.000106946360085146, 0.000106946360085146, 0.000106946360085146, 
    0.000106946360085146, 0.000106946360085146, 0.000106946360085146, 
    0.000106946360085146, 0.000106946360085146, 0.000106946360085146, 
    0.000106946360085146, 0.000106946360085146, 0.000106946360085146, 
    0.000106946360085146, 0.000106946360085146, 0.000106946360085146, 
    0.000106946360085146, 0.000106946360085146, 0.000106946360085146, 
    0.000106946360085146, 0.000106946360085146, 0.000106946360085146, 
    0.000106946360085146, 0.000106946360085146, 0.000106946360085146, 
    0.000106946360085146, 0.000106946360085146, 0.000106946360085146, 
    0.000106946360085146, 0.000106946360085146, 0.000106946360085146, 
    0.000106946360085146, 0.000106946360085146, 0.000106946360085146, 
    0.000106946360085146, 0.000106946360085146, 0.000106946360085146, 
    0.000106946360085146, 0.000106946360085146, 0.000106946360085146, 
    0.000106946360085146, 0.000106946360085146, 0.000106946360085146, 
    0.000106946360085146, 0.000106946360085146, 0.000106946360085146, 
    0.000106946360085146, 0.000106946360085146, 0.000106946360085146, 
    0.000106946360085146, 0.000106946360085146, 0.000106946360085146, 
    0.000106946360085146, 0.000106946360085146, 0.000106946360085146, 
    0.000106946360085146, 0.000106946360085146,
  0.000107518016350839, 0.000107518016350839, 0.000107518016350839, 
    0.000107518016350839, 0.000107518016350839, 0.000107518016350839, 
    0.000107518016350839, 0.000107518016350839, 0.000107518016350839, 
    0.000107518016350839, 0.000107518016350839, 0.000107518016350839, 
    0.000107518016350839, 0.000107518016350839, 0.000107518016350839, 
    0.000107518016350839, 0.000107518016350839, 0.000107518016350839, 
    0.000107518016350839, 0.000107518016350839, 0.000107518016350839, 
    0.000107518016350839, 0.000107518016350839, 0.000107518016350839, 
    0.000107518016350839, 0.000107518016350839, 0.000107518016350839, 
    0.000107518016350839, 0.000107518016350839, 0.000107518016350839, 
    0.000107518016350839, 0.000107518016350839, 0.000107518016350839, 
    0.000107518016350839, 0.000107518016350839, 0.000107518016350839, 
    0.000107518016350839, 0.000107518016350839, 0.000107518016350839, 
    0.000107518016350839, 0.000107518016350839, 0.000107518016350839, 
    0.000107518016350839, 0.000107518016350839, 0.000107518016350839, 
    0.000107518016350839, 0.000107518016350839, 0.000107518016350839, 
    0.000107518016350839, 0.000107518016350839, 0.000107518016350839, 
    0.000107518016350839, 0.000107518016350839, 0.000107518016350839, 
    0.000107518016350839, 0.000107518016350839,
  0.00010808603353116, 0.00010808603353116, 0.00010808603353116, 
    0.00010808603353116, 0.00010808603353116, 0.00010808603353116, 
    0.00010808603353116, 0.00010808603353116, 0.00010808603353116, 
    0.00010808603353116, 0.00010808603353116, 0.00010808603353116, 
    0.00010808603353116, 0.00010808603353116, 0.00010808603353116, 
    0.00010808603353116, 0.00010808603353116, 0.00010808603353116, 
    0.00010808603353116, 0.00010808603353116, 0.00010808603353116, 
    0.00010808603353116, 0.00010808603353116, 0.00010808603353116, 
    0.00010808603353116, 0.00010808603353116, 0.00010808603353116, 
    0.00010808603353116, 0.00010808603353116, 0.00010808603353116, 
    0.00010808603353116, 0.00010808603353116, 0.00010808603353116, 
    0.00010808603353116, 0.00010808603353116, 0.00010808603353116, 
    0.00010808603353116, 0.00010808603353116, 0.00010808603353116, 
    0.00010808603353116, 0.00010808603353116, 0.00010808603353116, 
    0.00010808603353116, 0.00010808603353116, 0.00010808603353116, 
    0.00010808603353116, 0.00010808603353116, 0.00010808603353116, 
    0.00010808603353116, 0.00010808603353116, 0.00010808603353116, 
    0.00010808603353116, 0.00010808603353116, 0.00010808603353116, 
    0.00010808603353116, 0.00010808603353116 ;

 pm =
  3.11708294538134e-05, 3.11708294538134e-05, 3.11708294538134e-05, 
    3.1170829453808e-05, 3.11708294538134e-05, 3.11708294538134e-05, 
    3.1170829453808e-05, 3.11708294538134e-05, 3.11708294538134e-05, 
    3.1170829453808e-05, 3.11708294538134e-05, 3.11708294538134e-05, 
    3.1170829453808e-05, 3.11708294538134e-05, 3.11708294538134e-05, 
    3.1170829453808e-05, 3.11708294538134e-05, 3.11708294538134e-05, 
    3.11708294538107e-05, 3.11708294538107e-05, 3.11708294538107e-05, 
    3.11708294538134e-05, 3.11708294538107e-05, 3.11708294538107e-05, 
    3.11708294538134e-05, 3.11708294538107e-05, 3.11708294538107e-05, 
    3.11708294538134e-05, 3.11708294538107e-05, 3.11708294538107e-05, 
    3.11708294538134e-05, 3.11708294538107e-05, 3.11708294538107e-05, 
    3.11708294538134e-05, 3.11708294538107e-05, 3.11708294538107e-05, 
    3.11708294538134e-05, 3.11708294538107e-05, 3.11708294538107e-05, 
    3.11708294538134e-05, 3.11708294538107e-05, 3.11708294538107e-05, 
    3.11708294538134e-05, 3.11708294538107e-05, 3.11708294538107e-05, 
    3.11708294538134e-05, 3.11708294538107e-05, 3.11708294538107e-05, 
    3.11708294538134e-05, 3.11708294538107e-05, 3.1170829453812e-05, 
    3.1170829453812e-05, 3.11708294538107e-05, 3.1170829453812e-05, 
    3.1170829453812e-05, 3.1170829453812e-05,
  3.12764123356491e-05, 3.12764123356491e-05, 3.12764123356491e-05, 
    3.12764123356438e-05, 3.12764123356491e-05, 3.12764123356491e-05, 
    3.12764123356438e-05, 3.12764123356491e-05, 3.12764123356491e-05, 
    3.12764123356438e-05, 3.12764123356491e-05, 3.12764123356491e-05, 
    3.12764123356438e-05, 3.12764123356491e-05, 3.12764123356491e-05, 
    3.12764123356438e-05, 3.12764123356491e-05, 3.12764123356491e-05, 
    3.12764123356464e-05, 3.12764123356464e-05, 3.12764123356464e-05, 
    3.12764123356491e-05, 3.12764123356464e-05, 3.12764123356464e-05, 
    3.12764123356491e-05, 3.12764123356464e-05, 3.12764123356464e-05, 
    3.12764123356491e-05, 3.12764123356464e-05, 3.12764123356464e-05, 
    3.12764123356491e-05, 3.12764123356464e-05, 3.12764123356464e-05, 
    3.12764123356491e-05, 3.12764123356464e-05, 3.12764123356464e-05, 
    3.12764123356491e-05, 3.12764123356464e-05, 3.12764123356464e-05, 
    3.12764123356491e-05, 3.12764123356464e-05, 3.12764123356464e-05, 
    3.12764123356491e-05, 3.12764123356464e-05, 3.12764123356464e-05, 
    3.12764123356491e-05, 3.12764123356464e-05, 3.12764123356464e-05, 
    3.12764123356491e-05, 3.12764123356464e-05, 3.12764123356478e-05, 
    3.12764123356478e-05, 3.12764123356464e-05, 3.12764123356478e-05, 
    3.12764123356478e-05, 3.12764123356478e-05,
  3.13837787507492e-05, 3.13837787507492e-05, 3.13837787507492e-05, 
    3.13837787507439e-05, 3.13837787507492e-05, 3.13837787507492e-05, 
    3.13837787507439e-05, 3.13837787507492e-05, 3.13837787507492e-05, 
    3.13837787507439e-05, 3.13837787507492e-05, 3.13837787507492e-05, 
    3.13837787507439e-05, 3.13837787507492e-05, 3.13837787507492e-05, 
    3.13837787507439e-05, 3.13837787507492e-05, 3.13837787507492e-05, 
    3.13837787507465e-05, 3.13837787507465e-05, 3.13837787507465e-05, 
    3.13837787507492e-05, 3.13837787507465e-05, 3.13837787507465e-05, 
    3.13837787507492e-05, 3.13837787507465e-05, 3.13837787507465e-05, 
    3.13837787507492e-05, 3.13837787507465e-05, 3.13837787507465e-05, 
    3.13837787507492e-05, 3.13837787507465e-05, 3.13837787507465e-05, 
    3.13837787507492e-05, 3.13837787507465e-05, 3.13837787507465e-05, 
    3.13837787507492e-05, 3.13837787507465e-05, 3.13837787507465e-05, 
    3.13837787507492e-05, 3.13837787507465e-05, 3.13837787507465e-05, 
    3.13837787507492e-05, 3.13837787507465e-05, 3.13837787507465e-05, 
    3.13837787507492e-05, 3.13837787507465e-05, 3.13837787507465e-05, 
    3.13837787507492e-05, 3.13837787507465e-05, 3.13837787507479e-05, 
    3.13837787507479e-05, 3.13837787507465e-05, 3.13837787507479e-05, 
    3.13837787507479e-05, 3.13837787507479e-05,
  3.14929544361165e-05, 3.14929544361165e-05, 3.14929544361165e-05, 
    3.14929544361111e-05, 3.14929544361165e-05, 3.14929544361165e-05, 
    3.14929544361111e-05, 3.14929544361165e-05, 3.14929544361165e-05, 
    3.14929544361111e-05, 3.14929544361165e-05, 3.14929544361165e-05, 
    3.14929544361111e-05, 3.14929544361165e-05, 3.14929544361165e-05, 
    3.14929544361111e-05, 3.14929544361165e-05, 3.14929544361165e-05, 
    3.14929544361138e-05, 3.14929544361138e-05, 3.14929544361138e-05, 
    3.14929544361165e-05, 3.14929544361138e-05, 3.14929544361138e-05, 
    3.14929544361165e-05, 3.14929544361138e-05, 3.14929544361138e-05, 
    3.14929544361165e-05, 3.14929544361138e-05, 3.14929544361138e-05, 
    3.14929544361165e-05, 3.14929544361138e-05, 3.14929544361138e-05, 
    3.14929544361165e-05, 3.14929544361138e-05, 3.14929544361138e-05, 
    3.14929544361165e-05, 3.14929544361138e-05, 3.14929544361138e-05, 
    3.14929544361165e-05, 3.14929544361138e-05, 3.14929544361138e-05, 
    3.14929544361165e-05, 3.14929544361138e-05, 3.14929544361138e-05, 
    3.14929544361165e-05, 3.14929544361138e-05, 3.14929544361138e-05, 
    3.14929544361165e-05, 3.14929544361138e-05, 3.14929544361151e-05, 
    3.14929544361151e-05, 3.14929544361138e-05, 3.14929544361151e-05, 
    3.14929544361151e-05, 3.14929544361151e-05,
  3.16039657692524e-05, 3.16039657692524e-05, 3.16039657692524e-05, 
    3.1603965769247e-05, 3.16039657692524e-05, 3.16039657692524e-05, 
    3.1603965769247e-05, 3.16039657692524e-05, 3.16039657692524e-05, 
    3.1603965769247e-05, 3.16039657692524e-05, 3.16039657692524e-05, 
    3.1603965769247e-05, 3.16039657692524e-05, 3.16039657692524e-05, 
    3.1603965769247e-05, 3.16039657692524e-05, 3.16039657692524e-05, 
    3.16039657692497e-05, 3.16039657692497e-05, 3.16039657692497e-05, 
    3.16039657692524e-05, 3.16039657692497e-05, 3.16039657692497e-05, 
    3.16039657692524e-05, 3.16039657692497e-05, 3.16039657692497e-05, 
    3.16039657692524e-05, 3.16039657692497e-05, 3.16039657692497e-05, 
    3.16039657692524e-05, 3.16039657692497e-05, 3.16039657692497e-05, 
    3.16039657692524e-05, 3.16039657692497e-05, 3.16039657692497e-05, 
    3.16039657692524e-05, 3.16039657692497e-05, 3.16039657692497e-05, 
    3.16039657692524e-05, 3.16039657692497e-05, 3.16039657692497e-05, 
    3.16039657692524e-05, 3.16039657692497e-05, 3.16039657692497e-05, 
    3.16039657692524e-05, 3.16039657692497e-05, 3.16039657692497e-05, 
    3.16039657692524e-05, 3.16039657692497e-05, 3.1603965769251e-05, 
    3.1603965769251e-05, 3.16039657692497e-05, 3.1603965769251e-05, 
    3.1603965769251e-05, 3.1603965769251e-05,
  3.17168397857176e-05, 3.17168397857176e-05, 3.17168397857176e-05, 
    3.17168397857122e-05, 3.17168397857176e-05, 3.17168397857176e-05, 
    3.17168397857122e-05, 3.17168397857176e-05, 3.17168397857176e-05, 
    3.17168397857122e-05, 3.17168397857176e-05, 3.17168397857176e-05, 
    3.17168397857122e-05, 3.17168397857176e-05, 3.17168397857176e-05, 
    3.17168397857122e-05, 3.17168397857176e-05, 3.17168397857176e-05, 
    3.17168397857149e-05, 3.17168397857149e-05, 3.17168397857149e-05, 
    3.17168397857176e-05, 3.17168397857149e-05, 3.17168397857149e-05, 
    3.17168397857176e-05, 3.17168397857149e-05, 3.17168397857149e-05, 
    3.17168397857176e-05, 3.17168397857149e-05, 3.17168397857149e-05, 
    3.17168397857176e-05, 3.17168397857149e-05, 3.17168397857149e-05, 
    3.17168397857176e-05, 3.17168397857149e-05, 3.17168397857149e-05, 
    3.17168397857176e-05, 3.17168397857149e-05, 3.17168397857149e-05, 
    3.17168397857176e-05, 3.17168397857149e-05, 3.17168397857149e-05, 
    3.17168397857176e-05, 3.17168397857149e-05, 3.17168397857149e-05, 
    3.17168397857176e-05, 3.17168397857149e-05, 3.17168397857149e-05, 
    3.17168397857176e-05, 3.17168397857149e-05, 3.17168397857162e-05, 
    3.17168397857162e-05, 3.17168397857149e-05, 3.17168397857162e-05, 
    3.17168397857162e-05, 3.17168397857162e-05,
  3.18316041973105e-05, 3.18316041973105e-05, 3.18316041973105e-05, 
    3.1831604197305e-05, 3.18316041973105e-05, 3.18316041973105e-05, 
    3.1831604197305e-05, 3.18316041973105e-05, 3.18316041973105e-05, 
    3.1831604197305e-05, 3.18316041973105e-05, 3.18316041973105e-05, 
    3.1831604197305e-05, 3.18316041973105e-05, 3.18316041973105e-05, 
    3.1831604197305e-05, 3.18316041973105e-05, 3.18316041973105e-05, 
    3.18316041973078e-05, 3.18316041973078e-05, 3.18316041973078e-05, 
    3.18316041973105e-05, 3.18316041973078e-05, 3.18316041973078e-05, 
    3.18316041973105e-05, 3.18316041973078e-05, 3.18316041973078e-05, 
    3.18316041973105e-05, 3.18316041973078e-05, 3.18316041973078e-05, 
    3.18316041973105e-05, 3.18316041973078e-05, 3.18316041973078e-05, 
    3.18316041973105e-05, 3.18316041973078e-05, 3.18316041973078e-05, 
    3.18316041973105e-05, 3.18316041973078e-05, 3.18316041973078e-05, 
    3.18316041973105e-05, 3.18316041973078e-05, 3.18316041973078e-05, 
    3.18316041973105e-05, 3.18316041973078e-05, 3.18316041973078e-05, 
    3.18316041973105e-05, 3.18316041973078e-05, 3.18316041973078e-05, 
    3.18316041973105e-05, 3.18316041973078e-05, 3.18316041973091e-05, 
    3.18316041973091e-05, 3.18316041973078e-05, 3.18316041973091e-05, 
    3.18316041973091e-05, 3.18316041973091e-05,
  3.19482874108883e-05, 3.19482874108883e-05, 3.19482874108883e-05, 
    3.19482874108828e-05, 3.19482874108883e-05, 3.19482874108883e-05, 
    3.19482874108828e-05, 3.19482874108883e-05, 3.19482874108883e-05, 
    3.19482874108828e-05, 3.19482874108883e-05, 3.19482874108883e-05, 
    3.19482874108828e-05, 3.19482874108883e-05, 3.19482874108883e-05, 
    3.19482874108828e-05, 3.19482874108883e-05, 3.19482874108883e-05, 
    3.19482874108856e-05, 3.19482874108856e-05, 3.19482874108856e-05, 
    3.19482874108883e-05, 3.19482874108856e-05, 3.19482874108856e-05, 
    3.19482874108883e-05, 3.19482874108856e-05, 3.19482874108856e-05, 
    3.19482874108883e-05, 3.19482874108856e-05, 3.19482874108856e-05, 
    3.19482874108883e-05, 3.19482874108856e-05, 3.19482874108856e-05, 
    3.19482874108883e-05, 3.19482874108856e-05, 3.19482874108856e-05, 
    3.19482874108883e-05, 3.19482874108856e-05, 3.19482874108856e-05, 
    3.19482874108883e-05, 3.19482874108856e-05, 3.19482874108856e-05, 
    3.19482874108883e-05, 3.19482874108856e-05, 3.19482874108856e-05, 
    3.19482874108883e-05, 3.19482874108856e-05, 3.19482874108856e-05, 
    3.19482874108883e-05, 3.19482874108856e-05, 3.19482874108869e-05, 
    3.19482874108869e-05, 3.19482874108856e-05, 3.19482874108869e-05, 
    3.19482874108869e-05, 3.19482874108869e-05,
  3.20669185478576e-05, 3.20669185478576e-05, 3.20669185478576e-05, 
    3.20669185478521e-05, 3.20669185478576e-05, 3.20669185478576e-05, 
    3.20669185478521e-05, 3.20669185478576e-05, 3.20669185478576e-05, 
    3.20669185478521e-05, 3.20669185478576e-05, 3.20669185478576e-05, 
    3.20669185478521e-05, 3.20669185478576e-05, 3.20669185478576e-05, 
    3.20669185478521e-05, 3.20669185478576e-05, 3.20669185478576e-05, 
    3.20669185478548e-05, 3.20669185478548e-05, 3.20669185478548e-05, 
    3.20669185478576e-05, 3.20669185478548e-05, 3.20669185478548e-05, 
    3.20669185478576e-05, 3.20669185478548e-05, 3.20669185478548e-05, 
    3.20669185478576e-05, 3.20669185478548e-05, 3.20669185478548e-05, 
    3.20669185478576e-05, 3.20669185478548e-05, 3.20669185478548e-05, 
    3.20669185478576e-05, 3.20669185478548e-05, 3.20669185478548e-05, 
    3.20669185478576e-05, 3.20669185478548e-05, 3.20669185478548e-05, 
    3.20669185478576e-05, 3.20669185478548e-05, 3.20669185478548e-05, 
    3.20669185478576e-05, 3.20669185478548e-05, 3.20669185478548e-05, 
    3.20669185478576e-05, 3.20669185478548e-05, 3.20669185478548e-05, 
    3.20669185478576e-05, 3.20669185478548e-05, 3.20669185478562e-05, 
    3.20669185478562e-05, 3.20669185478548e-05, 3.20669185478562e-05, 
    3.20669185478562e-05, 3.20669185478562e-05,
  3.21875274643601e-05, 3.21875274643601e-05, 3.21875274643601e-05, 
    3.21875274643546e-05, 3.21875274643601e-05, 3.21875274643601e-05, 
    3.21875274643546e-05, 3.21875274643601e-05, 3.21875274643601e-05, 
    3.21875274643546e-05, 3.21875274643601e-05, 3.21875274643601e-05, 
    3.21875274643546e-05, 3.21875274643601e-05, 3.21875274643601e-05, 
    3.21875274643546e-05, 3.21875274643601e-05, 3.21875274643601e-05, 
    3.21875274643573e-05, 3.21875274643573e-05, 3.21875274643573e-05, 
    3.21875274643601e-05, 3.21875274643573e-05, 3.21875274643573e-05, 
    3.21875274643601e-05, 3.21875274643573e-05, 3.21875274643573e-05, 
    3.21875274643601e-05, 3.21875274643573e-05, 3.21875274643573e-05, 
    3.21875274643601e-05, 3.21875274643573e-05, 3.21875274643573e-05, 
    3.21875274643601e-05, 3.21875274643573e-05, 3.21875274643573e-05, 
    3.21875274643601e-05, 3.21875274643573e-05, 3.21875274643573e-05, 
    3.21875274643601e-05, 3.21875274643573e-05, 3.21875274643573e-05, 
    3.21875274643601e-05, 3.21875274643573e-05, 3.21875274643573e-05, 
    3.21875274643601e-05, 3.21875274643573e-05, 3.21875274643573e-05, 
    3.21875274643601e-05, 3.21875274643573e-05, 3.21875274643587e-05, 
    3.21875274643587e-05, 3.21875274643573e-05, 3.21875274643587e-05, 
    3.21875274643587e-05, 3.21875274643587e-05,
  3.23101447721831e-05, 3.23101447721831e-05, 3.23101447721831e-05, 
    3.23101447721776e-05, 3.23101447721831e-05, 3.23101447721831e-05, 
    3.23101447721776e-05, 3.23101447721831e-05, 3.23101447721831e-05, 
    3.23101447721776e-05, 3.23101447721831e-05, 3.23101447721831e-05, 
    3.23101447721776e-05, 3.23101447721831e-05, 3.23101447721831e-05, 
    3.23101447721776e-05, 3.23101447721831e-05, 3.23101447721831e-05, 
    3.23101447721804e-05, 3.23101447721804e-05, 3.23101447721804e-05, 
    3.23101447721831e-05, 3.23101447721804e-05, 3.23101447721804e-05, 
    3.23101447721831e-05, 3.23101447721804e-05, 3.23101447721804e-05, 
    3.23101447721831e-05, 3.23101447721804e-05, 3.23101447721804e-05, 
    3.23101447721831e-05, 3.23101447721804e-05, 3.23101447721804e-05, 
    3.23101447721831e-05, 3.23101447721804e-05, 3.23101447721804e-05, 
    3.23101447721831e-05, 3.23101447721804e-05, 3.23101447721804e-05, 
    3.23101447721831e-05, 3.23101447721804e-05, 3.23101447721804e-05, 
    3.23101447721831e-05, 3.23101447721804e-05, 3.23101447721804e-05, 
    3.23101447721831e-05, 3.23101447721804e-05, 3.23101447721804e-05, 
    3.23101447721831e-05, 3.23101447721804e-05, 3.23101447721818e-05, 
    3.23101447721818e-05, 3.23101447721804e-05, 3.23101447721818e-05, 
    3.23101447721818e-05, 3.23101447721818e-05,
  3.24348018604244e-05, 3.24348018604244e-05, 3.24348018604244e-05, 
    3.24348018604188e-05, 3.24348018604244e-05, 3.24348018604244e-05, 
    3.24348018604188e-05, 3.24348018604244e-05, 3.24348018604244e-05, 
    3.24348018604188e-05, 3.24348018604244e-05, 3.24348018604244e-05, 
    3.24348018604188e-05, 3.24348018604244e-05, 3.24348018604244e-05, 
    3.24348018604188e-05, 3.24348018604244e-05, 3.24348018604244e-05, 
    3.24348018604216e-05, 3.24348018604216e-05, 3.24348018604216e-05, 
    3.24348018604244e-05, 3.24348018604216e-05, 3.24348018604216e-05, 
    3.24348018604244e-05, 3.24348018604216e-05, 3.24348018604216e-05, 
    3.24348018604244e-05, 3.24348018604216e-05, 3.24348018604216e-05, 
    3.24348018604244e-05, 3.24348018604216e-05, 3.24348018604216e-05, 
    3.24348018604244e-05, 3.24348018604216e-05, 3.24348018604216e-05, 
    3.24348018604244e-05, 3.24348018604216e-05, 3.24348018604216e-05, 
    3.24348018604244e-05, 3.24348018604216e-05, 3.24348018604216e-05, 
    3.24348018604244e-05, 3.24348018604216e-05, 3.24348018604216e-05, 
    3.24348018604244e-05, 3.24348018604216e-05, 3.24348018604216e-05, 
    3.24348018604244e-05, 3.24348018604216e-05, 3.2434801860423e-05, 
    3.2434801860423e-05, 3.24348018604216e-05, 3.2434801860423e-05, 
    3.2434801860423e-05, 3.2434801860423e-05,
  3.25615309179415e-05, 3.25615309179415e-05, 3.25615309179415e-05, 
    3.25615309179359e-05, 3.25615309179415e-05, 3.25615309179415e-05, 
    3.25615309179359e-05, 3.25615309179415e-05, 3.25615309179415e-05, 
    3.25615309179359e-05, 3.25615309179415e-05, 3.25615309179415e-05, 
    3.25615309179359e-05, 3.25615309179415e-05, 3.25615309179415e-05, 
    3.25615309179359e-05, 3.25615309179415e-05, 3.25615309179415e-05, 
    3.25615309179387e-05, 3.25615309179387e-05, 3.25615309179387e-05, 
    3.25615309179415e-05, 3.25615309179387e-05, 3.25615309179387e-05, 
    3.25615309179415e-05, 3.25615309179387e-05, 3.25615309179387e-05, 
    3.25615309179415e-05, 3.25615309179387e-05, 3.25615309179387e-05, 
    3.25615309179415e-05, 3.25615309179387e-05, 3.25615309179387e-05, 
    3.25615309179415e-05, 3.25615309179387e-05, 3.25615309179387e-05, 
    3.25615309179415e-05, 3.25615309179387e-05, 3.25615309179387e-05, 
    3.25615309179415e-05, 3.25615309179387e-05, 3.25615309179387e-05, 
    3.25615309179415e-05, 3.25615309179387e-05, 3.25615309179387e-05, 
    3.25615309179415e-05, 3.25615309179387e-05, 3.25615309179387e-05, 
    3.25615309179415e-05, 3.25615309179387e-05, 3.25615309179401e-05, 
    3.25615309179401e-05, 3.25615309179387e-05, 3.25615309179401e-05, 
    3.25615309179401e-05, 3.25615309179401e-05,
  3.26903649566202e-05, 3.26903649566202e-05, 3.26903649566202e-05, 
    3.26903649566147e-05, 3.26903649566202e-05, 3.26903649566202e-05, 
    3.26903649566147e-05, 3.26903649566202e-05, 3.26903649566202e-05, 
    3.26903649566147e-05, 3.26903649566202e-05, 3.26903649566202e-05, 
    3.26903649566147e-05, 3.26903649566202e-05, 3.26903649566202e-05, 
    3.26903649566147e-05, 3.26903649566202e-05, 3.26903649566202e-05, 
    3.26903649566174e-05, 3.26903649566174e-05, 3.26903649566174e-05, 
    3.26903649566202e-05, 3.26903649566174e-05, 3.26903649566174e-05, 
    3.26903649566202e-05, 3.26903649566174e-05, 3.26903649566174e-05, 
    3.26903649566202e-05, 3.26903649566174e-05, 3.26903649566174e-05, 
    3.26903649566202e-05, 3.26903649566174e-05, 3.26903649566174e-05, 
    3.26903649566202e-05, 3.26903649566174e-05, 3.26903649566174e-05, 
    3.26903649566202e-05, 3.26903649566174e-05, 3.26903649566174e-05, 
    3.26903649566202e-05, 3.26903649566174e-05, 3.26903649566174e-05, 
    3.26903649566202e-05, 3.26903649566174e-05, 3.26903649566174e-05, 
    3.26903649566202e-05, 3.26903649566174e-05, 3.26903649566174e-05, 
    3.26903649566202e-05, 3.26903649566174e-05, 3.26903649566188e-05, 
    3.26903649566188e-05, 3.26903649566174e-05, 3.26903649566188e-05, 
    3.26903649566188e-05, 3.26903649566188e-05,
  3.28213378354946e-05, 3.28213378354946e-05, 3.28213378354946e-05, 
    3.2821337835489e-05, 3.28213378354946e-05, 3.28213378354946e-05, 
    3.2821337835489e-05, 3.28213378354946e-05, 3.28213378354946e-05, 
    3.2821337835489e-05, 3.28213378354946e-05, 3.28213378354946e-05, 
    3.2821337835489e-05, 3.28213378354946e-05, 3.28213378354946e-05, 
    3.2821337835489e-05, 3.28213378354946e-05, 3.28213378354946e-05, 
    3.28213378354918e-05, 3.28213378354918e-05, 3.28213378354918e-05, 
    3.28213378354946e-05, 3.28213378354918e-05, 3.28213378354918e-05, 
    3.28213378354946e-05, 3.28213378354918e-05, 3.28213378354918e-05, 
    3.28213378354946e-05, 3.28213378354918e-05, 3.28213378354918e-05, 
    3.28213378354946e-05, 3.28213378354918e-05, 3.28213378354918e-05, 
    3.28213378354946e-05, 3.28213378354918e-05, 3.28213378354918e-05, 
    3.28213378354946e-05, 3.28213378354918e-05, 3.28213378354918e-05, 
    3.28213378354946e-05, 3.28213378354918e-05, 3.28213378354918e-05, 
    3.28213378354946e-05, 3.28213378354918e-05, 3.28213378354918e-05, 
    3.28213378354946e-05, 3.28213378354918e-05, 3.28213378354918e-05, 
    3.28213378354946e-05, 3.28213378354918e-05, 3.28213378354932e-05, 
    3.28213378354932e-05, 3.28213378354918e-05, 3.28213378354932e-05, 
    3.28213378354932e-05, 3.28213378354932e-05,
  3.29544842857554e-05, 3.29544842857554e-05, 3.29544842857554e-05, 
    3.29544842857498e-05, 3.29544842857554e-05, 3.29544842857554e-05, 
    3.29544842857498e-05, 3.29544842857554e-05, 3.29544842857554e-05, 
    3.29544842857498e-05, 3.29544842857554e-05, 3.29544842857554e-05, 
    3.29544842857498e-05, 3.29544842857554e-05, 3.29544842857554e-05, 
    3.29544842857498e-05, 3.29544842857554e-05, 3.29544842857554e-05, 
    3.29544842857526e-05, 3.29544842857526e-05, 3.29544842857526e-05, 
    3.29544842857554e-05, 3.29544842857526e-05, 3.29544842857526e-05, 
    3.29544842857554e-05, 3.29544842857526e-05, 3.29544842857526e-05, 
    3.29544842857554e-05, 3.29544842857526e-05, 3.29544842857526e-05, 
    3.29544842857554e-05, 3.29544842857526e-05, 3.29544842857526e-05, 
    3.29544842857554e-05, 3.29544842857526e-05, 3.29544842857526e-05, 
    3.29544842857554e-05, 3.29544842857526e-05, 3.29544842857526e-05, 
    3.29544842857554e-05, 3.29544842857526e-05, 3.29544842857526e-05, 
    3.29544842857554e-05, 3.29544842857526e-05, 3.29544842857526e-05, 
    3.29544842857554e-05, 3.29544842857526e-05, 3.29544842857526e-05, 
    3.29544842857554e-05, 3.29544842857526e-05, 3.2954484285754e-05, 
    3.2954484285754e-05, 3.29544842857526e-05, 3.2954484285754e-05, 
    3.2954484285754e-05, 3.2954484285754e-05,
  3.30898399366848e-05, 3.30898399366848e-05, 3.30898399366848e-05, 
    3.30898399366792e-05, 3.30898399366848e-05, 3.30898399366848e-05, 
    3.30898399366792e-05, 3.30898399366848e-05, 3.30898399366848e-05, 
    3.30898399366792e-05, 3.30898399366848e-05, 3.30898399366848e-05, 
    3.30898399366792e-05, 3.30898399366848e-05, 3.30898399366848e-05, 
    3.30898399366792e-05, 3.30898399366848e-05, 3.30898399366848e-05, 
    3.3089839936682e-05, 3.3089839936682e-05, 3.3089839936682e-05, 
    3.30898399366848e-05, 3.3089839936682e-05, 3.3089839936682e-05, 
    3.30898399366848e-05, 3.3089839936682e-05, 3.3089839936682e-05, 
    3.30898399366848e-05, 3.3089839936682e-05, 3.3089839936682e-05, 
    3.30898399366848e-05, 3.3089839936682e-05, 3.3089839936682e-05, 
    3.30898399366848e-05, 3.3089839936682e-05, 3.3089839936682e-05, 
    3.30898399366848e-05, 3.3089839936682e-05, 3.3089839936682e-05, 
    3.30898399366848e-05, 3.3089839936682e-05, 3.3089839936682e-05, 
    3.30898399366848e-05, 3.3089839936682e-05, 3.3089839936682e-05, 
    3.30898399366848e-05, 3.3089839936682e-05, 3.3089839936682e-05, 
    3.30898399366848e-05, 3.3089839936682e-05, 3.30898399366834e-05, 
    3.30898399366834e-05, 3.3089839936682e-05, 3.30898399366834e-05, 
    3.30898399366834e-05, 3.30898399366834e-05,
  3.32274413425564e-05, 3.32274413425564e-05, 3.32274413425564e-05, 
    3.32274413425507e-05, 3.32274413425564e-05, 3.32274413425564e-05, 
    3.32274413425507e-05, 3.32274413425564e-05, 3.32274413425564e-05, 
    3.32274413425507e-05, 3.32274413425564e-05, 3.32274413425564e-05, 
    3.32274413425507e-05, 3.32274413425564e-05, 3.32274413425564e-05, 
    3.32274413425507e-05, 3.32274413425564e-05, 3.32274413425564e-05, 
    3.32274413425535e-05, 3.32274413425535e-05, 3.32274413425535e-05, 
    3.32274413425564e-05, 3.32274413425535e-05, 3.32274413425535e-05, 
    3.32274413425564e-05, 3.32274413425535e-05, 3.32274413425535e-05, 
    3.32274413425564e-05, 3.32274413425535e-05, 3.32274413425535e-05, 
    3.32274413425564e-05, 3.32274413425535e-05, 3.32274413425535e-05, 
    3.32274413425564e-05, 3.32274413425535e-05, 3.32274413425535e-05, 
    3.32274413425564e-05, 3.32274413425535e-05, 3.32274413425535e-05, 
    3.32274413425564e-05, 3.32274413425535e-05, 3.32274413425535e-05, 
    3.32274413425564e-05, 3.32274413425535e-05, 3.32274413425535e-05, 
    3.32274413425564e-05, 3.32274413425535e-05, 3.32274413425535e-05, 
    3.32274413425564e-05, 3.32274413425535e-05, 3.3227441342555e-05, 
    3.3227441342555e-05, 3.32274413425535e-05, 3.3227441342555e-05, 
    3.3227441342555e-05, 3.3227441342555e-05,
  3.33673260105419e-05, 3.33673260105419e-05, 3.33673260105419e-05, 
    3.33673260105362e-05, 3.33673260105419e-05, 3.33673260105419e-05, 
    3.33673260105362e-05, 3.33673260105419e-05, 3.33673260105419e-05, 
    3.33673260105362e-05, 3.33673260105419e-05, 3.33673260105419e-05, 
    3.33673260105362e-05, 3.33673260105419e-05, 3.33673260105419e-05, 
    3.33673260105362e-05, 3.33673260105419e-05, 3.33673260105419e-05, 
    3.33673260105391e-05, 3.33673260105391e-05, 3.33673260105391e-05, 
    3.33673260105419e-05, 3.33673260105391e-05, 3.33673260105391e-05, 
    3.33673260105419e-05, 3.33673260105391e-05, 3.33673260105391e-05, 
    3.33673260105419e-05, 3.33673260105391e-05, 3.33673260105391e-05, 
    3.33673260105419e-05, 3.33673260105391e-05, 3.33673260105391e-05, 
    3.33673260105419e-05, 3.33673260105391e-05, 3.33673260105391e-05, 
    3.33673260105419e-05, 3.33673260105391e-05, 3.33673260105391e-05, 
    3.33673260105419e-05, 3.33673260105391e-05, 3.33673260105391e-05, 
    3.33673260105419e-05, 3.33673260105391e-05, 3.33673260105391e-05, 
    3.33673260105419e-05, 3.33673260105391e-05, 3.33673260105391e-05, 
    3.33673260105419e-05, 3.33673260105391e-05, 3.33673260105405e-05, 
    3.33673260105405e-05, 3.33673260105391e-05, 3.33673260105405e-05, 
    3.33673260105405e-05, 3.33673260105405e-05,
  3.35095324296697e-05, 3.35095324296697e-05, 3.35095324296697e-05, 
    3.3509532429664e-05, 3.35095324296697e-05, 3.35095324296697e-05, 
    3.3509532429664e-05, 3.35095324296697e-05, 3.35095324296697e-05, 
    3.3509532429664e-05, 3.35095324296697e-05, 3.35095324296697e-05, 
    3.3509532429664e-05, 3.35095324296697e-05, 3.35095324296697e-05, 
    3.3509532429664e-05, 3.35095324296697e-05, 3.35095324296697e-05, 
    3.35095324296669e-05, 3.35095324296669e-05, 3.35095324296669e-05, 
    3.35095324296697e-05, 3.35095324296669e-05, 3.35095324296669e-05, 
    3.35095324296697e-05, 3.35095324296669e-05, 3.35095324296669e-05, 
    3.35095324296697e-05, 3.35095324296669e-05, 3.35095324296669e-05, 
    3.35095324296697e-05, 3.35095324296669e-05, 3.35095324296669e-05, 
    3.35095324296697e-05, 3.35095324296669e-05, 3.35095324296669e-05, 
    3.35095324296697e-05, 3.35095324296669e-05, 3.35095324296669e-05, 
    3.35095324296697e-05, 3.35095324296669e-05, 3.35095324296669e-05, 
    3.35095324296697e-05, 3.35095324296669e-05, 3.35095324296669e-05, 
    3.35095324296697e-05, 3.35095324296669e-05, 3.35095324296669e-05, 
    3.35095324296697e-05, 3.35095324296669e-05, 3.35095324296683e-05, 
    3.35095324296683e-05, 3.35095324296669e-05, 3.35095324296683e-05, 
    3.35095324296683e-05, 3.35095324296683e-05,
  3.36541001008783e-05, 3.36541001008783e-05, 3.36541001008783e-05, 
    3.36541001008726e-05, 3.36541001008783e-05, 3.36541001008783e-05, 
    3.36541001008726e-05, 3.36541001008783e-05, 3.36541001008783e-05, 
    3.36541001008726e-05, 3.36541001008783e-05, 3.36541001008783e-05, 
    3.36541001008726e-05, 3.36541001008783e-05, 3.36541001008783e-05, 
    3.36541001008726e-05, 3.36541001008783e-05, 3.36541001008783e-05, 
    3.36541001008754e-05, 3.36541001008754e-05, 3.36541001008754e-05, 
    3.36541001008783e-05, 3.36541001008754e-05, 3.36541001008754e-05, 
    3.36541001008783e-05, 3.36541001008754e-05, 3.36541001008754e-05, 
    3.36541001008783e-05, 3.36541001008754e-05, 3.36541001008754e-05, 
    3.36541001008783e-05, 3.36541001008754e-05, 3.36541001008754e-05, 
    3.36541001008783e-05, 3.36541001008754e-05, 3.36541001008754e-05, 
    3.36541001008783e-05, 3.36541001008754e-05, 3.36541001008754e-05, 
    3.36541001008783e-05, 3.36541001008754e-05, 3.36541001008754e-05, 
    3.36541001008783e-05, 3.36541001008754e-05, 3.36541001008754e-05, 
    3.36541001008783e-05, 3.36541001008754e-05, 3.36541001008754e-05, 
    3.36541001008783e-05, 3.36541001008754e-05, 3.36541001008769e-05, 
    3.36541001008769e-05, 3.36541001008754e-05, 3.36541001008769e-05, 
    3.36541001008769e-05, 3.36541001008769e-05,
  3.38010695682153e-05, 3.38010695682153e-05, 3.38010695682153e-05, 
    3.38010695682095e-05, 3.38010695682153e-05, 3.38010695682153e-05, 
    3.38010695682095e-05, 3.38010695682153e-05, 3.38010695682153e-05, 
    3.38010695682095e-05, 3.38010695682153e-05, 3.38010695682153e-05, 
    3.38010695682095e-05, 3.38010695682153e-05, 3.38010695682153e-05, 
    3.38010695682095e-05, 3.38010695682153e-05, 3.38010695682153e-05, 
    3.38010695682124e-05, 3.38010695682124e-05, 3.38010695682124e-05, 
    3.38010695682153e-05, 3.38010695682124e-05, 3.38010695682124e-05, 
    3.38010695682153e-05, 3.38010695682124e-05, 3.38010695682124e-05, 
    3.38010695682153e-05, 3.38010695682124e-05, 3.38010695682124e-05, 
    3.38010695682153e-05, 3.38010695682124e-05, 3.38010695682124e-05, 
    3.38010695682153e-05, 3.38010695682124e-05, 3.38010695682124e-05, 
    3.38010695682153e-05, 3.38010695682124e-05, 3.38010695682124e-05, 
    3.38010695682153e-05, 3.38010695682124e-05, 3.38010695682124e-05, 
    3.38010695682153e-05, 3.38010695682124e-05, 3.38010695682124e-05, 
    3.38010695682153e-05, 3.38010695682124e-05, 3.38010695682124e-05, 
    3.38010695682153e-05, 3.38010695682124e-05, 3.38010695682139e-05, 
    3.38010695682139e-05, 3.38010695682124e-05, 3.38010695682139e-05, 
    3.38010695682139e-05, 3.38010695682139e-05,
  3.39504824512312e-05, 3.39504824512312e-05, 3.39504824512312e-05, 
    3.39504824512254e-05, 3.39504824512312e-05, 3.39504824512312e-05, 
    3.39504824512254e-05, 3.39504824512312e-05, 3.39504824512312e-05, 
    3.39504824512254e-05, 3.39504824512312e-05, 3.39504824512312e-05, 
    3.39504824512254e-05, 3.39504824512312e-05, 3.39504824512312e-05, 
    3.39504824512254e-05, 3.39504824512312e-05, 3.39504824512312e-05, 
    3.39504824512283e-05, 3.39504824512283e-05, 3.39504824512283e-05, 
    3.39504824512312e-05, 3.39504824512283e-05, 3.39504824512283e-05, 
    3.39504824512312e-05, 3.39504824512283e-05, 3.39504824512283e-05, 
    3.39504824512312e-05, 3.39504824512283e-05, 3.39504824512283e-05, 
    3.39504824512312e-05, 3.39504824512283e-05, 3.39504824512283e-05, 
    3.39504824512312e-05, 3.39504824512283e-05, 3.39504824512283e-05, 
    3.39504824512312e-05, 3.39504824512283e-05, 3.39504824512283e-05, 
    3.39504824512312e-05, 3.39504824512283e-05, 3.39504824512283e-05, 
    3.39504824512312e-05, 3.39504824512283e-05, 3.39504824512283e-05, 
    3.39504824512312e-05, 3.39504824512283e-05, 3.39504824512283e-05, 
    3.39504824512312e-05, 3.39504824512283e-05, 3.39504824512297e-05, 
    3.39504824512297e-05, 3.39504824512283e-05, 3.39504824512297e-05, 
    3.39504824512297e-05, 3.39504824512297e-05,
  3.4102381478621e-05, 3.4102381478621e-05, 3.4102381478621e-05, 
    3.41023814786152e-05, 3.4102381478621e-05, 3.4102381478621e-05, 
    3.41023814786152e-05, 3.4102381478621e-05, 3.4102381478621e-05, 
    3.41023814786152e-05, 3.4102381478621e-05, 3.4102381478621e-05, 
    3.41023814786152e-05, 3.4102381478621e-05, 3.4102381478621e-05, 
    3.41023814786152e-05, 3.4102381478621e-05, 3.4102381478621e-05, 
    3.41023814786181e-05, 3.41023814786181e-05, 3.41023814786181e-05, 
    3.4102381478621e-05, 3.41023814786181e-05, 3.41023814786181e-05, 
    3.4102381478621e-05, 3.41023814786181e-05, 3.41023814786181e-05, 
    3.4102381478621e-05, 3.41023814786181e-05, 3.41023814786181e-05, 
    3.4102381478621e-05, 3.41023814786181e-05, 3.41023814786181e-05, 
    3.4102381478621e-05, 3.41023814786181e-05, 3.41023814786181e-05, 
    3.4102381478621e-05, 3.41023814786181e-05, 3.41023814786181e-05, 
    3.4102381478621e-05, 3.41023814786181e-05, 3.41023814786181e-05, 
    3.4102381478621e-05, 3.41023814786181e-05, 3.41023814786181e-05, 
    3.4102381478621e-05, 3.41023814786181e-05, 3.41023814786181e-05, 
    3.4102381478621e-05, 3.41023814786181e-05, 3.41023814786196e-05, 
    3.41023814786196e-05, 3.41023814786181e-05, 3.41023814786196e-05, 
    3.41023814786196e-05, 3.41023814786196e-05,
  3.42568105231701e-05, 3.42568105231701e-05, 3.42568105231701e-05, 
    3.42568105231643e-05, 3.42568105231701e-05, 3.42568105231701e-05, 
    3.42568105231643e-05, 3.42568105231701e-05, 3.42568105231701e-05, 
    3.42568105231643e-05, 3.42568105231701e-05, 3.42568105231701e-05, 
    3.42568105231643e-05, 3.42568105231701e-05, 3.42568105231701e-05, 
    3.42568105231643e-05, 3.42568105231701e-05, 3.42568105231701e-05, 
    3.42568105231672e-05, 3.42568105231672e-05, 3.42568105231672e-05, 
    3.42568105231701e-05, 3.42568105231672e-05, 3.42568105231672e-05, 
    3.42568105231701e-05, 3.42568105231672e-05, 3.42568105231672e-05, 
    3.42568105231701e-05, 3.42568105231672e-05, 3.42568105231672e-05, 
    3.42568105231701e-05, 3.42568105231672e-05, 3.42568105231672e-05, 
    3.42568105231701e-05, 3.42568105231672e-05, 3.42568105231672e-05, 
    3.42568105231701e-05, 3.42568105231672e-05, 3.42568105231672e-05, 
    3.42568105231701e-05, 3.42568105231672e-05, 3.42568105231672e-05, 
    3.42568105231701e-05, 3.42568105231672e-05, 3.42568105231672e-05, 
    3.42568105231701e-05, 3.42568105231672e-05, 3.42568105231672e-05, 
    3.42568105231701e-05, 3.42568105231672e-05, 3.42568105231687e-05, 
    3.42568105231687e-05, 3.42568105231672e-05, 3.42568105231687e-05, 
    3.42568105231687e-05, 3.42568105231687e-05,
  3.44138146380627e-05, 3.44138146380627e-05, 3.44138146380627e-05, 
    3.44138146380568e-05, 3.44138146380627e-05, 3.44138146380627e-05, 
    3.44138146380568e-05, 3.44138146380627e-05, 3.44138146380627e-05, 
    3.44138146380568e-05, 3.44138146380627e-05, 3.44138146380627e-05, 
    3.44138146380568e-05, 3.44138146380627e-05, 3.44138146380627e-05, 
    3.44138146380568e-05, 3.44138146380627e-05, 3.44138146380627e-05, 
    3.44138146380598e-05, 3.44138146380598e-05, 3.44138146380598e-05, 
    3.44138146380627e-05, 3.44138146380598e-05, 3.44138146380598e-05, 
    3.44138146380627e-05, 3.44138146380598e-05, 3.44138146380598e-05, 
    3.44138146380627e-05, 3.44138146380598e-05, 3.44138146380598e-05, 
    3.44138146380627e-05, 3.44138146380598e-05, 3.44138146380598e-05, 
    3.44138146380627e-05, 3.44138146380598e-05, 3.44138146380598e-05, 
    3.44138146380627e-05, 3.44138146380598e-05, 3.44138146380598e-05, 
    3.44138146380627e-05, 3.44138146380598e-05, 3.44138146380598e-05, 
    3.44138146380627e-05, 3.44138146380598e-05, 3.44138146380598e-05, 
    3.44138146380627e-05, 3.44138146380598e-05, 3.44138146380598e-05, 
    3.44138146380627e-05, 3.44138146380598e-05, 3.44138146380612e-05, 
    3.44138146380612e-05, 3.44138146380598e-05, 3.44138146380612e-05, 
    3.44138146380612e-05, 3.44138146380612e-05,
  3.45734400946144e-05, 3.45734400946144e-05, 3.45734400946144e-05, 
    3.45734400946086e-05, 3.45734400946144e-05, 3.45734400946144e-05, 
    3.45734400946086e-05, 3.45734400946144e-05, 3.45734400946144e-05, 
    3.45734400946086e-05, 3.45734400946144e-05, 3.45734400946144e-05, 
    3.45734400946086e-05, 3.45734400946144e-05, 3.45734400946144e-05, 
    3.45734400946086e-05, 3.45734400946144e-05, 3.45734400946144e-05, 
    3.45734400946115e-05, 3.45734400946115e-05, 3.45734400946115e-05, 
    3.45734400946144e-05, 3.45734400946115e-05, 3.45734400946115e-05, 
    3.45734400946144e-05, 3.45734400946115e-05, 3.45734400946115e-05, 
    3.45734400946144e-05, 3.45734400946115e-05, 3.45734400946115e-05, 
    3.45734400946144e-05, 3.45734400946115e-05, 3.45734400946115e-05, 
    3.45734400946144e-05, 3.45734400946115e-05, 3.45734400946115e-05, 
    3.45734400946144e-05, 3.45734400946115e-05, 3.45734400946115e-05, 
    3.45734400946144e-05, 3.45734400946115e-05, 3.45734400946115e-05, 
    3.45734400946144e-05, 3.45734400946115e-05, 3.45734400946115e-05, 
    3.45734400946144e-05, 3.45734400946115e-05, 3.45734400946115e-05, 
    3.45734400946144e-05, 3.45734400946115e-05, 3.4573440094613e-05, 
    3.4573440094613e-05, 3.45734400946115e-05, 3.4573440094613e-05, 
    3.4573440094613e-05, 3.4573440094613e-05,
  3.47357344214949e-05, 3.47357344214949e-05, 3.47357344214949e-05, 
    3.4735734421489e-05, 3.47357344214949e-05, 3.47357344214949e-05, 
    3.4735734421489e-05, 3.47357344214949e-05, 3.47357344214949e-05, 
    3.4735734421489e-05, 3.47357344214949e-05, 3.47357344214949e-05, 
    3.4735734421489e-05, 3.47357344214949e-05, 3.47357344214949e-05, 
    3.4735734421489e-05, 3.47357344214949e-05, 3.47357344214949e-05, 
    3.47357344214919e-05, 3.47357344214919e-05, 3.47357344214919e-05, 
    3.47357344214949e-05, 3.47357344214919e-05, 3.47357344214919e-05, 
    3.47357344214949e-05, 3.47357344214919e-05, 3.47357344214919e-05, 
    3.47357344214949e-05, 3.47357344214919e-05, 3.47357344214919e-05, 
    3.47357344214949e-05, 3.47357344214919e-05, 3.47357344214919e-05, 
    3.47357344214949e-05, 3.47357344214919e-05, 3.47357344214919e-05, 
    3.47357344214949e-05, 3.47357344214919e-05, 3.47357344214919e-05, 
    3.47357344214949e-05, 3.47357344214919e-05, 3.47357344214919e-05, 
    3.47357344214949e-05, 3.47357344214919e-05, 3.47357344214919e-05, 
    3.47357344214949e-05, 3.47357344214919e-05, 3.47357344214919e-05, 
    3.47357344214949e-05, 3.47357344214919e-05, 3.47357344214934e-05, 
    3.47357344214934e-05, 3.47357344214919e-05, 3.47357344214934e-05, 
    3.47357344214934e-05, 3.47357344214934e-05,
  3.49007464455074e-05, 3.49007464455074e-05, 3.49007464455074e-05, 
    3.49007464455014e-05, 3.49007464455074e-05, 3.49007464455074e-05, 
    3.49007464455014e-05, 3.49007464455074e-05, 3.49007464455074e-05, 
    3.49007464455014e-05, 3.49007464455074e-05, 3.49007464455074e-05, 
    3.49007464455014e-05, 3.49007464455074e-05, 3.49007464455074e-05, 
    3.49007464455014e-05, 3.49007464455074e-05, 3.49007464455074e-05, 
    3.49007464455044e-05, 3.49007464455044e-05, 3.49007464455044e-05, 
    3.49007464455074e-05, 3.49007464455044e-05, 3.49007464455044e-05, 
    3.49007464455074e-05, 3.49007464455044e-05, 3.49007464455044e-05, 
    3.49007464455074e-05, 3.49007464455044e-05, 3.49007464455044e-05, 
    3.49007464455074e-05, 3.49007464455044e-05, 3.49007464455044e-05, 
    3.49007464455074e-05, 3.49007464455044e-05, 3.49007464455044e-05, 
    3.49007464455074e-05, 3.49007464455044e-05, 3.49007464455044e-05, 
    3.49007464455074e-05, 3.49007464455044e-05, 3.49007464455044e-05, 
    3.49007464455074e-05, 3.49007464455044e-05, 3.49007464455044e-05, 
    3.49007464455074e-05, 3.49007464455044e-05, 3.49007464455044e-05, 
    3.49007464455074e-05, 3.49007464455044e-05, 3.49007464455059e-05, 
    3.49007464455059e-05, 3.49007464455044e-05, 3.49007464455059e-05, 
    3.49007464455059e-05, 3.49007464455059e-05,
  3.50685263339989e-05, 3.50685263339989e-05, 3.50685263339989e-05, 
    3.50685263339929e-05, 3.50685263339989e-05, 3.50685263339989e-05, 
    3.50685263339929e-05, 3.50685263339989e-05, 3.50685263339989e-05, 
    3.50685263339929e-05, 3.50685263339989e-05, 3.50685263339989e-05, 
    3.50685263339929e-05, 3.50685263339989e-05, 3.50685263339989e-05, 
    3.50685263339929e-05, 3.50685263339989e-05, 3.50685263339989e-05, 
    3.50685263339959e-05, 3.50685263339959e-05, 3.50685263339959e-05, 
    3.50685263339989e-05, 3.50685263339959e-05, 3.50685263339959e-05, 
    3.50685263339989e-05, 3.50685263339959e-05, 3.50685263339959e-05, 
    3.50685263339989e-05, 3.50685263339959e-05, 3.50685263339959e-05, 
    3.50685263339989e-05, 3.50685263339959e-05, 3.50685263339959e-05, 
    3.50685263339989e-05, 3.50685263339959e-05, 3.50685263339959e-05, 
    3.50685263339989e-05, 3.50685263339959e-05, 3.50685263339959e-05, 
    3.50685263339989e-05, 3.50685263339959e-05, 3.50685263339959e-05, 
    3.50685263339989e-05, 3.50685263339959e-05, 3.50685263339959e-05, 
    3.50685263339989e-05, 3.50685263339959e-05, 3.50685263339959e-05, 
    3.50685263339989e-05, 3.50685263339959e-05, 3.50685263339974e-05, 
    3.50685263339974e-05, 3.50685263339959e-05, 3.50685263339974e-05, 
    3.50685263339974e-05, 3.50685263339974e-05,
  3.52391256389759e-05, 3.52391256389759e-05, 3.52391256389759e-05, 
    3.52391256389699e-05, 3.52391256389759e-05, 3.52391256389759e-05, 
    3.52391256389699e-05, 3.52391256389759e-05, 3.52391256389759e-05, 
    3.52391256389699e-05, 3.52391256389759e-05, 3.52391256389759e-05, 
    3.52391256389699e-05, 3.52391256389759e-05, 3.52391256389759e-05, 
    3.52391256389699e-05, 3.52391256389759e-05, 3.52391256389759e-05, 
    3.52391256389729e-05, 3.52391256389729e-05, 3.52391256389729e-05, 
    3.52391256389759e-05, 3.52391256389729e-05, 3.52391256389729e-05, 
    3.52391256389759e-05, 3.52391256389729e-05, 3.52391256389729e-05, 
    3.52391256389759e-05, 3.52391256389729e-05, 3.52391256389729e-05, 
    3.52391256389759e-05, 3.52391256389729e-05, 3.52391256389729e-05, 
    3.52391256389759e-05, 3.52391256389729e-05, 3.52391256389729e-05, 
    3.52391256389759e-05, 3.52391256389729e-05, 3.52391256389729e-05, 
    3.52391256389759e-05, 3.52391256389729e-05, 3.52391256389729e-05, 
    3.52391256389759e-05, 3.52391256389729e-05, 3.52391256389729e-05, 
    3.52391256389759e-05, 3.52391256389729e-05, 3.52391256389729e-05, 
    3.52391256389759e-05, 3.52391256389729e-05, 3.52391256389744e-05, 
    3.52391256389744e-05, 3.52391256389729e-05, 3.52391256389744e-05, 
    3.52391256389744e-05, 3.52391256389744e-05,
  3.54125973430055e-05, 3.54125973430055e-05, 3.54125973430055e-05, 
    3.54125973429995e-05, 3.54125973430055e-05, 3.54125973430055e-05, 
    3.54125973429995e-05, 3.54125973430055e-05, 3.54125973430055e-05, 
    3.54125973429995e-05, 3.54125973430055e-05, 3.54125973430055e-05, 
    3.54125973429995e-05, 3.54125973430055e-05, 3.54125973430055e-05, 
    3.54125973429995e-05, 3.54125973430055e-05, 3.54125973430055e-05, 
    3.54125973430025e-05, 3.54125973430025e-05, 3.54125973430025e-05, 
    3.54125973430055e-05, 3.54125973430025e-05, 3.54125973430025e-05, 
    3.54125973430055e-05, 3.54125973430025e-05, 3.54125973430025e-05, 
    3.54125973430055e-05, 3.54125973430025e-05, 3.54125973430025e-05, 
    3.54125973430055e-05, 3.54125973430025e-05, 3.54125973430025e-05, 
    3.54125973430055e-05, 3.54125973430025e-05, 3.54125973430025e-05, 
    3.54125973430055e-05, 3.54125973430025e-05, 3.54125973430025e-05, 
    3.54125973430055e-05, 3.54125973430025e-05, 3.54125973430025e-05, 
    3.54125973430055e-05, 3.54125973430025e-05, 3.54125973430025e-05, 
    3.54125973430055e-05, 3.54125973430025e-05, 3.54125973430025e-05, 
    3.54125973430055e-05, 3.54125973430025e-05, 3.5412597343004e-05, 
    3.5412597343004e-05, 3.54125973430025e-05, 3.5412597343004e-05, 
    3.5412597343004e-05, 3.5412597343004e-05,
  3.55889959069871e-05, 3.55889959069871e-05, 3.55889959069871e-05, 
    3.5588995906981e-05, 3.55889959069871e-05, 3.55889959069871e-05, 
    3.5588995906981e-05, 3.55889959069871e-05, 3.55889959069871e-05, 
    3.5588995906981e-05, 3.55889959069871e-05, 3.55889959069871e-05, 
    3.5588995906981e-05, 3.55889959069871e-05, 3.55889959069871e-05, 
    3.5588995906981e-05, 3.55889959069871e-05, 3.55889959069871e-05, 
    3.55889959069841e-05, 3.55889959069841e-05, 3.55889959069841e-05, 
    3.55889959069871e-05, 3.55889959069841e-05, 3.55889959069841e-05, 
    3.55889959069871e-05, 3.55889959069841e-05, 3.55889959069841e-05, 
    3.55889959069871e-05, 3.55889959069841e-05, 3.55889959069841e-05, 
    3.55889959069871e-05, 3.55889959069841e-05, 3.55889959069841e-05, 
    3.55889959069871e-05, 3.55889959069841e-05, 3.55889959069841e-05, 
    3.55889959069871e-05, 3.55889959069841e-05, 3.55889959069841e-05, 
    3.55889959069871e-05, 3.55889959069841e-05, 3.55889959069841e-05, 
    3.55889959069871e-05, 3.55889959069841e-05, 3.55889959069841e-05, 
    3.55889959069871e-05, 3.55889959069841e-05, 3.55889959069841e-05, 
    3.55889959069871e-05, 3.55889959069841e-05, 3.55889959069856e-05, 
    3.55889959069856e-05, 3.55889959069841e-05, 3.55889959069856e-05, 
    3.55889959069856e-05, 3.55889959069856e-05,
  3.57683773198826e-05, 3.57683773198826e-05, 3.57683773198826e-05, 
    3.57683773198765e-05, 3.57683773198826e-05, 3.57683773198826e-05, 
    3.57683773198765e-05, 3.57683773198826e-05, 3.57683773198826e-05, 
    3.57683773198765e-05, 3.57683773198826e-05, 3.57683773198826e-05, 
    3.57683773198765e-05, 3.57683773198826e-05, 3.57683773198826e-05, 
    3.57683773198765e-05, 3.57683773198826e-05, 3.57683773198826e-05, 
    3.57683773198796e-05, 3.57683773198796e-05, 3.57683773198796e-05, 
    3.57683773198826e-05, 3.57683773198796e-05, 3.57683773198796e-05, 
    3.57683773198826e-05, 3.57683773198796e-05, 3.57683773198796e-05, 
    3.57683773198826e-05, 3.57683773198796e-05, 3.57683773198796e-05, 
    3.57683773198826e-05, 3.57683773198796e-05, 3.57683773198796e-05, 
    3.57683773198826e-05, 3.57683773198796e-05, 3.57683773198796e-05, 
    3.57683773198826e-05, 3.57683773198796e-05, 3.57683773198796e-05, 
    3.57683773198826e-05, 3.57683773198796e-05, 3.57683773198796e-05, 
    3.57683773198826e-05, 3.57683773198796e-05, 3.57683773198796e-05, 
    3.57683773198826e-05, 3.57683773198796e-05, 3.57683773198796e-05, 
    3.57683773198826e-05, 3.57683773198796e-05, 3.57683773198811e-05, 
    3.57683773198811e-05, 3.57683773198796e-05, 3.57683773198811e-05, 
    3.57683773198811e-05, 3.57683773198811e-05,
  3.59507991504995e-05, 3.59507991504995e-05, 3.59507991504995e-05, 
    3.59507991504933e-05, 3.59507991504995e-05, 3.59507991504995e-05, 
    3.59507991504933e-05, 3.59507991504995e-05, 3.59507991504995e-05, 
    3.59507991504933e-05, 3.59507991504995e-05, 3.59507991504995e-05, 
    3.59507991504933e-05, 3.59507991504995e-05, 3.59507991504995e-05, 
    3.59507991504933e-05, 3.59507991504995e-05, 3.59507991504995e-05, 
    3.59507991504964e-05, 3.59507991504964e-05, 3.59507991504964e-05, 
    3.59507991504995e-05, 3.59507991504964e-05, 3.59507991504964e-05, 
    3.59507991504995e-05, 3.59507991504964e-05, 3.59507991504964e-05, 
    3.59507991504995e-05, 3.59507991504964e-05, 3.59507991504964e-05, 
    3.59507991504995e-05, 3.59507991504964e-05, 3.59507991504964e-05, 
    3.59507991504995e-05, 3.59507991504964e-05, 3.59507991504964e-05, 
    3.59507991504995e-05, 3.59507991504964e-05, 3.59507991504964e-05, 
    3.59507991504995e-05, 3.59507991504964e-05, 3.59507991504964e-05, 
    3.59507991504995e-05, 3.59507991504964e-05, 3.59507991504964e-05, 
    3.59507991504995e-05, 3.59507991504964e-05, 3.59507991504964e-05, 
    3.59507991504995e-05, 3.59507991504964e-05, 3.59507991504979e-05, 
    3.59507991504979e-05, 3.59507991504964e-05, 3.59507991504979e-05, 
    3.59507991504979e-05, 3.59507991504979e-05,
  3.61363206014253e-05, 3.61363206014253e-05, 3.61363206014253e-05, 
    3.61363206014191e-05, 3.61363206014253e-05, 3.61363206014253e-05, 
    3.61363206014191e-05, 3.61363206014253e-05, 3.61363206014253e-05, 
    3.61363206014191e-05, 3.61363206014253e-05, 3.61363206014253e-05, 
    3.61363206014191e-05, 3.61363206014253e-05, 3.61363206014253e-05, 
    3.61363206014191e-05, 3.61363206014253e-05, 3.61363206014253e-05, 
    3.61363206014222e-05, 3.61363206014222e-05, 3.61363206014222e-05, 
    3.61363206014253e-05, 3.61363206014222e-05, 3.61363206014222e-05, 
    3.61363206014253e-05, 3.61363206014222e-05, 3.61363206014222e-05, 
    3.61363206014253e-05, 3.61363206014222e-05, 3.61363206014222e-05, 
    3.61363206014253e-05, 3.61363206014222e-05, 3.61363206014222e-05, 
    3.61363206014253e-05, 3.61363206014222e-05, 3.61363206014222e-05, 
    3.61363206014253e-05, 3.61363206014222e-05, 3.61363206014222e-05, 
    3.61363206014253e-05, 3.61363206014222e-05, 3.61363206014222e-05, 
    3.61363206014253e-05, 3.61363206014222e-05, 3.61363206014222e-05, 
    3.61363206014253e-05, 3.61363206014222e-05, 3.61363206014222e-05, 
    3.61363206014253e-05, 3.61363206014222e-05, 3.61363206014237e-05, 
    3.61363206014237e-05, 3.61363206014222e-05, 3.61363206014237e-05, 
    3.61363206014237e-05, 3.61363206014237e-05,
  3.63250025652185e-05, 3.63250025652185e-05, 3.63250025652185e-05, 
    3.63250025652123e-05, 3.63250025652185e-05, 3.63250025652185e-05, 
    3.63250025652123e-05, 3.63250025652185e-05, 3.63250025652185e-05, 
    3.63250025652123e-05, 3.63250025652185e-05, 3.63250025652185e-05, 
    3.63250025652123e-05, 3.63250025652185e-05, 3.63250025652185e-05, 
    3.63250025652123e-05, 3.63250025652185e-05, 3.63250025652185e-05, 
    3.63250025652154e-05, 3.63250025652154e-05, 3.63250025652154e-05, 
    3.63250025652185e-05, 3.63250025652154e-05, 3.63250025652154e-05, 
    3.63250025652185e-05, 3.63250025652154e-05, 3.63250025652154e-05, 
    3.63250025652185e-05, 3.63250025652154e-05, 3.63250025652154e-05, 
    3.63250025652185e-05, 3.63250025652154e-05, 3.63250025652154e-05, 
    3.63250025652185e-05, 3.63250025652154e-05, 3.63250025652154e-05, 
    3.63250025652185e-05, 3.63250025652154e-05, 3.63250025652154e-05, 
    3.63250025652185e-05, 3.63250025652154e-05, 3.63250025652154e-05, 
    3.63250025652185e-05, 3.63250025652154e-05, 3.63250025652154e-05, 
    3.63250025652185e-05, 3.63250025652154e-05, 3.63250025652154e-05, 
    3.63250025652185e-05, 3.63250025652154e-05, 3.6325002565217e-05, 
    3.6325002565217e-05, 3.63250025652154e-05, 3.6325002565217e-05, 
    3.6325002565217e-05, 3.6325002565217e-05,
  3.65169076829657e-05, 3.65169076829657e-05, 3.65169076829657e-05, 
    3.65169076829595e-05, 3.65169076829657e-05, 3.65169076829657e-05, 
    3.65169076829595e-05, 3.65169076829657e-05, 3.65169076829657e-05, 
    3.65169076829595e-05, 3.65169076829657e-05, 3.65169076829657e-05, 
    3.65169076829595e-05, 3.65169076829657e-05, 3.65169076829657e-05, 
    3.65169076829595e-05, 3.65169076829657e-05, 3.65169076829657e-05, 
    3.65169076829626e-05, 3.65169076829626e-05, 3.65169076829626e-05, 
    3.65169076829657e-05, 3.65169076829626e-05, 3.65169076829626e-05, 
    3.65169076829657e-05, 3.65169076829626e-05, 3.65169076829626e-05, 
    3.65169076829657e-05, 3.65169076829626e-05, 3.65169076829626e-05, 
    3.65169076829657e-05, 3.65169076829626e-05, 3.65169076829626e-05, 
    3.65169076829657e-05, 3.65169076829626e-05, 3.65169076829626e-05, 
    3.65169076829657e-05, 3.65169076829626e-05, 3.65169076829626e-05, 
    3.65169076829657e-05, 3.65169076829626e-05, 3.65169076829626e-05, 
    3.65169076829657e-05, 3.65169076829626e-05, 3.65169076829626e-05, 
    3.65169076829657e-05, 3.65169076829626e-05, 3.65169076829626e-05, 
    3.65169076829657e-05, 3.65169076829626e-05, 3.65169076829642e-05, 
    3.65169076829642e-05, 3.65169076829626e-05, 3.65169076829642e-05, 
    3.65169076829642e-05, 3.65169076829642e-05,
  3.67121004053212e-05, 3.67121004053212e-05, 3.67121004053212e-05, 
    3.6712100405315e-05, 3.67121004053212e-05, 3.67121004053212e-05, 
    3.6712100405315e-05, 3.67121004053212e-05, 3.67121004053212e-05, 
    3.6712100405315e-05, 3.67121004053212e-05, 3.67121004053212e-05, 
    3.6712100405315e-05, 3.67121004053212e-05, 3.67121004053212e-05, 
    3.6712100405315e-05, 3.67121004053212e-05, 3.67121004053212e-05, 
    3.67121004053181e-05, 3.67121004053181e-05, 3.67121004053181e-05, 
    3.67121004053212e-05, 3.67121004053181e-05, 3.67121004053181e-05, 
    3.67121004053212e-05, 3.67121004053181e-05, 3.67121004053181e-05, 
    3.67121004053212e-05, 3.67121004053181e-05, 3.67121004053181e-05, 
    3.67121004053212e-05, 3.67121004053181e-05, 3.67121004053181e-05, 
    3.67121004053212e-05, 3.67121004053181e-05, 3.67121004053181e-05, 
    3.67121004053212e-05, 3.67121004053181e-05, 3.67121004053181e-05, 
    3.67121004053212e-05, 3.67121004053181e-05, 3.67121004053181e-05, 
    3.67121004053212e-05, 3.67121004053181e-05, 3.67121004053181e-05, 
    3.67121004053212e-05, 3.67121004053181e-05, 3.67121004053181e-05, 
    3.67121004053212e-05, 3.67121004053181e-05, 3.67121004053197e-05, 
    3.67121004053197e-05, 3.67121004053181e-05, 3.67121004053197e-05, 
    3.67121004053197e-05, 3.67121004053197e-05,
  3.69106470561529e-05, 3.69106470561529e-05, 3.69106470561529e-05, 
    3.69106470561466e-05, 3.69106470561529e-05, 3.69106470561529e-05, 
    3.69106470561466e-05, 3.69106470561529e-05, 3.69106470561529e-05, 
    3.69106470561466e-05, 3.69106470561529e-05, 3.69106470561529e-05, 
    3.69106470561466e-05, 3.69106470561529e-05, 3.69106470561529e-05, 
    3.69106470561466e-05, 3.69106470561529e-05, 3.69106470561529e-05, 
    3.69106470561498e-05, 3.69106470561498e-05, 3.69106470561498e-05, 
    3.69106470561529e-05, 3.69106470561498e-05, 3.69106470561498e-05, 
    3.69106470561529e-05, 3.69106470561498e-05, 3.69106470561498e-05, 
    3.69106470561529e-05, 3.69106470561498e-05, 3.69106470561498e-05, 
    3.69106470561529e-05, 3.69106470561498e-05, 3.69106470561498e-05, 
    3.69106470561529e-05, 3.69106470561498e-05, 3.69106470561498e-05, 
    3.69106470561529e-05, 3.69106470561498e-05, 3.69106470561498e-05, 
    3.69106470561529e-05, 3.69106470561498e-05, 3.69106470561498e-05, 
    3.69106470561529e-05, 3.69106470561498e-05, 3.69106470561498e-05, 
    3.69106470561529e-05, 3.69106470561498e-05, 3.69106470561498e-05, 
    3.69106470561529e-05, 3.69106470561498e-05, 3.69106470561514e-05, 
    3.69106470561514e-05, 3.69106470561498e-05, 3.69106470561514e-05, 
    3.69106470561514e-05, 3.69106470561514e-05,
  3.71126158989245e-05, 3.71126158989245e-05, 3.71126158989245e-05, 
    3.71126158989182e-05, 3.71126158989245e-05, 3.71126158989245e-05, 
    3.71126158989182e-05, 3.71126158989245e-05, 3.71126158989245e-05, 
    3.71126158989182e-05, 3.71126158989245e-05, 3.71126158989245e-05, 
    3.71126158989182e-05, 3.71126158989245e-05, 3.71126158989245e-05, 
    3.71126158989182e-05, 3.71126158989245e-05, 3.71126158989245e-05, 
    3.71126158989213e-05, 3.71126158989213e-05, 3.71126158989213e-05, 
    3.71126158989245e-05, 3.71126158989213e-05, 3.71126158989213e-05, 
    3.71126158989245e-05, 3.71126158989213e-05, 3.71126158989213e-05, 
    3.71126158989245e-05, 3.71126158989213e-05, 3.71126158989213e-05, 
    3.71126158989245e-05, 3.71126158989213e-05, 3.71126158989213e-05, 
    3.71126158989245e-05, 3.71126158989213e-05, 3.71126158989213e-05, 
    3.71126158989245e-05, 3.71126158989213e-05, 3.71126158989213e-05, 
    3.71126158989245e-05, 3.71126158989213e-05, 3.71126158989213e-05, 
    3.71126158989245e-05, 3.71126158989213e-05, 3.71126158989213e-05, 
    3.71126158989245e-05, 3.71126158989213e-05, 3.71126158989213e-05, 
    3.71126158989245e-05, 3.71126158989213e-05, 3.71126158989229e-05, 
    3.71126158989229e-05, 3.71126158989213e-05, 3.71126158989229e-05, 
    3.71126158989229e-05, 3.71126158989229e-05,
  3.73180772059509e-05, 3.73180772059509e-05, 3.73180772059509e-05, 
    3.73180772059446e-05, 3.73180772059509e-05, 3.73180772059509e-05, 
    3.73180772059446e-05, 3.73180772059509e-05, 3.73180772059509e-05, 
    3.73180772059446e-05, 3.73180772059509e-05, 3.73180772059509e-05, 
    3.73180772059446e-05, 3.73180772059509e-05, 3.73180772059509e-05, 
    3.73180772059446e-05, 3.73180772059509e-05, 3.73180772059509e-05, 
    3.73180772059478e-05, 3.73180772059478e-05, 3.73180772059478e-05, 
    3.73180772059509e-05, 3.73180772059478e-05, 3.73180772059478e-05, 
    3.73180772059509e-05, 3.73180772059478e-05, 3.73180772059478e-05, 
    3.73180772059509e-05, 3.73180772059478e-05, 3.73180772059478e-05, 
    3.73180772059509e-05, 3.73180772059478e-05, 3.73180772059478e-05, 
    3.73180772059509e-05, 3.73180772059478e-05, 3.73180772059478e-05, 
    3.73180772059509e-05, 3.73180772059478e-05, 3.73180772059478e-05, 
    3.73180772059509e-05, 3.73180772059478e-05, 3.73180772059478e-05, 
    3.73180772059509e-05, 3.73180772059478e-05, 3.73180772059478e-05, 
    3.73180772059509e-05, 3.73180772059478e-05, 3.73180772059478e-05, 
    3.73180772059509e-05, 3.73180772059478e-05, 3.73180772059494e-05, 
    3.73180772059494e-05, 3.73180772059478e-05, 3.73180772059494e-05, 
    3.73180772059494e-05, 3.73180772059494e-05,
  3.75271033306738e-05, 3.75271033306738e-05, 3.75271033306738e-05, 
    3.75271033306674e-05, 3.75271033306738e-05, 3.75271033306738e-05, 
    3.75271033306674e-05, 3.75271033306738e-05, 3.75271033306738e-05, 
    3.75271033306674e-05, 3.75271033306738e-05, 3.75271033306738e-05, 
    3.75271033306674e-05, 3.75271033306738e-05, 3.75271033306738e-05, 
    3.75271033306674e-05, 3.75271033306738e-05, 3.75271033306738e-05, 
    3.75271033306706e-05, 3.75271033306706e-05, 3.75271033306706e-05, 
    3.75271033306738e-05, 3.75271033306706e-05, 3.75271033306706e-05, 
    3.75271033306738e-05, 3.75271033306706e-05, 3.75271033306706e-05, 
    3.75271033306738e-05, 3.75271033306706e-05, 3.75271033306706e-05, 
    3.75271033306738e-05, 3.75271033306706e-05, 3.75271033306706e-05, 
    3.75271033306738e-05, 3.75271033306706e-05, 3.75271033306706e-05, 
    3.75271033306738e-05, 3.75271033306706e-05, 3.75271033306706e-05, 
    3.75271033306738e-05, 3.75271033306706e-05, 3.75271033306706e-05, 
    3.75271033306738e-05, 3.75271033306706e-05, 3.75271033306706e-05, 
    3.75271033306738e-05, 3.75271033306706e-05, 3.75271033306706e-05, 
    3.75271033306738e-05, 3.75271033306706e-05, 3.75271033306722e-05, 
    3.75271033306722e-05, 3.75271033306706e-05, 3.75271033306722e-05, 
    3.75271033306722e-05, 3.75271033306722e-05,
  3.77397687831096e-05, 3.77397687831096e-05, 3.77397687831096e-05, 
    3.77397687831032e-05, 3.77397687831096e-05, 3.77397687831096e-05, 
    3.77397687831032e-05, 3.77397687831096e-05, 3.77397687831096e-05, 
    3.77397687831032e-05, 3.77397687831096e-05, 3.77397687831096e-05, 
    3.77397687831032e-05, 3.77397687831096e-05, 3.77397687831096e-05, 
    3.77397687831032e-05, 3.77397687831096e-05, 3.77397687831096e-05, 
    3.77397687831064e-05, 3.77397687831064e-05, 3.77397687831064e-05, 
    3.77397687831096e-05, 3.77397687831064e-05, 3.77397687831064e-05, 
    3.77397687831096e-05, 3.77397687831064e-05, 3.77397687831064e-05, 
    3.77397687831096e-05, 3.77397687831064e-05, 3.77397687831064e-05, 
    3.77397687831096e-05, 3.77397687831064e-05, 3.77397687831064e-05, 
    3.77397687831096e-05, 3.77397687831064e-05, 3.77397687831064e-05, 
    3.77397687831096e-05, 3.77397687831064e-05, 3.77397687831064e-05, 
    3.77397687831096e-05, 3.77397687831064e-05, 3.77397687831064e-05, 
    3.77397687831096e-05, 3.77397687831064e-05, 3.77397687831064e-05, 
    3.77397687831096e-05, 3.77397687831064e-05, 3.77397687831064e-05, 
    3.77397687831096e-05, 3.77397687831064e-05, 3.7739768783108e-05, 
    3.7739768783108e-05, 3.77397687831064e-05, 3.7739768783108e-05, 
    3.7739768783108e-05, 3.7739768783108e-05,
  3.79561503086355e-05, 3.79561503086355e-05, 3.79561503086355e-05, 
    3.7956150308629e-05, 3.79561503086355e-05, 3.79561503086355e-05, 
    3.7956150308629e-05, 3.79561503086355e-05, 3.79561503086355e-05, 
    3.7956150308629e-05, 3.79561503086355e-05, 3.79561503086355e-05, 
    3.7956150308629e-05, 3.79561503086355e-05, 3.79561503086355e-05, 
    3.7956150308629e-05, 3.79561503086355e-05, 3.79561503086355e-05, 
    3.79561503086323e-05, 3.79561503086323e-05, 3.79561503086323e-05, 
    3.79561503086355e-05, 3.79561503086323e-05, 3.79561503086323e-05, 
    3.79561503086355e-05, 3.79561503086323e-05, 3.79561503086323e-05, 
    3.79561503086355e-05, 3.79561503086323e-05, 3.79561503086323e-05, 
    3.79561503086355e-05, 3.79561503086323e-05, 3.79561503086323e-05, 
    3.79561503086355e-05, 3.79561503086323e-05, 3.79561503086323e-05, 
    3.79561503086355e-05, 3.79561503086323e-05, 3.79561503086323e-05, 
    3.79561503086355e-05, 3.79561503086323e-05, 3.79561503086323e-05, 
    3.79561503086355e-05, 3.79561503086323e-05, 3.79561503086323e-05, 
    3.79561503086355e-05, 3.79561503086323e-05, 3.79561503086323e-05, 
    3.79561503086355e-05, 3.79561503086323e-05, 3.79561503086339e-05, 
    3.79561503086339e-05, 3.79561503086323e-05, 3.79561503086339e-05, 
    3.79561503086339e-05, 3.79561503086339e-05,
  3.81763269702841e-05, 3.81763269702841e-05, 3.81763269702841e-05, 
    3.81763269702775e-05, 3.81763269702841e-05, 3.81763269702841e-05, 
    3.81763269702775e-05, 3.81763269702841e-05, 3.81763269702841e-05, 
    3.81763269702775e-05, 3.81763269702841e-05, 3.81763269702841e-05, 
    3.81763269702775e-05, 3.81763269702841e-05, 3.81763269702841e-05, 
    3.81763269702775e-05, 3.81763269702841e-05, 3.81763269702841e-05, 
    3.81763269702808e-05, 3.81763269702808e-05, 3.81763269702808e-05, 
    3.81763269702841e-05, 3.81763269702808e-05, 3.81763269702808e-05, 
    3.81763269702841e-05, 3.81763269702808e-05, 3.81763269702808e-05, 
    3.81763269702841e-05, 3.81763269702808e-05, 3.81763269702808e-05, 
    3.81763269702841e-05, 3.81763269702808e-05, 3.81763269702808e-05, 
    3.81763269702841e-05, 3.81763269702808e-05, 3.81763269702808e-05, 
    3.81763269702841e-05, 3.81763269702808e-05, 3.81763269702808e-05, 
    3.81763269702841e-05, 3.81763269702808e-05, 3.81763269702808e-05, 
    3.81763269702841e-05, 3.81763269702808e-05, 3.81763269702808e-05, 
    3.81763269702841e-05, 3.81763269702808e-05, 3.81763269702808e-05, 
    3.81763269702841e-05, 3.81763269702808e-05, 3.81763269702824e-05, 
    3.81763269702824e-05, 3.81763269702808e-05, 3.81763269702824e-05, 
    3.81763269702824e-05, 3.81763269702824e-05,
  3.8400380234731e-05, 3.8400380234731e-05, 3.8400380234731e-05, 
    3.84003802347244e-05, 3.8400380234731e-05, 3.8400380234731e-05, 
    3.84003802347244e-05, 3.8400380234731e-05, 3.8400380234731e-05, 
    3.84003802347244e-05, 3.8400380234731e-05, 3.8400380234731e-05, 
    3.84003802347244e-05, 3.8400380234731e-05, 3.8400380234731e-05, 
    3.84003802347244e-05, 3.8400380234731e-05, 3.8400380234731e-05, 
    3.84003802347277e-05, 3.84003802347277e-05, 3.84003802347277e-05, 
    3.8400380234731e-05, 3.84003802347277e-05, 3.84003802347277e-05, 
    3.8400380234731e-05, 3.84003802347277e-05, 3.84003802347277e-05, 
    3.8400380234731e-05, 3.84003802347277e-05, 3.84003802347277e-05, 
    3.8400380234731e-05, 3.84003802347277e-05, 3.84003802347277e-05, 
    3.8400380234731e-05, 3.84003802347277e-05, 3.84003802347277e-05, 
    3.8400380234731e-05, 3.84003802347277e-05, 3.84003802347277e-05, 
    3.8400380234731e-05, 3.84003802347277e-05, 3.84003802347277e-05, 
    3.8400380234731e-05, 3.84003802347277e-05, 3.84003802347277e-05, 
    3.8400380234731e-05, 3.84003802347277e-05, 3.84003802347277e-05, 
    3.8400380234731e-05, 3.84003802347277e-05, 3.84003802347294e-05, 
    3.84003802347294e-05, 3.84003802347277e-05, 3.84003802347294e-05, 
    3.84003802347294e-05, 3.84003802347294e-05,
  3.86283940621702e-05, 3.86283940621702e-05, 3.86283940621702e-05, 
    3.86283940621636e-05, 3.86283940621702e-05, 3.86283940621702e-05, 
    3.86283940621636e-05, 3.86283940621702e-05, 3.86283940621702e-05, 
    3.86283940621636e-05, 3.86283940621702e-05, 3.86283940621702e-05, 
    3.86283940621636e-05, 3.86283940621702e-05, 3.86283940621702e-05, 
    3.86283940621636e-05, 3.86283940621702e-05, 3.86283940621702e-05, 
    3.86283940621669e-05, 3.86283940621669e-05, 3.86283940621669e-05, 
    3.86283940621702e-05, 3.86283940621669e-05, 3.86283940621669e-05, 
    3.86283940621702e-05, 3.86283940621669e-05, 3.86283940621669e-05, 
    3.86283940621702e-05, 3.86283940621669e-05, 3.86283940621669e-05, 
    3.86283940621702e-05, 3.86283940621669e-05, 3.86283940621669e-05, 
    3.86283940621702e-05, 3.86283940621669e-05, 3.86283940621669e-05, 
    3.86283940621702e-05, 3.86283940621669e-05, 3.86283940621669e-05, 
    3.86283940621702e-05, 3.86283940621669e-05, 3.86283940621669e-05, 
    3.86283940621702e-05, 3.86283940621669e-05, 3.86283940621669e-05, 
    3.86283940621702e-05, 3.86283940621669e-05, 3.86283940621669e-05, 
    3.86283940621702e-05, 3.86283940621669e-05, 3.86283940621685e-05, 
    3.86283940621685e-05, 3.86283940621669e-05, 3.86283940621685e-05, 
    3.86283940621685e-05, 3.86283940621685e-05,
  3.88604550002813e-05, 3.88604550002813e-05, 3.88604550002813e-05, 
    3.88604550002747e-05, 3.88604550002813e-05, 3.88604550002813e-05, 
    3.88604550002747e-05, 3.88604550002813e-05, 3.88604550002813e-05, 
    3.88604550002747e-05, 3.88604550002813e-05, 3.88604550002813e-05, 
    3.88604550002747e-05, 3.88604550002813e-05, 3.88604550002813e-05, 
    3.88604550002747e-05, 3.88604550002813e-05, 3.88604550002813e-05, 
    3.8860455000278e-05, 3.8860455000278e-05, 3.8860455000278e-05, 
    3.88604550002813e-05, 3.8860455000278e-05, 3.8860455000278e-05, 
    3.88604550002813e-05, 3.8860455000278e-05, 3.8860455000278e-05, 
    3.88604550002813e-05, 3.8860455000278e-05, 3.8860455000278e-05, 
    3.88604550002813e-05, 3.8860455000278e-05, 3.8860455000278e-05, 
    3.88604550002813e-05, 3.8860455000278e-05, 3.8860455000278e-05, 
    3.88604550002813e-05, 3.8860455000278e-05, 3.8860455000278e-05, 
    3.88604550002813e-05, 3.8860455000278e-05, 3.8860455000278e-05, 
    3.88604550002813e-05, 3.8860455000278e-05, 3.8860455000278e-05, 
    3.88604550002813e-05, 3.8860455000278e-05, 3.8860455000278e-05, 
    3.88604550002813e-05, 3.8860455000278e-05, 3.88604550002797e-05, 
    3.88604550002797e-05, 3.8860455000278e-05, 3.88604550002797e-05, 
    3.88604550002797e-05, 3.88604550002797e-05,
  3.90966522825095e-05, 3.90966522825095e-05, 3.90966522825095e-05, 
    3.90966522825028e-05, 3.90966522825095e-05, 3.90966522825095e-05, 
    3.90966522825028e-05, 3.90966522825095e-05, 3.90966522825095e-05, 
    3.90966522825028e-05, 3.90966522825095e-05, 3.90966522825095e-05, 
    3.90966522825028e-05, 3.90966522825095e-05, 3.90966522825095e-05, 
    3.90966522825028e-05, 3.90966522825095e-05, 3.90966522825095e-05, 
    3.90966522825061e-05, 3.90966522825061e-05, 3.90966522825061e-05, 
    3.90966522825095e-05, 3.90966522825061e-05, 3.90966522825061e-05, 
    3.90966522825095e-05, 3.90966522825061e-05, 3.90966522825061e-05, 
    3.90966522825095e-05, 3.90966522825061e-05, 3.90966522825061e-05, 
    3.90966522825095e-05, 3.90966522825061e-05, 3.90966522825061e-05, 
    3.90966522825095e-05, 3.90966522825061e-05, 3.90966522825061e-05, 
    3.90966522825095e-05, 3.90966522825061e-05, 3.90966522825061e-05, 
    3.90966522825095e-05, 3.90966522825061e-05, 3.90966522825061e-05, 
    3.90966522825095e-05, 3.90966522825061e-05, 3.90966522825061e-05, 
    3.90966522825095e-05, 3.90966522825061e-05, 3.90966522825061e-05, 
    3.90966522825095e-05, 3.90966522825061e-05, 3.90966522825078e-05, 
    3.90966522825078e-05, 3.90966522825061e-05, 3.90966522825078e-05, 
    3.90966522825078e-05, 3.90966522825078e-05,
  3.93370779308883e-05, 3.93370779308883e-05, 3.93370779308883e-05, 
    3.93370779308816e-05, 3.93370779308883e-05, 3.93370779308883e-05, 
    3.93370779308816e-05, 3.93370779308883e-05, 3.93370779308883e-05, 
    3.93370779308816e-05, 3.93370779308883e-05, 3.93370779308883e-05, 
    3.93370779308816e-05, 3.93370779308883e-05, 3.93370779308883e-05, 
    3.93370779308816e-05, 3.93370779308883e-05, 3.93370779308883e-05, 
    3.93370779308849e-05, 3.93370779308849e-05, 3.93370779308849e-05, 
    3.93370779308883e-05, 3.93370779308849e-05, 3.93370779308849e-05, 
    3.93370779308883e-05, 3.93370779308849e-05, 3.93370779308849e-05, 
    3.93370779308883e-05, 3.93370779308849e-05, 3.93370779308849e-05, 
    3.93370779308883e-05, 3.93370779308849e-05, 3.93370779308849e-05, 
    3.93370779308883e-05, 3.93370779308849e-05, 3.93370779308849e-05, 
    3.93370779308883e-05, 3.93370779308849e-05, 3.93370779308849e-05, 
    3.93370779308883e-05, 3.93370779308849e-05, 3.93370779308849e-05, 
    3.93370779308883e-05, 3.93370779308849e-05, 3.93370779308849e-05, 
    3.93370779308883e-05, 3.93370779308849e-05, 3.93370779308849e-05, 
    3.93370779308883e-05, 3.93370779308849e-05, 3.93370779308866e-05, 
    3.93370779308866e-05, 3.93370779308849e-05, 3.93370779308866e-05, 
    3.93370779308866e-05, 3.93370779308866e-05,
  3.9581826863653e-05, 3.9581826863653e-05, 3.9581826863653e-05, 
    3.95818268636462e-05, 3.9581826863653e-05, 3.9581826863653e-05, 
    3.95818268636462e-05, 3.9581826863653e-05, 3.9581826863653e-05, 
    3.95818268636462e-05, 3.9581826863653e-05, 3.9581826863653e-05, 
    3.95818268636462e-05, 3.9581826863653e-05, 3.9581826863653e-05, 
    3.95818268636462e-05, 3.9581826863653e-05, 3.9581826863653e-05, 
    3.95818268636496e-05, 3.95818268636496e-05, 3.95818268636496e-05, 
    3.9581826863653e-05, 3.95818268636496e-05, 3.95818268636496e-05, 
    3.9581826863653e-05, 3.95818268636496e-05, 3.95818268636496e-05, 
    3.9581826863653e-05, 3.95818268636496e-05, 3.95818268636496e-05, 
    3.9581826863653e-05, 3.95818268636496e-05, 3.95818268636496e-05, 
    3.9581826863653e-05, 3.95818268636496e-05, 3.95818268636496e-05, 
    3.9581826863653e-05, 3.95818268636496e-05, 3.95818268636496e-05, 
    3.9581826863653e-05, 3.95818268636496e-05, 3.95818268636496e-05, 
    3.9581826863653e-05, 3.95818268636496e-05, 3.95818268636496e-05, 
    3.9581826863653e-05, 3.95818268636496e-05, 3.95818268636496e-05, 
    3.9581826863653e-05, 3.95818268636496e-05, 3.95818268636513e-05, 
    3.95818268636513e-05, 3.95818268636496e-05, 3.95818268636513e-05, 
    3.95818268636513e-05, 3.95818268636513e-05,
  3.98309970079057e-05, 3.98309970079057e-05, 3.98309970079057e-05, 
    3.98309970078989e-05, 3.98309970079057e-05, 3.98309970079057e-05, 
    3.98309970078989e-05, 3.98309970079057e-05, 3.98309970079057e-05, 
    3.98309970078989e-05, 3.98309970079057e-05, 3.98309970079057e-05, 
    3.98309970078989e-05, 3.98309970079057e-05, 3.98309970079057e-05, 
    3.98309970078989e-05, 3.98309970079057e-05, 3.98309970079057e-05, 
    3.98309970079023e-05, 3.98309970079023e-05, 3.98309970079023e-05, 
    3.98309970079057e-05, 3.98309970079023e-05, 3.98309970079023e-05, 
    3.98309970079057e-05, 3.98309970079023e-05, 3.98309970079023e-05, 
    3.98309970079057e-05, 3.98309970079023e-05, 3.98309970079023e-05, 
    3.98309970079057e-05, 3.98309970079023e-05, 3.98309970079023e-05, 
    3.98309970079057e-05, 3.98309970079023e-05, 3.98309970079023e-05, 
    3.98309970079057e-05, 3.98309970079023e-05, 3.98309970079023e-05, 
    3.98309970079057e-05, 3.98309970079023e-05, 3.98309970079023e-05, 
    3.98309970079057e-05, 3.98309970079023e-05, 3.98309970079023e-05, 
    3.98309970079057e-05, 3.98309970079023e-05, 3.98309970079023e-05, 
    3.98309970079057e-05, 3.98309970079023e-05, 3.9830997007904e-05, 
    3.9830997007904e-05, 3.98309970079023e-05, 3.9830997007904e-05, 
    3.9830997007904e-05, 3.9830997007904e-05,
  4.00846894176107e-05, 4.00846894176107e-05, 4.00846894176107e-05, 
    4.00846894176039e-05, 4.00846894176107e-05, 4.00846894176107e-05, 
    4.00846894176039e-05, 4.00846894176107e-05, 4.00846894176107e-05, 
    4.00846894176039e-05, 4.00846894176107e-05, 4.00846894176107e-05, 
    4.00846894176039e-05, 4.00846894176107e-05, 4.00846894176107e-05, 
    4.00846894176039e-05, 4.00846894176107e-05, 4.00846894176107e-05, 
    4.00846894176073e-05, 4.00846894176073e-05, 4.00846894176073e-05, 
    4.00846894176107e-05, 4.00846894176073e-05, 4.00846894176073e-05, 
    4.00846894176107e-05, 4.00846894176073e-05, 4.00846894176073e-05, 
    4.00846894176107e-05, 4.00846894176073e-05, 4.00846894176073e-05, 
    4.00846894176107e-05, 4.00846894176073e-05, 4.00846894176073e-05, 
    4.00846894176107e-05, 4.00846894176073e-05, 4.00846894176073e-05, 
    4.00846894176107e-05, 4.00846894176073e-05, 4.00846894176073e-05, 
    4.00846894176107e-05, 4.00846894176073e-05, 4.00846894176073e-05, 
    4.00846894176107e-05, 4.00846894176073e-05, 4.00846894176073e-05, 
    4.00846894176107e-05, 4.00846894176073e-05, 4.00846894176073e-05, 
    4.00846894176107e-05, 4.00846894176073e-05, 4.0084689417609e-05, 
    4.0084689417609e-05, 4.00846894176073e-05, 4.0084689417609e-05, 
    4.0084689417609e-05, 4.0084689417609e-05,
  4.03430083972161e-05, 4.03430083972161e-05, 4.03430083972161e-05, 
    4.03430083972093e-05, 4.03430083972161e-05, 4.03430083972161e-05, 
    4.03430083972093e-05, 4.03430083972161e-05, 4.03430083972161e-05, 
    4.03430083972093e-05, 4.03430083972161e-05, 4.03430083972161e-05, 
    4.03430083972093e-05, 4.03430083972161e-05, 4.03430083972161e-05, 
    4.03430083972093e-05, 4.03430083972161e-05, 4.03430083972161e-05, 
    4.03430083972127e-05, 4.03430083972127e-05, 4.03430083972127e-05, 
    4.03430083972161e-05, 4.03430083972127e-05, 4.03430083972127e-05, 
    4.03430083972161e-05, 4.03430083972127e-05, 4.03430083972127e-05, 
    4.03430083972161e-05, 4.03430083972127e-05, 4.03430083972127e-05, 
    4.03430083972161e-05, 4.03430083972127e-05, 4.03430083972127e-05, 
    4.03430083972161e-05, 4.03430083972127e-05, 4.03430083972127e-05, 
    4.03430083972161e-05, 4.03430083972127e-05, 4.03430083972127e-05, 
    4.03430083972161e-05, 4.03430083972127e-05, 4.03430083972127e-05, 
    4.03430083972161e-05, 4.03430083972127e-05, 4.03430083972127e-05, 
    4.03430083972161e-05, 4.03430083972127e-05, 4.03430083972127e-05, 
    4.03430083972161e-05, 4.03430083972127e-05, 4.03430083972144e-05, 
    4.03430083972144e-05, 4.03430083972127e-05, 4.03430083972144e-05, 
    4.03430083972144e-05, 4.03430083972144e-05 ;

 pn =
  2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05,
  2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05,
  2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05,
  2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05,
  2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05,
  2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05,
  2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05,
  2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05,
  2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05,
  2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05,
  2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05,
  2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05,
  2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05,
  2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05,
  2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05,
  2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05,
  2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05,
  2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05,
  2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05,
  2.69947206465744e-05, 2.69947206465744e-05, 2.69947206465744e-05, 
    2.69947206465744e-05, 2.69947206465744e-05, 2.69947206465744e-05, 
    2.69947206465744e-05, 2.69947206465744e-05, 2.69947206465744e-05, 
    2.69947206465744e-05, 2.69947206465744e-05, 2.69947206465744e-05, 
    2.69947206465744e-05, 2.69947206465744e-05, 2.69947206465744e-05, 
    2.69947206465744e-05, 2.69947206465744e-05, 2.69947206465744e-05, 
    2.69947206465744e-05, 2.69947206465744e-05, 2.69947206465744e-05, 
    2.69947206465744e-05, 2.69947206465744e-05, 2.69947206465744e-05, 
    2.69947206465744e-05, 2.69947206465744e-05, 2.69947206465744e-05, 
    2.69947206465744e-05, 2.69947206465744e-05, 2.69947206465744e-05, 
    2.69947206465744e-05, 2.69947206465744e-05, 2.69947206465744e-05, 
    2.69947206465744e-05, 2.69947206465744e-05, 2.69947206465744e-05, 
    2.69947206465744e-05, 2.69947206465744e-05, 2.69947206465744e-05, 
    2.69947206465744e-05, 2.69947206465744e-05, 2.69947206465744e-05, 
    2.69947206465744e-05, 2.69947206465744e-05, 2.69947206465744e-05, 
    2.69947206465744e-05, 2.69947206465744e-05, 2.69947206465744e-05, 
    2.69947206465744e-05, 2.69947206465744e-05, 2.69947206465744e-05, 
    2.69947206465744e-05, 2.69947206465744e-05, 2.69947206465744e-05, 
    2.69947206465744e-05, 2.69947206465744e-05,
  2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05,
  2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05,
  2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05,
  2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05,
  2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05,
  2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05,
  2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05,
  2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05, 2.69947206465726e-05, 
    2.69947206465726e-05, 2.69947206465726e-05,
  2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05, 2.69947206465739e-05, 
    2.69947206465739e-05, 2.69947206465739e-05,
  2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05,
  2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05,
  2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05,
  2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05,
  2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05,
  2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05,
  2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05,
  2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05,
  2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05,
  2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05,
  2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05,
  2.69947206465747e-05, 2.69947206465747e-05, 2.69947206465747e-05, 
    2.69947206465747e-05, 2.69947206465747e-05, 2.69947206465747e-05, 
    2.69947206465747e-05, 2.69947206465747e-05, 2.69947206465747e-05, 
    2.69947206465747e-05, 2.69947206465747e-05, 2.69947206465747e-05, 
    2.69947206465747e-05, 2.69947206465747e-05, 2.69947206465747e-05, 
    2.69947206465747e-05, 2.69947206465747e-05, 2.69947206465747e-05, 
    2.69947206465747e-05, 2.69947206465747e-05, 2.69947206465747e-05, 
    2.69947206465747e-05, 2.69947206465747e-05, 2.69947206465747e-05, 
    2.69947206465747e-05, 2.69947206465747e-05, 2.69947206465747e-05, 
    2.69947206465747e-05, 2.69947206465747e-05, 2.69947206465747e-05, 
    2.69947206465747e-05, 2.69947206465747e-05, 2.69947206465747e-05, 
    2.69947206465747e-05, 2.69947206465747e-05, 2.69947206465747e-05, 
    2.69947206465747e-05, 2.69947206465747e-05, 2.69947206465747e-05, 
    2.69947206465747e-05, 2.69947206465747e-05, 2.69947206465747e-05, 
    2.69947206465747e-05, 2.69947206465747e-05, 2.69947206465747e-05, 
    2.69947206465747e-05, 2.69947206465747e-05, 2.69947206465747e-05, 
    2.69947206465747e-05, 2.69947206465747e-05, 2.69947206465747e-05, 
    2.69947206465747e-05, 2.69947206465747e-05, 2.69947206465747e-05, 
    2.69947206465747e-05, 2.69947206465747e-05,
  2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05, 2.69947206465729e-05, 
    2.69947206465729e-05, 2.69947206465729e-05,
  2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05,
  2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05,
  2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05,
  2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05,
  2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05,
  2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05,
  2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05, 2.69947206465731e-05, 
    2.69947206465731e-05, 2.69947206465731e-05,
  2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05,
  2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05, 2.69947206465736e-05, 
    2.69947206465736e-05, 2.69947206465736e-05,
  2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05, 2.69947206465742e-05, 
    2.69947206465742e-05, 2.69947206465742e-05,
  2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05,
  2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05,
  2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05, 2.69947206465734e-05, 
    2.69947206465734e-05, 2.69947206465734e-05 ;

 dndx =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0 ;

 dmde =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0 ;

 x_rho =
  0, 32081.2765499785, 64162.5530999569, 96243.8296499381, 128325.106199919, 
    160406.382749898, 192487.659299879, 224568.93584986, 256650.212399839, 
    288731.48894982, 320812.765499801, 352894.042049779, 384975.318599761, 
    417056.595149742, 449137.87169972, 481219.148249701, 513300.424799683, 
    545381.701349661, 577462.977899641, 609544.254449622, 641625.530999603, 
    673706.807549583, 705788.084099563, 737869.360649544, 769950.637199524, 
    802031.913749504, 834113.190299485, 866194.466849465, 898275.743399445, 
    930357.019949426, 962438.296499406, 994519.573049385, 1026600.84959937, 
    1058682.12614935, 1090763.40269933, 1122844.67924931, 1154925.95579929, 
    1187007.23234927, 1219088.50889925, 1251169.78544923, 1283251.06199921, 
    1315332.33854919, 1347413.61509917, 1379494.89164915, 1411576.16819913, 
    1443657.44474911, 1475738.72129909, 1507819.99784907, 1539901.27439905, 
    1571982.55094903, 1604063.82749901, 1636145.10404899, 1668226.38059897, 
    1700307.65714895, 1732388.93369893, 1764470.21024891,
  0, 31972.9766083239, 63945.9532166477, 95918.9298249743, 127891.906433301, 
    159864.883041625, 191837.859649951, 223810.836258278, 255783.812866602, 
    287756.789474928, 319729.766083255, 351702.742691579, 383675.719299905, 
    415648.695908232, 447621.672516556, 479594.649124882, 511567.625733209, 
    543540.602341533, 575513.578949858, 607486.555558185, 639459.532166511, 
    671432.508774836, 703405.485383162, 735378.461991488, 767351.438599813, 
    799324.415208139, 831297.391816465, 863270.368424791, 895243.345033116, 
    927216.321641442, 959189.298249768, 991162.274858093, 1023135.25146642, 
    1055108.22807474, 1087081.20468307, 1119054.1812914, 1151027.15789972, 
    1183000.13450805, 1214973.11111637, 1246946.0877247, 1278919.06433302, 
    1310892.04094135, 1342865.01754968, 1374837.994158, 1406810.97076633, 
    1438783.94737465, 1470756.92398298, 1502729.90059131, 1534702.87719963, 
    1566675.85380796, 1598648.83041628, 1630621.80702461, 1662594.78363293, 
    1694567.76024126, 1726540.73684958, 1758513.71345791,
  0, 31863.594500268, 63727.189000536, 95590.7835008067, 127454.378001077, 
    159317.972501345, 191181.567001616, 223045.161501887, 254908.756002155, 
    286772.350502426, 318635.945002696, 350499.539502964, 382363.134003235, 
    414226.728503506, 446090.323003774, 477953.917504045, 509817.512004315, 
    541681.106504583, 573544.701004853, 605408.295505123, 637271.890005394, 
    669135.484505663, 700999.079005933, 732862.673506203, 764726.268006473, 
    796589.862506742, 828453.457007013, 860317.051507282, 892180.646007552, 
    924044.240507822, 955907.835008092, 987771.429508361, 1019635.02400863, 
    1051498.6185089, 1083362.21300917, 1115225.80750944, 1147089.40200971, 
    1178952.99650998, 1210816.59101025, 1242680.18551052, 1274543.78001079, 
    1306407.37451106, 1338270.96901133, 1370134.5635116, 1401998.15801187, 
    1433861.75251214, 1465725.34701241, 1497588.94151268, 1529452.53601295, 
    1561316.13051322, 1593179.72501349, 1625043.31951376, 1656906.91401403, 
    1688770.5085143, 1720634.10301457, 1752497.69751483,
  0, 31753.1339280506, 63506.2678561011, 95259.4017841544, 127012.535712208, 
    158765.669640258, 190518.803568312, 222271.937496365, 254025.071424415, 
    285778.205352469, 317531.339280522, 349284.473208573, 381037.607136626, 
    412790.741064679, 444543.87499273, 476297.008920783, 508050.142848836, 
    539803.276776887, 571556.410704939, 603309.544632992, 635062.678561045, 
    666815.812489097, 698568.946417149, 730322.080345202, 762075.214273254, 
    793828.348201306, 825581.48212936, 857334.616057411, 889087.749985463, 
    920840.883913517, 952594.017841569, 984347.15176962, 1016100.28569767, 
    1047853.41962573, 1079606.55355378, 1111359.68748183, 1143112.82140988, 
    1174865.95533793, 1206619.08926599, 1238372.22319404, 1270125.35712209, 
    1301878.49105015, 1333631.6249782, 1365384.75890625, 1397137.8928343, 
    1428891.02676235, 1460644.16069041, 1492397.29461846, 1524150.42854651, 
    1555903.56247456, 1587656.69640262, 1619409.83033067, 1651162.96425872, 
    1682916.09818677, 1714669.23211483, 1746422.36604288,
  0, 31641.5986304132, 63283.1972608263, 94924.7958912422, 126566.394521658, 
    158207.993152071, 189849.591782487, 221491.190412903, 253132.789043316, 
    284774.387673732, 316415.986304148, 348057.584934561, 379699.183564977, 
    411340.782195393, 442982.380825806, 474623.979456222, 506265.578086638, 
    537907.176717051, 569548.775347465, 601190.373977881, 632831.972608297, 
    664473.571238711, 696115.169869126, 727756.768499542, 759398.367129956, 
    791039.965760371, 822681.564390786, 854323.163021201, 885964.761651615, 
    917606.360282031, 949247.958912446, 980889.55754286, 1012531.15617328, 
    1044172.75480369, 1075814.3534341, 1107455.95206452, 1139097.55069494, 
    1170739.14932535, 1202380.74795577, 1234022.34658618, 1265663.94521659, 
    1297305.54384701, 1328947.14247743, 1360588.74110784, 1392230.33973826, 
    1423871.93836867, 1455513.53699908, 1487155.1356295, 1518796.73425991, 
    1550438.33289033, 1582079.93152074, 1613721.53015116, 1645363.12878157, 
    1677004.72741199, 1708646.3260424, 1740287.92467282,
  0, 31528.9923824728, 63057.9847649456, 94586.977147421, 126115.969529897, 
    157644.961912369, 189173.954294845, 220702.94667732, 252231.939059793, 
    283760.931442268, 315289.923824744, 346818.916207217, 378347.908589692, 
    409876.900972168, 441405.89335464, 472934.885737116, 504463.878119591, 
    535992.870502064, 567521.862884538, 599050.855267014, 630579.847649489, 
    662108.840031963, 693637.832414438, 725166.824796913, 756695.817179387, 
    788224.809561861, 819753.801944337, 851282.794326811, 882811.786709285, 
    914340.779091761, 945869.771474235, 977398.763856709, 1008927.75623918, 
    1040456.74862166, 1071985.74100413, 1103514.73338661, 1135043.72576908, 
    1166572.71815156, 1198101.71053403, 1229630.70291651, 1261159.69529898, 
    1292688.68768146, 1324217.68006393, 1355746.6724464, 1387275.66482888, 
    1418804.65721135, 1450333.64959383, 1481862.6419763, 1513391.63435878, 
    1544920.62674125, 1576449.61912373, 1607978.6115062, 1639507.60388868, 
    1671036.59627115, 1702565.58865362, 1734094.5810361,
  0, 31415.3189955941, 62830.6379911882, 94245.9569867849, 125661.275982382, 
    157076.594977976, 188491.913973573, 219907.232969169, 251322.551964763, 
    282737.87096036, 314153.189955957, 345568.508951551, 376983.827947148, 
    408399.146942745, 439814.465938339, 471229.784933936, 502645.103929532, 
    534060.422925126, 565475.741920722, 596891.060916319, 628306.379911915, 
    659721.698907511, 691137.017903106, 722552.336898703, 753967.655894298, 
    785382.974889894, 816798.293885491, 848213.612881086, 879628.931876681, 
    911044.250872278, 942459.569867874, 973874.888863469, 1005290.20785907, 
    1036705.52685466, 1068120.84585026, 1099536.16484585, 1130951.48384145, 
    1162366.80283704, 1193782.12183264, 1225197.44082824, 1256612.75982383, 
    1288028.07881943, 1319443.39781502, 1350858.71681062, 1382274.03580622, 
    1413689.35480181, 1445104.67379741, 1476519.992793, 1507935.3117886, 
    1539350.6307842, 1570765.94977979, 1602181.26877539, 1633596.58777098, 
    1665011.90676658, 1696427.22576217, 1727842.54475777,
  0, 31300.5823172603, 62601.1646345206, 93901.7469517836, 125202.329269047, 
    156502.911586307, 187803.49390357, 219104.076220833, 250404.658538093, 
    281705.240855356, 313005.823172619, 344306.405489879, 375606.987807142, 
    406907.570124405, 438208.152441666, 469508.734758929, 500809.317076192, 
    532109.899393452, 563410.481710714, 594711.064027977, 626011.64634524, 
    657312.228662501, 688612.810979763, 719913.393297026, 751213.975614288, 
    782514.557931549, 813815.140248812, 845115.722566074, 876416.304883335, 
    907716.887200598, 939017.46951786, 970318.051835122, 1001618.63415238, 
    1032919.21646965, 1064219.79878691, 1095520.38110417, 1126820.96342143, 
    1158121.54573869, 1189422.12805596, 1220722.71037322, 1252023.29269048, 
    1283323.87500774, 1314624.45732501, 1345925.03964227, 1377225.62195953, 
    1408526.20427679, 1439826.78659405, 1471127.36891132, 1502427.95122858, 
    1533728.53354584, 1565029.1158631, 1596329.69818036, 1627630.28049763, 
    1658930.86281489, 1690231.44513215, 1721532.02744941,
  0, 31184.786230943, 62369.572461886, 93554.3586928317, 124739.144923777, 
    155923.93115472, 187108.717385666, 218293.503616612, 249478.289847555, 
    280663.0760785, 311847.862309446, 343032.648540389, 374217.434771335, 
    405402.22100228, 436587.007233224, 467771.793464169, 498956.579695115, 
    530141.365926058, 561326.152157002, 592510.938387948, 623695.724618894, 
    654880.510849838, 686065.297080782, 717250.083311728, 748434.869542672, 
    779619.655773617, 810804.442004562, 841989.228235507, 873174.014466451, 
    904358.800697397, 935543.586928341, 966728.373159286, 997913.159390231, 
    1029097.94562118, 1060282.73185212, 1091467.51808307, 1122652.30431401, 
    1153837.09054495, 1185021.8767759, 1216206.66300684, 1247391.44923779, 
    1278576.23546873, 1309761.02169968, 1340945.80793062, 1372130.59416157, 
    1403315.38039251, 1434500.16662346, 1465684.9528544, 1496869.73908535, 
    1528054.52531629, 1559239.31154724, 1590424.09777818, 1621608.88400913, 
    1652793.67024007, 1683978.45647102, 1715163.24270196,
  0, 31067.9346559707, 62135.8693119414, 93203.8039679147, 124271.738623888, 
    155339.673279859, 186407.607935832, 217475.542591805, 248543.477247776, 
    279611.411903749, 310679.346559723, 341747.281215693, 372815.215871667, 
    403883.15052764, 434951.085183611, 466019.019839584, 497086.954495557, 
    528154.889151528, 559222.8238075, 590290.758463474, 621358.693119447, 
    652426.627775419, 683494.562431391, 714562.497087364, 745630.431743336, 
    776698.366399308, 807766.301055282, 838834.235711254, 869902.170367226, 
    900970.105023199, 932038.039679171, 963105.974335143, 994173.908991117, 
    1025241.84364709, 1056309.77830306, 1087377.71295903, 1118445.64761501, 
    1149513.58227098, 1180581.51692695, 1211649.45158292, 1242717.3862389, 
    1273785.32089487, 1304853.25555084, 1335921.19020681, 1366989.12486279, 
    1398057.05951876, 1429124.99417473, 1460192.9288307, 1491260.86348668, 
    1522328.79814265, 1553396.73279862, 1584464.66745459, 1615532.60211056, 
    1646600.53676654, 1677668.47142251, 1708736.40607848,
  0, 30950.031547396, 61900.063094792, 92850.0946421907, 123800.126189589, 
    154750.157736985, 185700.189284384, 216650.220831783, 247600.252379179, 
    278550.283926577, 309500.315473976, 340450.347021372, 371400.378568771, 
    402350.410116169, 433300.441663565, 464250.473210964, 495200.504758363, 
    526150.536305759, 557100.567853156, 588050.599400555, 619000.630947953, 
    649950.662495351, 680900.694042748, 711850.725590147, 742800.757137544, 
    773750.788684941, 804700.82023234, 835650.851779737, 866600.883327135, 
    897550.914874533, 928500.946421931, 959450.977969328, 990401.009516727, 
    1021351.04106412, 1052301.07261152, 1083251.10415892, 1114201.13570632, 
    1145151.16725371, 1176101.19880111, 1207051.23034851, 1238001.26189591, 
    1268951.29344331, 1299901.3249907, 1330851.3565381, 1361801.3880855, 
    1392751.4196329, 1423701.45118029, 1454651.48272769, 1485601.51427509, 
    1516551.54582249, 1547501.57736989, 1578451.60891728, 1609401.64046468, 
    1640351.67201208, 1671301.70355948, 1702251.73510687,
  0, 30831.080895862, 61662.1617917241, 92493.2426875887, 123324.323583453, 
    154155.404479315, 184986.48537518, 215817.566271045, 246648.647166907, 
    277479.728062771, 308310.808958636, 339141.889854498, 369972.970750363, 
    400804.051646227, 431635.13254209, 462466.213437954, 493297.294333819, 
    524128.375229681, 554959.456125544, 585790.537021409, 616621.617917273, 
    647452.698813137, 678283.779709, 709114.860604865, 739945.941500728, 
    770777.022396591, 801608.103292456, 832439.184188319, 863270.265084183, 
    894101.345980047, 924932.426875911, 955763.507771774, 986594.588667639, 
    1017425.6695635, 1048256.75045937, 1079087.83135523, 1109918.91225109, 
    1140749.99314696, 1171581.07404282, 1202412.15493868, 1233243.23583455, 
    1264074.31673041, 1294905.39762628, 1325736.47852214, 1356567.559418, 
    1387398.64031387, 1418229.72120973, 1449060.80210559, 1479891.88300146, 
    1510722.96389732, 1541554.04479319, 1572385.12568905, 1603216.20658491, 
    1634047.28748078, 1664878.36837664, 1695709.4492725,
  0, 30711.086727467, 61422.173454934, 92133.2601824037, 122844.346909873, 
    153555.43363734, 184266.52036481, 214977.60709228, 245688.693819747, 
    276399.780547216, 307110.867274686, 337821.954002153, 368533.040729623, 
    399244.127457092, 429955.214184559, 460666.300912029, 491377.387639499, 
    522088.474366966, 552799.561094434, 583510.647821904, 614221.734549373, 
    644932.821276842, 675643.90800431, 706354.99473178, 737066.081459248, 
    767777.168186716, 798488.254914186, 829199.341641654, 859910.428369122, 
    890621.515096592, 921332.60182406, 952043.688551529, 982754.775278998, 
    1013465.86200647, 1044176.94873394, 1074888.0354614, 1105599.12218887, 
    1136310.20891634, 1167021.29564381, 1197732.38237128, 1228443.46909875, 
    1259154.55582622, 1289865.64255369, 1320576.72928115, 1351287.81600862, 
    1381998.90273609, 1412709.98946356, 1443421.07619103, 1474132.1629185, 
    1504843.24964597, 1535554.33637344, 1566265.4231009, 1596976.50982837, 
    1627687.59655584, 1658398.68328331, 1689109.77001078,
  0, 30590.0531036282, 61180.1062072564, 91770.1593108873, 122360.212414518, 
    152950.265518146, 183540.318621777, 214130.371725408, 244720.424829036, 
    275310.477932667, 305900.531036298, 336490.584139926, 367080.637243557, 
    397670.690347188, 428260.743450816, 458850.796554447, 489440.849658078, 
    520030.902761706, 550620.955865335, 581211.008968966, 611801.062072597, 
    642391.115176227, 672981.168279856, 703571.221383487, 734161.274487117, 
    764751.327590746, 795341.380694377, 825931.433798007, 856521.486901636, 
    887111.540005267, 917701.593108896, 948291.646212526, 978881.699316157, 
    1009471.75241979, 1040061.80552342, 1070651.85862705, 1101241.91173068, 
    1131831.96483431, 1162422.01793794, 1193012.07104157, 1223602.1241452, 
    1254192.17724883, 1284782.23035246, 1315372.28345609, 1345962.33655972, 
    1376552.38966335, 1407142.44276698, 1437732.49587061, 1468322.54897424, 
    1498912.60207787, 1529502.6551815, 1560092.70828512, 1590682.76138876, 
    1621272.81449239, 1651862.86759601, 1682452.92069964,
  0, 30467.9841209444, 60935.9682418887, 91403.9523628357, 121871.936483783, 
    152339.920604727, 182807.904725674, 213275.888846621, 243743.872967565, 
    274211.857088512, 304679.841209459, 335147.825330404, 365615.809451351, 
    396083.793572298, 426551.777693242, 457019.761814189, 487487.745935136, 
    517955.73005608, 548423.714177026, 578891.698297973, 609359.68241892, 
    639827.666539866, 670295.650660811, 700763.634781758, 731231.618902704, 
    761699.60302365, 792167.587144597, 822635.571265542, 853103.555386488, 
    883571.539507435, 914039.52362838, 944507.507749326, 974975.491870273, 
    1005443.47599122, 1035911.46011216, 1066379.44423311, 1096847.42835406, 
    1127315.412475, 1157783.39659595, 1188251.3807169, 1218719.36483784, 
    1249187.34895879, 1279655.33307973, 1310123.31720068, 1340591.30132163, 
    1371059.28544257, 1401527.26956352, 1431995.25368447, 1462463.23780541, 
    1492931.22192636, 1523399.2060473, 1553867.19016825, 1584335.1742892, 
    1614803.15841014, 1645271.14253109, 1675739.12665203,
  0, 30344.883911057, 60689.767822114, 91034.6517331736, 121379.535644233, 
    151724.41955529, 182069.30346635, 212414.187377409, 242759.071288466, 
    273103.955199526, 303448.839110585, 333793.723021642, 364138.606932702, 
    394483.490843762, 424828.374754819, 455173.258665878, 485518.142576938, 
    515863.026487995, 546207.910399053, 576552.794310113, 606897.678221172, 
    637242.56213223, 667587.446043289, 697932.329954348, 728277.213865407, 
    758622.097776465, 788966.981687525, 819311.865598583, 849656.749509641, 
    880001.633420701, 910346.517331759, 940691.401242817, 971036.285153877, 
    1001381.16906494, 1031726.05297599, 1062070.93688705, 1092415.82079811, 
    1122760.70470917, 1153105.58862023, 1183450.47253129, 1213795.35644235, 
    1244140.24035341, 1274485.12426446, 1304830.00817552, 1335174.89208658, 
    1365519.77599764, 1395864.6599087, 1426209.54381976, 1456554.42773082, 
    1486899.31164187, 1517244.19555293, 1547589.07946399, 1577933.96337505, 
    1608278.84728611, 1638623.73119717, 1668968.61510823,
  0, 30220.7566405106, 60441.5132810211, 90662.2699215342, 120883.026562047, 
    151103.783202558, 181324.539843071, 211545.296483584, 241766.053124095, 
    271986.809764608, 302207.566405121, 332428.323045632, 362649.079686145, 
    392869.836326658, 423090.592967168, 453311.349607682, 483532.106248195, 
    513752.862888705, 543973.619529217, 574194.37616973, 604415.132810243, 
    634635.889450755, 664856.646091267, 695077.40273178, 725298.159372292, 
    755518.916012804, 785739.672653317, 815960.429293829, 846181.185934341, 
    876401.942574854, 906622.699215366, 936843.455855877, 967064.212496391, 
    997284.969136902, 1027505.72577741, 1057726.48241793, 1087947.23905844, 
    1118167.99569895, 1148388.75233946, 1178609.50897998, 1208830.26562049, 
    1239051.022261, 1269271.77890151, 1299492.53554202, 1329713.29218254, 
    1359934.04882305, 1390154.80546356, 1420375.56210407, 1450596.31874459, 
    1480817.0753851, 1511037.83202561, 1541258.58866612, 1571479.34530663, 
    1601700.10194715, 1631920.85858766, 1662141.61522817,
  0, 30095.6065106115, 60191.2130212229, 90286.819531837, 120382.426042451, 
    150478.032553062, 180573.639063676, 210669.245574291, 240764.852084902, 
    270860.458595516, 300956.06510613, 331051.671616742, 361147.278127356, 
    391242.88463797, 421338.491148581, 451434.097659195, 481529.704169809, 
    511625.310680421, 541720.917191033, 571816.523701648, 601912.130212262, 
    632007.736722874, 662103.343233487, 692198.949744101, 722294.556254714, 
    752390.162765327, 782485.769275941, 812581.375786553, 842676.982297166, 
    872772.58880778, 902868.195318393, 932963.801829006, 963059.40833962, 
    993155.014850233, 1023250.62136085, 1053346.22787146, 1083441.83438207, 
    1113537.44089268, 1143633.0474033, 1173728.65391391, 1203824.26042452, 
    1233919.86693514, 1264015.47344575, 1294111.07995636, 1324206.68646698, 
    1354302.29297759, 1384397.8994882, 1414493.50599882, 1444589.11250943, 
    1474684.71902004, 1504780.32553066, 1534875.93204127, 1564971.53855188, 
    1595067.14506249, 1625162.75157311, 1655258.35808372,
  0, 29969.4377572858, 59938.8755145716, 89908.3132718599, 119877.751029148, 
    149847.188786434, 179816.626543722, 209786.064301011, 239755.502058297, 
    269724.939815585, 299694.377572873, 329663.815330159, 359633.253087447, 
    389602.690844736, 419572.128602021, 449541.56635931, 479511.004116598, 
    509480.441873884, 539449.879631171, 569419.317388459, 599388.755145748, 
    629358.192903035, 659327.630660322, 689297.06841761, 719266.506174897, 
    749235.943932184, 779205.381689473, 809174.81944676, 839144.257204047, 
    869113.694961335, 899083.132718622, 929052.570475909, 959022.008233197, 
    988991.445990485, 1018960.88374777, 1048930.32150506, 1078899.75926235, 
    1108869.19701963, 1138838.63477692, 1168808.07253421, 1198777.5102915, 
    1228746.94804879, 1258716.38580607, 1288685.82356336, 1318655.26132065, 
    1348624.69907794, 1378594.13683522, 1408563.57459251, 1438533.0123498, 
    1468502.45010709, 1498471.88786437, 1528441.32562166, 1558410.76337895, 
    1588380.20113624, 1618349.63889352, 1648319.07665081,
  0, 29842.2546509359, 59684.5093018719, 89526.7639528104, 119369.018603749, 
    149211.273254685, 179053.527905623, 208895.782556562, 238738.037207498, 
    268580.291858436, 298422.546509375, 328264.801160311, 358107.055811249, 
    387949.310462188, 417791.565113124, 447633.819764062, 477476.074415001, 
    507318.329065937, 537160.583716874, 567002.838367812, 596845.093018751, 
    626687.347669688, 656529.602320625, 686371.856971563, 716214.111622501, 
    746056.366273438, 775898.620924376, 805740.875575314, 835583.130226251, 
    865425.384877189, 895267.639528126, 925109.894179064, 954952.148830002, 
    984794.403480939, 1014636.65813188, 1044478.91278281, 1074321.16743375, 
    1104163.42208469, 1134005.67673563, 1163847.93138657, 1193690.1860375, 
    1223532.44068844, 1253374.69533938, 1283216.94999032, 1313059.20464125, 
    1342901.45929219, 1372743.71394313, 1402585.96859407, 1432428.223245, 
    1462270.47789594, 1492112.73254688, 1521954.98719782, 1551797.24184875, 
    1581639.49649969, 1611481.75115063, 1641324.00580157,
  0, 29714.061496296, 59428.1229925921, 89142.1844888906, 118856.245985189, 
    148570.307481485, 178284.368977784, 207998.430474082, 237712.491970378, 
    267426.553466677, 297140.614962975, 326854.676459272, 356568.73795557, 
    386282.799451869, 415996.860948165, 445710.922444463, 475424.983940762, 
    505139.045437058, 534853.106933355, 564567.168429654, 594281.229925952, 
    623995.29142225, 653709.352918547, 683423.414414845, 713137.475911143, 
    742851.53740744, 772565.598903738, 802279.660400036, 831993.721896333, 
    861707.783392631, 891421.844888929, 921135.906385226, 950849.967881524, 
    980564.029377822, 1010278.09087412, 1039992.15237042, 1069706.21386671, 
    1099420.27536301, 1129134.33685931, 1158848.39835561, 1188562.45985191, 
    1218276.5213482, 1247990.5828445, 1277704.6443408, 1307418.7058371, 
    1337132.76733339, 1366846.82882969, 1396560.89032599, 1426274.95182229, 
    1455989.01331858, 1485703.07481488, 1515417.13631118, 1545131.19780748, 
    1574845.25930378, 1604559.32080007, 1634273.38229637,
  0, 29584.8626322862, 59169.7252645724, 88754.5878968612, 118339.45052915, 
    147924.313161436, 177509.175793725, 207094.038426014, 236678.9010583, 
    266263.763690589, 295848.626322877, 325433.488955164, 355018.351587452, 
    384603.214219741, 414188.076852027, 443772.939484316, 473357.802116605, 
    502942.664748891, 532527.527381179, 562112.390013467, 591697.252645756, 
    621282.115278043, 650866.977910331, 680451.84054262, 710036.703174907, 
    739621.565807194, 769206.428439483, 798791.291071771, 828376.153704058, 
    857961.016336347, 887545.878968634, 917130.741600922, 946715.60423321, 
    976300.466865498, 1005885.32949779, 1035470.19213007, 1065055.05476236, 
    1094639.91739465, 1124224.78002694, 1153809.64265923, 1183394.50529151, 
    1212979.3679238, 1242564.23055609, 1272149.09318838, 1301733.95582066, 
    1331318.81845295, 1360903.68108524, 1390488.54371753, 1420073.40634982, 
    1449658.2689821, 1479243.13161439, 1508827.99424668, 1538412.85687897, 
    1567997.71951126, 1597582.58214354, 1627167.44477583,
  0, 29454.6624318658, 58909.3248637317, 88363.9872956, 117818.649727468, 
    147273.312159334, 176727.974591203, 206182.637023071, 235637.299454937, 
    265091.961886805, 294546.624318673, 324001.286750539, 353455.949182408, 
    382910.611614276, 412365.274046142, 441819.93647801, 471274.598909878, 
    500729.261341744, 530183.923773611, 559638.58620548, 589093.248637348, 
    618547.911069215, 648002.573501082, 677457.235932951, 706911.898364818, 
    736366.560796685, 765821.223228553, 795275.88566042, 824730.548092287, 
    854185.210524156, 883639.872956023, 913094.53538789, 942549.197819758, 
    972003.860251625, 1001458.52268349, 1030913.18511536, 1060367.84754723, 
    1089822.50997909, 1119277.17241096, 1148731.83484283, 1178186.4972747, 
    1207641.15970657, 1237095.82213843, 1266550.4845703, 1296005.14700217, 
    1325459.80943404, 1354914.4718659, 1384369.13429777, 1413823.79672964, 
    1443278.4591615, 1472733.12159337, 1502187.78402524, 1531642.44645711, 
    1561097.10888898, 1590551.77132084, 1620006.43375271,
  0, 29323.4653018853, 58646.9306037707, 87970.3959056585, 117293.861207546, 
    146617.326509432, 175940.791811319, 205264.257113207, 234587.722415093, 
    263911.18771698, 293234.653018868, 322558.118320754, 351881.583622641, 
    381205.048924529, 410528.514226415, 439851.979528302, 469175.44483019, 
    498498.910132076, 527822.375433962, 557145.84073585, 586469.306037738, 
    615792.771339624, 645116.236641511, 674439.701943399, 703763.167245285, 
    733086.632547172, 762410.09784906, 791733.563150946, 821057.028452833, 
    850380.493754721, 879703.959056607, 909027.424358494, 938350.889660382, 
    967674.354962268, 996997.820264155, 1026321.28556604, 1055644.75086793, 
    1084968.21616982, 1114291.6814717, 1143615.14677359, 1172938.61207548, 
    1202262.07737736, 1231585.54267925, 1260909.00798114, 1290232.47328303, 
    1319555.93858491, 1348879.4038868, 1378202.86918869, 1407526.33449057, 
    1436849.79979246, 1466173.26509435, 1495496.73039623, 1524820.19569812, 
    1554143.66100001, 1583467.1263019, 1612790.59160378,
  0, 29191.2756829371, 58382.5513658742, 87573.8270488138, 116765.102731753, 
    145956.378414691, 175147.65409763, 204338.92978057, 233530.205463507, 
    262721.481146446, 291912.756829386, 321104.032512323, 350295.308195263, 
    379486.583878202, 408677.85956114, 437869.135244079, 467060.410927019, 
    496251.686609956, 525442.962292894, 554634.237975834, 583825.513658773, 
    613016.789341712, 642208.06502465, 671399.34070759, 700590.616390528, 
    729781.892073467, 758973.167756406, 788164.443439345, 817355.719122283, 
    846546.994805222, 875738.270488161, 904929.546171099, 934120.821854039, 
    963312.097536977, 992503.373219916, 1021694.64890286, 1050885.92458579, 
    1080077.20026873, 1109268.47595167, 1138459.75163461, 1167651.02731755, 
    1196842.30300049, 1226033.57868343, 1255224.85436636, 1284416.1300493, 
    1313607.40573224, 1342798.68141518, 1371989.95709812, 1401181.23278106, 
    1430372.508464, 1459563.78414694, 1488755.05982987, 1517946.33551281, 
    1547137.61119575, 1576328.88687869, 1605520.16256163,
  0, 29058.0980492052, 58116.1960984105, 87174.2941476182, 116232.392196826, 
    145290.490246031, 174348.588295239, 203406.686344447, 232464.784393652, 
    261522.88244286, 290580.980492067, 319639.078541273, 348697.17659048, 
    377755.274639688, 406813.372688893, 435871.470738101, 464929.568787309, 
    493987.666836514, 523045.76488572, 552103.862934928, 581161.960984136, 
    610220.059033342, 639278.157082549, 668336.255131756, 697394.353180963, 
    726452.451230169, 755510.549279377, 784568.647328583, 813626.74537779, 
    842684.843426998, 871742.941476204, 900801.03952541, 929859.137574618, 
    958917.235623825, 987975.333673031, 1017033.43172224, 1046091.52977145, 
    1075149.62782065, 1104207.72586986, 1133265.82391907, 1162323.92196827, 
    1191382.02001748, 1220440.11806669, 1249498.21611589, 1278556.3141651, 
    1307614.41221431, 1336672.51026351, 1365730.60831272, 1394788.70636193, 
    1423846.80441113, 1452904.90246034, 1481963.00050955, 1511021.09855875, 
    1540079.19660796, 1569137.29465717, 1598195.39270637,
  0, 28923.9369083139, 57847.8738166279, 86771.8107249443, 115695.747633261, 
    144619.684541575, 173543.621449891, 202467.558358208, 231391.495266521, 
    260315.432174838, 289239.369083154, 318163.305991468, 347087.242899785, 
    376011.179808101, 404935.116716415, 433859.053624731, 462782.990533048, 
    491706.927441362, 520630.864349677, 549554.801257993, 578478.73816631, 
    607402.675074625, 636326.61198294, 665250.548891257, 694174.485799572, 
    723098.422707887, 752022.359616203, 780946.296524519, 809870.233432834, 
    838794.17034115, 867718.107249465, 896642.04415778, 925565.981066097, 
    954489.917974412, 983413.854882727, 1012337.79179104, 1041261.72869936, 
    1070185.66560767, 1099109.60251599, 1128033.53942431, 1156957.47633262, 
    1185881.41324094, 1214805.35014925, 1243729.28705757, 1272653.22396588, 
    1301577.1608742, 1330501.09778251, 1359425.03469083, 1388348.97159915, 
    1417272.90850746, 1446196.84541578, 1475120.78232409, 1504044.71923241, 
    1532968.65614072, 1561892.59304904, 1590816.52995735,
  0, 28788.7968011751, 57577.5936023502, 86366.3904035278, 115155.187204705, 
    143943.98400588, 172732.780807058, 201521.577608236, 230310.374409411, 
    259099.171210588, 287887.968011766, 316676.764812941, 345465.561614118, 
    374254.358415296, 403043.155216471, 431831.952017649, 460620.748818826, 
    489409.545620001, 518198.342421178, 546987.139222355, 575775.936023533, 
    604564.732824709, 633353.529625885, 662142.326427063, 690931.123228239, 
    719719.920029415, 748508.716830593, 777297.513631769, 806086.310432945, 
    834875.107234123, 863663.904035299, 892452.700836476, 921241.497637653, 
    950030.294438829, 978819.091240006, 1007607.88804118, 1036396.68484236, 
    1065185.48164354, 1093974.27844471, 1122763.07524589, 1151551.87204707, 
    1180340.66884824, 1209129.46564942, 1237918.2624506, 1266707.05925177, 
    1295495.85605295, 1324284.65285413, 1353073.4496553, 1381862.24645648, 
    1410651.04325766, 1439439.84005883, 1468228.63686001, 1497017.43366119, 
    1525806.23046236, 1554595.02726354, 1583383.82406472,
  0, 28652.6823018344, 57305.3646036689, 85958.0469055058, 114610.729207343, 
    143263.411509177, 171916.093811014, 200568.776112851, 229221.458414685, 
    257874.140716522, 286526.823018359, 315179.505320193, 343832.18762203, 
    372484.869923867, 401137.552225702, 429790.234527539, 458442.916829376, 
    487095.59913121, 515748.281433046, 544400.963734883, 573053.646036719, 
    601706.328338555, 630359.010640391, 659011.692942228, 687664.375244063, 
    716317.057545899, 744969.739847736, 773622.422149571, 802275.104451407, 
    830927.786753244, 859580.46905508, 888233.151356915, 916885.833658752, 
    945538.515960588, 974191.198262423, 1002843.88056426, 1031496.5628661, 
    1060149.24516793, 1088801.92746977, 1117454.6097716, 1146107.29207344, 
    1174759.97437528, 1203412.65667711, 1232065.33897895, 1260718.02128078, 
    1289370.70358262, 1318023.38588446, 1346676.06818629, 1375328.75048813, 
    1403981.43278996, 1432634.1150918, 1461286.79739364, 1489939.47969547, 
    1518592.16199731, 1547244.84429914, 1575897.52660098,
  0, 28515.5980173168, 57031.1960346336, 85546.7940519528, 114062.392069272, 
    142577.990086589, 171093.588103908, 199609.186121227, 228124.784138544, 
    256640.382155863, 285155.980173182, 313671.578190499, 342187.176207818, 
    370702.774225138, 399218.372242454, 427733.970259774, 456249.568277093, 
    484765.16629441, 513280.764311728, 541796.362329047, 570311.960346366, 
    598827.558363684, 627343.156381002, 655858.754398321, 684374.352415639, 
    712889.950432957, 741405.548450276, 769921.146467594, 798436.744484912, 
    826952.342502231, 855467.940519549, 883983.538536867, 912499.136554186, 
    941014.734571504, 969530.332588822, 998045.930606142, 1026561.52862346, 
    1055077.12664078, 1083592.7246581, 1112108.32267541, 1140623.92069273, 
    1169139.51871005, 1197655.11672737, 1226170.71474469, 1254686.31276201, 
    1283201.91077932, 1311717.50879664, 1340233.10681396, 1368748.70483128, 
    1397264.3028486, 1425779.90086592, 1454295.49888323, 1482811.09690055, 
    1511326.69491787, 1539842.29293519, 1568357.89095251,
  0, 28377.5485874701, 56755.0971749401, 85132.6457624126, 113510.194349885, 
    141887.742937355, 170265.291524828, 198642.8401123, 227020.38869977, 
    255397.937287243, 283775.485874715, 312153.034462185, 340530.583049658, 
    368908.13163713, 397285.6802246, 425663.228812073, 454040.777399545, 
    482418.325987015, 510795.874574487, 539173.423161959, 567550.971749432, 
    595928.520336903, 624306.068924374, 652683.617511847, 681061.166099318, 
    709438.714686789, 737816.263274262, 766193.811861733, 794571.360449204, 
    822948.909036677, 851326.457624148, 879704.006211619, 908081.554799092, 
    936459.103386563, 964836.651974034, 993214.200561507, 1021591.74914898, 
    1049969.29773645, 1078346.84632392, 1106724.39491139, 1135101.94349886, 
    1163479.49208634, 1191857.04067381, 1220234.58926128, 1248612.13784875, 
    1276989.68643622, 1305367.23502369, 1333744.78361117, 1362122.33219864, 
    1390499.88078611, 1418877.42937358, 1447254.97796105, 1475632.52654852, 
    1504010.075136, 1532387.62372347, 1560765.17231094,
  0, 28238.5386848083, 56477.0773696166, 84715.6160544273, 112954.154739238, 
    141192.693424046, 169431.232108857, 197669.770793668, 225908.309478476, 
    254146.848163287, 282385.386848097, 310623.925532906, 338862.464217716, 
    367101.002902527, 395339.541587335, 423578.080272146, 451816.618956957, 
    480055.157641765, 508293.696326574, 536532.235011385, 564770.773696196, 
    593009.312381005, 621247.851065815, 649486.389750626, 677724.928435435, 
    705963.467120245, 734202.005805055, 762440.544489865, 790679.083174674, 
    818917.621859485, 847156.160544294, 875394.699229104, 903633.237913915, 
    931871.776598724, 960110.315283534, 988348.853968344, 1016587.39265315, 
    1044825.93133796, 1073064.47002277, 1101303.00870758, 1129541.54739239, 
    1157780.0860772, 1186018.62476201, 1214257.16344682, 1242495.70213163, 
    1270734.24081644, 1298972.77950125, 1327211.31818606, 1355449.85687087, 
    1383688.39555568, 1411926.93424049, 1440165.4729253, 1468404.01161011, 
    1496642.55029492, 1524881.08897973, 1553119.62766454,
  0, 28098.5730143534, 56197.1460287067, 84295.7190430625, 112394.292057418, 
    140492.865071772, 168591.438086127, 196690.011100483, 224788.584114836, 
    252887.157129192, 280985.730143548, 309084.303157901, 337182.876172257, 
    365281.449186613, 393380.022200966, 421478.595215322, 449577.168229678, 
    477675.741244031, 505774.314258385, 533872.887272741, 561971.460287097, 
    590070.033301451, 618168.606315806, 646267.179330162, 674365.752344516, 
    702464.325358871, 730562.898373227, 758661.471387581, 786760.044401936, 
    814858.617416291, 842957.190430646, 871055.763445001, 899154.336459356, 
    927252.909473711, 955351.482488065, 983450.055502421, 1011548.62851678, 
    1039647.20153113, 1067745.77454549, 1095844.34755984, 1123942.9205742, 
    1152041.49358855, 1180140.06660291, 1208238.63961726, 1236337.21263162, 
    1264435.78564597, 1292534.35866032, 1320632.93167468, 1348731.50468904, 
    1376830.07770339, 1404928.65071774, 1433027.2237321, 1461125.79674645, 
    1489224.36976081, 1517322.94277516, 1545421.51578952,
  0, 27957.6563134758, 55915.3126269515, 83872.9689404297, 111830.625253908, 
    139788.281567384, 167745.937880862, 195703.59419434, 223661.250507816, 
    251618.906821294, 279576.563134772, 307534.219448248, 335491.875761726, 
    363449.532075204, 391407.18838868, 419364.844702158, 447322.501015636, 
    475280.157329112, 503237.813642589, 531195.469956067, 559153.126269545, 
    587110.782583022, 615068.438896499, 643026.095209977, 670983.751523454, 
    698941.407836931, 726899.064150409, 754856.720463886, 782814.376777363, 
    810772.033090841, 838729.689404318, 866687.345717795, 894645.002031273, 
    922602.65834475, 950560.314658227, 978517.970971706, 1006475.62728518, 
    1034433.28359866, 1062390.93991214, 1090348.59622561, 1118306.25253909, 
    1146263.90885257, 1174221.56516605, 1202179.22147952, 1230136.877793, 
    1258094.53410648, 1286052.19041996, 1314009.84673343, 1341967.50304691, 
    1369925.15936039, 1397882.81567386, 1425840.47198734, 1453798.12830082, 
    1481755.7846143, 1509713.44092777, 1537671.09724125,
  0, 27815.7933517344, 55631.5867034687, 83447.3800552054, 111263.173406942, 
    139078.966758677, 166894.760110413, 194710.55346215, 222526.346813884, 
    250342.140165621, 278157.933517358, 305973.726869092, 333789.520220829, 
    361605.313572566, 389421.1069243, 417236.900276037, 445052.693627773, 
    472868.486979508, 500684.280331243, 528500.07368298, 556315.867034717, 
    584131.660386452, 611947.453738188, 639763.247089925, 667579.04044166, 
    695394.833793396, 723210.627145133, 751026.420496868, 778842.213848604, 
    806658.00720034, 834473.800552076, 862289.593903812, 890105.387255548, 
    917921.180607284, 945736.973959019, 973552.767310756, 1001368.56066249, 
    1029184.35401423, 1057000.14736596, 1084815.9407177, 1112631.73406943, 
    1140447.52742117, 1168263.32077291, 1196079.11412464, 1223894.90747638, 
    1251710.70082811, 1279526.49417985, 1307342.28753159, 1335158.08088332, 
    1362973.87423506, 1390789.66758679, 1418605.46093853, 1446421.25429027, 
    1474237.047642, 1502052.84099374, 1529868.63434547,
  0, 27672.9889307147, 55345.9778614295, 83018.9667921466, 110691.955722864, 
    138364.944653578, 166037.933584296, 193710.922515013, 221383.911445727, 
    249056.900376444, 276729.889307162, 304402.878237876, 332075.867168593, 
    359748.856099311, 387421.845030025, 415094.833960742, 442767.822891459, 
    470440.811822174, 498113.80075289, 525786.789683607, 553459.778614324, 
    581132.76754504, 608805.756475756, 636478.745406473, 664151.734337189, 
    691824.723267905, 719497.712198622, 747170.701129338, 774843.690060054, 
    802516.678990771, 830189.667921487, 857862.656852203, 885535.64578292, 
    913208.634713636, 940881.623644352, 968554.612575069, 996227.601505785, 
    1023900.5904365, 1051573.57936722, 1079246.56829793, 1106919.55722865, 
    1134592.54615937, 1162265.53509008, 1189938.5240208, 1217611.51295152, 
    1245284.50188223, 1272957.49081295, 1300630.47974367, 1328303.46867438, 
    1355976.4576051, 1383649.44653581, 1411322.43546653, 1438995.42439725, 
    1466668.41332796, 1494341.40225868, 1522014.39118939,
  0, 27529.2478838669, 55058.4957677337, 82587.7436516029, 110116.991535472, 
    137646.239419339, 165175.487303208, 192704.735187077, 220233.983070944, 
    247763.230954813, 275292.478838683, 302821.726722549, 330350.974606419, 
    357880.222490288, 385409.470374155, 412938.718258024, 440467.966141893, 
    467997.21402576, 495526.461909628, 523055.709793497, 550584.957677366, 
    578114.205561234, 605643.453445103, 633172.701328972, 660701.94921284, 
    688231.197096708, 715760.444980577, 743289.692864445, 770818.940748313, 
    798348.188632182, 825877.43651605, 853406.684399919, 880935.932283788, 
    908465.180167656, 935994.428051524, 963523.675935393, 991052.923819261, 
    1018582.17170313, 1046111.419587, 1073640.66747087, 1101169.91535473, 
    1128699.1632386, 1156228.41112247, 1183757.65900634, 1211286.90689021, 
    1238816.15477408, 1266345.40265794, 1293874.65054181, 1321403.89842568, 
    1348933.14630955, 1376462.39419342, 1403991.64207729, 1431520.88996115, 
    1459050.13784502, 1486579.38572889, 1514108.63361276,
  0, 27384.5750763413, 54769.1501526826, 82153.7252290263, 109538.30030537, 
    136922.875381711, 164307.450458055, 191692.025534398, 219076.60061074, 
    246461.175687083, 273845.750763427, 301230.325839768, 328614.900916112, 
    355999.475992456, 383384.051068797, 410768.626145141, 438153.201221484, 
    465537.776297825, 492922.351374168, 520306.926450511, 547691.501526855, 
    575076.076603198, 602460.65167954, 629845.226755884, 657229.801832226, 
    684614.376908569, 711998.951984912, 739383.527061255, 766768.102137597, 
    794152.677213941, 821537.252290283, 848921.827366626, 876306.402442969, 
    903690.977519312, 931075.552595654, 958460.127671998, 985844.70274834, 
    1013229.27782468, 1040613.85290103, 1067998.42797737, 1095383.00305371, 
    1122767.57813005, 1150152.1532064, 1177536.72828274, 1204921.30335908, 
    1232305.87843543, 1259690.45351177, 1287075.02858811, 1314459.60366446, 
    1341844.1787408, 1369228.75381714, 1396613.32889348, 1423997.90396983, 
    1451382.47904617, 1478767.05412251, 1506151.62919885,
  0, 27238.9754048247, 54477.9508096494, 81716.9262144765, 108955.901619303, 
    136194.877024128, 163433.852428955, 190672.827833782, 217911.803238607, 
    245150.778643434, 272389.754048261, 299628.729453086, 326867.704857913, 
    354106.68026274, 381345.655667565, 408584.631072392, 435823.606477219, 
    463062.581882043, 490301.557286869, 517540.532691696, 544779.508096523, 
    572018.483501349, 599257.458906175, 626496.434311002, 653735.409715828, 
    680974.385120654, 708213.360525481, 735452.335930307, 762691.311335133, 
    789930.28673996, 817169.262144785, 844408.237549611, 871647.212954438, 
    898886.188359264, 926125.16376409, 953364.139168917, 980603.114573743, 
    1007842.08997857, 1035081.0653834, 1062320.04078822, 1089559.01619305, 
    1116797.99159787, 1144036.9670027, 1171275.94240753, 1198514.91781235, 
    1225753.89321718, 1252992.868622, 1280231.84402683, 1307470.81943166, 
    1334709.79483648, 1361948.77024131, 1389187.74564614, 1416426.72105096, 
    1443665.69645579, 1470904.67186061, 1498143.64726544,
  0, 27092.453797374, 54184.9075947479, 81277.3613921242, 108369.8151895, 
    135462.268986874, 162554.722784251, 189647.176581627, 216739.630379001, 
    243832.084176377, 270924.537973753, 298016.991771127, 325109.445568504, 
    352201.89936588, 379294.353163254, 406386.80696063, 433479.260758006, 
    460571.71455538, 487664.168352755, 514756.622150132, 541849.075947508, 
    568941.529744883, 596033.983542258, 623126.437339634, 650218.891137009, 
    677311.344934385, 704403.798731761, 731496.252529136, 758588.706326511, 
    785681.160123887, 812773.613921262, 839866.067718637, 866958.521516014, 
    894050.975313389, 921143.429110764, 948235.88290814, 975328.336705515, 
    1002420.79050289, 1029513.24430027, 1056605.69809764, 1083698.15189502, 
    1110790.60569239, 1137883.05948977, 1164975.51328714, 1192067.96708452, 
    1219160.42088189, 1246252.87467927, 1273345.32847665, 1300437.78227402, 
    1327530.2360714, 1354622.68986877, 1381715.14366615, 1408807.59746352, 
    1435900.0512609, 1462992.50505827, 1490084.95885565,
  0, 26945.0152132493, 53890.0304264987, 80835.0456397503, 107780.060853002, 
    134725.076066251, 161670.091279503, 188615.106492755, 215560.121706004, 
    242505.136919256, 269450.152132507, 296395.167345757, 323340.182559008, 
    350285.19777226, 377230.212985509, 404175.228198761, 431120.243412013, 
    458065.258625262, 485010.273838512, 511955.289051764, 538900.304265016, 
    565845.319478266, 592790.334691517, 619735.349904768, 646680.365118019, 
    673625.380331269, 700570.395544521, 727515.410757772, 754460.425971022, 
    781405.441184274, 808350.456397524, 835295.471610775, 862240.486824027, 
    889185.502037277, 916130.517250528, 943075.532463779, 970020.54767703, 
    996965.562890281, 1023910.57810353, 1050855.59331678, 1077800.60853003, 
    1104745.62374328, 1131690.63895654, 1158635.65416979, 1185580.66938304, 
    1212525.68459629, 1239470.69980954, 1266415.71502279, 1293360.73023604, 
    1320305.74544929, 1347250.76066254, 1374195.77587579, 1401140.79108904, 
    1428085.80630229, 1455030.82151554, 1481975.83672879,
  0, 26796.6646427468, 53593.3292854935, 80389.9939282426, 107186.658570992, 
    133983.323213738, 160779.987856487, 187576.652499237, 214373.317141983, 
    241169.981784732, 267966.646427481, 294763.311070228, 321559.975712977, 
    348356.640355726, 375153.304998473, 401949.969641222, 428746.634283971, 
    455543.298926718, 482339.963569466, 509136.628212215, 535933.292854964, 
    562729.957497712, 589526.62214046, 616323.286783209, 643119.951425957, 
    669916.616068705, 696713.280711454, 723509.945354202, 750306.60999695, 
    777103.274639699, 803899.939282447, 830696.603925195, 857493.268567944, 
    884289.933210692, 911086.59785344, 937883.262496189, 964679.927138937, 
    991476.591781685, 1018273.25642443, 1045069.92106718, 1071866.58570993, 
    1098663.25035268, 1125459.91499543, 1152256.57963817, 1179053.24428092, 
    1205849.90892367, 1232646.57356642, 1259443.23820917, 1286239.90285192, 
    1313036.56749466, 1339833.23213741, 1366629.89678016, 1393426.56142291, 
    1420223.22606566, 1447019.89070841, 1473816.55535115,
  0, 26647.4071070288, 53294.8142140576, 79942.2213210886, 106589.62842812, 
    133237.035535148, 159884.44264218, 186531.849749211, 213179.256856239, 
    239826.66396327, 266474.071070302, 293121.47817733, 319768.885284361, 
    346416.292391393, 373063.699498421, 399711.106605452, 426358.513712483, 
    453005.920819512, 479653.327926542, 506300.735033573, 532948.142140604, 
    559595.549247634, 586242.956354664, 612890.363461695, 639537.770568725, 
    666185.177675755, 692832.584782786, 719479.991889816, 746127.398996846, 
    772774.806103877, 799422.213210907, 826069.620317937, 852717.027424968, 
    879364.434531998, 906011.841639028, 932659.248746059, 959306.655853089, 
    985954.062960119, 1012601.47006715, 1039248.87717418, 1065896.28428121, 
    1092543.69138824, 1119191.09849527, 1145838.5056023, 1172485.91270933, 
    1199133.31981636, 1225780.72692339, 1252428.13403042, 1279075.54113745, 
    1305722.94824448, 1332370.35535151, 1359017.76245854, 1385665.16956557, 
    1412312.5766726, 1438959.98377963, 1465607.39088666,
  0, 26497.2476579546, 52994.4953159093, 79491.7429738661, 105988.990631823, 
    132486.238289778, 158983.485947735, 185480.733605691, 211977.981263646, 
    238475.228921603, 264972.47657956, 291469.724237515, 317966.971895471, 
    344464.219553428, 370961.467211383, 397458.71486934, 423955.962527297, 
    450453.210185251, 476950.457843207, 503447.705501164, 529944.953159121, 
    556442.200817077, 582939.448475032, 609436.696132989, 635933.943790945, 
    662431.191448901, 688928.439106858, 715425.686764813, 741922.934422769, 
    768420.182080726, 794917.429738682, 821414.677396638, 847911.925054595, 
    874409.17271255, 900906.420370506, 927403.668028463, 953900.915686419, 
    980398.163344374, 1006895.41100233, 1033392.65866029, 1059889.90631824, 
    1086387.1539762, 1112884.40163416, 1139381.64929211, 1165878.89695007, 
    1192376.14460802, 1218873.39226598, 1245370.63992394, 1271867.88758189, 
    1298365.13523985, 1324862.3828978, 1351359.63055576, 1377856.87821372, 
    1404354.12587167, 1430851.37352963, 1457348.62118758,
  0, 26346.1913779092, 52692.3827558185, 79038.57413373, 105384.765511641, 
    131730.956889551, 158077.148267462, 184423.339645374, 210769.531023283, 
    237115.722401194, 263461.913779106, 289808.105157015, 316154.296534927, 
    342500.487912838, 368846.679290747, 395192.870668659, 421539.06204657, 
    447885.253424479, 474231.44480239, 500577.636180301, 526923.827558213, 
    553270.018936123, 579616.210314033, 605962.401691945, 632308.593069855, 
    658654.784447766, 685000.975825677, 711347.167203587, 737693.358581498, 
    764039.549959409, 790385.741337319, 816731.93271523, 843078.124093141, 
    869424.315471052, 895770.506848962, 922116.698226873, 948462.889604784, 
    974809.080982694, 1001155.27236061, 1027501.46373852, 1053847.65511643, 
    1080193.84649434, 1106540.03787225, 1132886.22925016, 1159232.42062807, 
    1185578.61200598, 1211924.80338389, 1238270.9947618, 1264617.18613971, 
    1290963.37751762, 1317309.56889553, 1343655.76027344, 1370001.95165136, 
    1396348.14302927, 1422694.33440718, 1449040.52578509,
  0, 26194.2433796312, 52388.4867592624, 78582.7301388959, 104776.973518529, 
    130971.216898161, 157165.460277794, 183359.703657428, 209553.947037059, 
    235748.190416692, 261942.433796326, 288136.677175957, 314330.92055559, 
    340525.163935224, 366719.407314855, 392913.650694488, 419107.894074122, 
    445302.137453753, 471496.380833386, 497690.624213019, 523884.867592652, 
    550079.110972285, 576273.354351917, 602467.597731551, 628661.841111183, 
    654856.084490815, 681050.327870449, 707244.571250081, 733438.814629713, 
    759633.058009347, 785827.301388979, 812021.544768612, 838215.788148245, 
    864410.031527877, 890604.27490751, 916798.518287143, 942992.761666775, 
    969187.005046408, 995381.248426041, 1021575.49180567, 1047769.73518531, 
    1073963.97856494, 1100158.22194457, 1126352.4653242, 1152546.70870384, 
    1178740.95208347, 1204935.1954631, 1231129.43884274, 1257323.68222237, 
    1283517.925602, 1309712.16898163, 1335906.41236126, 1362100.6557409, 
    1388294.89912053, 1414489.14250016, 1440683.3858798,
  0, 26041.4088060398, 52082.8176120796, 78124.2264181216, 104165.635224164, 
    130207.044030203, 156248.452836245, 182289.861642287, 208331.270448327, 
    234372.679254369, 260414.088060411, 286455.496866451, 312496.905672493, 
    338538.314478535, 364579.723284575, 390621.132090617, 416662.540896659, 
    442703.949702698, 468745.358508739, 494786.767314781, 520828.176120823, 
    546869.584926864, 572910.993732905, 598952.402538947, 624993.811344988, 
    651035.220151029, 677076.628957071, 703118.037763112, 729159.446569153, 
    755200.855375195, 781242.264181236, 807283.672987276, 833325.081793319, 
    859366.490599359, 885407.8994054, 911449.308211442, 937490.717017483, 
    963532.125823524, 989573.534629566, 1015614.94343561, 1041656.35224165, 
    1067697.76104769, 1093739.16985373, 1119780.57865977, 1145821.98746581, 
    1171863.39627185, 1197904.8050779, 1223946.21388394, 1249987.62268998, 
    1276029.03149602, 1302070.44030206, 1328111.8491081, 1354153.25791414, 
    1380194.66672018, 1406236.07552623, 1432277.48433227,
  0, 25887.6928300606, 51775.3856601213, 77663.0784901841, 103550.771320247, 
    129438.464150308, 155326.15698037, 181213.849810433, 207101.542640494, 
    232989.235470557, 258876.92830062, 284764.62113068, 310652.313960743, 
    336540.006790806, 362427.699620867, 388315.392450929, 414203.085280992, 
    440090.778111053, 465978.470941115, 491866.163771177, 517753.85660124, 
    543641.549431302, 569529.242261364, 595416.935091426, 621304.627921488, 
    647192.32075155, 673080.013581613, 698967.706411675, 724855.399241736, 
    750743.092071799, 776630.784901861, 802518.477731923, 828406.170561986, 
    854293.863392047, 880181.556222109, 906069.249052172, 931956.941882234, 
    957844.634712295, 983732.327542358, 1009620.02037242, 1035507.71320248, 
    1061395.40603254, 1087283.09886261, 1113170.79169267, 1139058.48452273, 
    1164946.17735279, 1190833.87018285, 1216721.56301292, 1242609.25584298, 
    1268496.94867304, 1294384.6415031, 1320272.33433317, 1346160.02716323, 
    1372047.71999329, 1397935.41282335, 1423823.10565341,
  0, 25733.1006544509, 51466.2013089019, 77199.301963355, 102932.402617808, 
    128665.503272259, 154398.603926712, 180131.704581165, 205864.805235616, 
    231597.905890069, 257331.006544523, 283064.107198973, 308797.207853427, 
    334530.30850788, 360263.409162331, 385996.509816784, 411729.610471237, 
    437462.711125688, 463195.81178014, 488928.912434593, 514662.013089046, 
    540395.113743498, 566128.21439795, 591861.315052403, 617594.415706855, 
    643327.516361307, 669060.617015761, 694793.717670213, 720526.818324665, 
    746259.918979118, 771993.01963357, 797726.120288022, 823459.220942475, 
    849192.321596927, 874925.422251379, 900658.522905832, 926391.623560284, 
    952124.724214736, 977857.824869189, 1003590.92552364, 1029324.02617809, 
    1055057.12683255, 1080790.227487, 1106523.32814145, 1132256.4287959, 
    1157989.52945036, 1183722.63010481, 1209455.73075926, 1235188.83141371, 
    1260921.93206816, 1286655.03272262, 1312388.13337707, 1338121.23403152, 
    1363854.33468597, 1389587.43534043, 1415320.53599488,
  0, 25577.6375116231, 51155.2750232462, 76732.9125348715, 102310.550046497, 
    127888.18755812, 153465.825069745, 179043.462581371, 204621.100092994, 
    230198.737604619, 255776.375116244, 281354.012627867, 306931.650139493, 
    332509.287651118, 358086.925162741, 383664.562674366, 409242.200185992, 
    434819.837697615, 460397.475209239, 485975.112720864, 511552.75023249, 
    537130.387744114, 562708.025255738, 588285.662767363, 613863.300278988, 
    639440.937790612, 665018.575302237, 690596.212813861, 716173.850325486, 
    741751.487837111, 767329.125348735, 792906.76286036, 818484.400371985, 
    844062.037883609, 869639.675395233, 895217.312906859, 920794.950418483, 
    946372.587930107, 971950.225441732, 997527.862953357, 1023105.50046498, 
    1048683.13797661, 1074260.77548823, 1099838.41299985, 1125416.05051148, 
    1150993.6880231, 1176571.32553473, 1202148.96304635, 1227726.60055798, 
    1253304.2380696, 1278881.87558123, 1304459.51309285, 1330037.15060448, 
    1355614.7881161, 1381192.42562773, 1406770.06313935,
  0, 25421.3086634678, 50842.6173269357, 76263.9259904057, 101685.234653876, 
    127106.543317344, 152527.851980814, 177949.160644284, 203370.469307751, 
    228791.777971221, 254213.086634692, 279634.395298159, 305055.703961629, 
    330477.012625099, 355898.321288567, 381319.629952037, 406740.938615507, 
    432162.247278975, 457583.555942444, 483004.864605914, 508426.173269384, 
    533847.481932853, 559268.790596322, 584690.099259792, 610111.407923261, 
    635532.71658673, 660954.0252502, 686375.333913669, 711796.642577138, 
    737217.951240608, 762639.259904077, 788060.568567546, 813481.877231015, 
    838903.185894484, 864324.494557953, 889745.803221423, 915167.111884892, 
    940588.420548361, 966009.729211831, 991431.0378753, 1016852.34653877, 
    1042273.65520224, 1067694.96386571, 1093116.27252918, 1118537.58119265, 
    1143958.88985612, 1169380.19851958, 1194801.50718305, 1220222.81584652, 
    1245644.12450999, 1271065.43317346, 1296486.74183693, 1321908.0505004, 
    1347329.35916387, 1372750.66782734, 1398171.97649081,
  0, 25264.1194011759, 50528.2388023518, 75792.3582035298, 101056.477604708, 
    126320.597005884, 151584.716407062, 176848.83580824, 202112.955209416, 
    227377.074610594, 252641.194011772, 277905.313412948, 303169.432814126, 
    328433.552215304, 353697.67161648, 378961.791017658, 404225.910418836, 
    429490.029820012, 454754.149221189, 480018.268622367, 505282.388023545, 
    530546.507424721, 555810.626825898, 581074.746227077, 606338.865628253, 
    631602.98502943, 656867.104430608, 682131.223831785, 707395.343232962, 
    732659.46263414, 757923.582035317, 783187.701436494, 808451.820837672, 
    833715.940238849, 858980.059640026, 884244.179041204, 909508.298442381, 
    934772.417843558, 960036.537244736, 985300.656645913, 1010564.77604709, 
    1035828.89544827, 1061093.01484945, 1086357.13425062, 1111621.2536518, 
    1136885.37305298, 1162149.49245415, 1187413.61185533, 1212677.73125651, 
    1237941.85065769, 1263205.97005886, 1288470.08946004, 1313734.20886122, 
    1338998.3282624, 1364262.44766357, 1389526.56706475,
  0, 25106.075045059, 50212.150090118, 75318.2251351791, 100424.30018024, 
    125530.375225299, 150636.45027036, 175742.525315422, 200848.600360481, 
    225954.675405542, 251060.750450603, 276166.825495662, 301272.900540723, 
    326378.975585784, 351485.050630843, 376591.125675904, 401697.200720965, 
    426803.275766024, 451909.350811084, 477015.425856145, 502121.500901207, 
    527227.575946267, 552333.650991327, 577439.726036388, 602545.801081448, 
    627651.876126508, 652757.951171569, 677864.026216629, 702970.101261689, 
    728076.17630675, 753182.25135181, 778288.32639687, 803394.401441931, 
    828500.476486991, 853606.551532051, 878712.626577113, 903818.701622173, 
    928924.776667233, 954030.851712294, 979136.926757354, 1004243.00180241, 
    1029349.07684748, 1054455.15189254, 1079561.2269376, 1104667.30198266, 
    1129773.37702772, 1154879.45207278, 1179985.52711784, 1205091.6021629, 
    1230197.67720796, 1255303.75225302, 1280409.82729808, 1305515.90234314, 
    1330621.9773882, 1355728.05243326, 1380834.12747832,
  0, 24947.1809443698, 49894.3618887396, 74841.5428331116, 99788.7237774835, 
    124735.904721853, 149683.085666225, 174630.266610597, 199577.447554967, 
    224524.628499339, 249471.809443711, 274418.990388081, 299366.171332453, 
    324313.352276825, 349260.533221194, 374207.714165566, 399154.895109938, 
    424102.076054308, 449049.256998679, 473996.437943051, 498943.618887423, 
    523890.799831794, 548837.980776165, 573785.161720537, 598732.342664908, 
    623679.523609278, 648626.70455365, 673573.885498021, 698521.066442392, 
    723468.247386764, 748415.428331135, 773362.609275506, 798309.790219878, 
    823256.971164249, 848204.15210862, 873151.333052992, 898098.513997363, 
    923045.694941734, 947992.875886106, 972940.056830477, 997887.237774848, 
    1022834.41871922, 1047781.59966359, 1072728.78060796, 1097675.96155233, 
    1122623.1424967, 1147570.32344107, 1172517.50438545, 1197464.68532982, 
    1222411.86627419, 1247359.04721856, 1272306.22816293, 1297253.4091073, 
    1322200.59005167, 1347147.77099604, 1372094.95194042,
  0, 24787.4424771209, 49574.8849542418, 74362.3274313648, 99149.7699084878, 
    123937.212385609, 148724.654862732, 173512.097339855, 198299.539816976, 
    223086.982294099, 247874.424771222, 272661.867248342, 297449.309725465, 
    322236.752202588, 347024.194679709, 371811.637156832, 396599.079633955, 
    421386.522111076, 446173.964588198, 470961.407065321, 495748.849542444, 
    520536.292019566, 545323.734496688, 570111.176973811, 594898.619450933, 
    619686.061928055, 644473.504405178, 669260.9468823, 694048.389359422, 
    718835.831836545, 743623.274313667, 768410.716790789, 793198.159267912, 
    817985.601745034, 842773.044222156, 867560.486699279, 892347.929176401, 
    917135.371653522, 941922.814130645, 966710.256607767, 991497.699084889, 
    1016285.14156201, 1041072.58403913, 1065860.02651626, 1090647.46899338, 
    1115434.9114705, 1140222.35394762, 1165009.79642475, 1189797.23890187, 
    1214584.68137899, 1239372.12385611, 1264159.56633323, 1288947.00881036, 
    1313734.45128748, 1338521.8937646, 1363309.33624172 ;

 x_u =
  16040.6382749892, 48121.9148249677, 80203.1913749475, 112284.467924929, 
    144365.744474909, 176447.021024888, 208528.297574869, 240609.574124849, 
    272690.850674829, 304772.12722481, 336853.40377479, 368934.68032477, 
    401015.956874751, 433097.233424731, 465178.509974711, 497259.786524692, 
    529341.063074672, 561422.339624651, 593503.616174632, 625584.892724613, 
    657666.169274593, 689747.445824573, 721828.722374554, 753909.998924534, 
    785991.275474514, 818072.552024494, 850153.828574475, 882235.105124455, 
    914316.381674435, 946397.658224416, 978478.934774396, 1010560.21132438, 
    1042641.48787436, 1074722.76442434, 1106804.04097432, 1138885.3175243, 
    1170966.59407428, 1203047.87062426, 1235129.14717424, 1267210.42372422, 
    1299291.7002742, 1331372.97682418, 1363454.25337416, 1395535.52992414, 
    1427616.80647412, 1459698.0830241, 1491779.35957408, 1523860.63612406, 
    1555941.91267404, 1588023.18922402, 1620104.465774, 1652185.74232398, 
    1684267.01887396, 1716348.29542394, 1748429.57197392,
  15986.4883041619, 47959.4649124858, 79932.441520811, 111905.418129138, 
    143878.394737463, 175851.371345788, 207824.347954115, 239797.32456244, 
    271770.301170765, 303743.277779092, 335716.254387417, 367689.230995742, 
    399662.207604069, 431635.184212394, 463608.160820719, 495581.137429046, 
    527554.114037371, 559527.090645695, 591500.067254021, 623473.043862348, 
    655446.020470674, 687418.997078999, 719391.973687325, 751364.950295651, 
    783337.926903976, 815310.903512302, 847283.880120628, 879256.856728953, 
    911229.833337279, 943202.809945605, 975175.78655393, 1007148.76316226, 
    1039121.73977058, 1071094.71637891, 1103067.69298723, 1135040.66959556, 
    1167013.64620388, 1198986.62281221, 1230959.59942054, 1262932.57602886, 
    1294905.55263719, 1326878.52924551, 1358851.50585384, 1390824.48246216, 
    1422797.45907049, 1454770.43567882, 1486743.41228714, 1518716.38889547, 
    1550689.36550379, 1582662.34211212, 1614635.31872044, 1646608.29532877, 
    1678581.2719371, 1710554.24854542, 1742527.22515375,
  15931.797250134, 47795.391750402, 79658.9862506714, 111522.580750942, 
    143386.175251211, 175249.769751481, 207113.364251752, 238976.958752021, 
    270840.55325229, 302704.147752561, 334567.74225283, 366431.3367531, 
    398294.93125337, 430158.52575364, 462022.120253909, 493885.71475418, 
    525749.309254449, 557612.903754718, 589476.498254988, 621340.092755259, 
    653203.687255529, 685067.281755798, 716930.876256068, 748794.470756338, 
    780658.065256607, 812521.659756878, 844385.254257148, 876248.848757417, 
    908112.443257687, 939976.037757957, 971839.632258226, 1003703.2267585, 
    1035566.82125877, 1067430.41575904, 1099294.01025931, 1131157.60475958, 
    1163021.19925985, 1194884.79376012, 1226748.38826039, 1258611.98276065, 
    1290475.57726092, 1322339.17176119, 1354202.76626146, 1386066.36076173, 
    1417929.955262, 1449793.54976227, 1481657.14426254, 1513520.73876281, 
    1545384.33326308, 1577247.92776335, 1609111.52226362, 1640975.11676389, 
    1672838.71126416, 1704702.30576443, 1736565.9002647,
  15876.5669640253, 47629.7008920759, 79382.8348201278, 111135.968748181, 
    142889.102676233, 174642.236604285, 206395.370532338, 238148.50446039, 
    269901.638388442, 301654.772316495, 333407.906244547, 365161.040172599, 
    396914.174100652, 428667.308028704, 460420.441956756, 492173.575884809, 
    523926.709812861, 555679.843740913, 587432.977668965, 619186.111597019, 
    650939.245525071, 682692.379453123, 714445.513381176, 746198.647309228, 
    777951.78123728, 809704.915165333, 841458.049093385, 873211.183021437, 
    904964.31694949, 936717.450877543, 968470.584805595, 1000223.71873365, 
    1031976.8526617, 1063729.98658975, 1095483.1205178, 1127236.25444586, 
    1158989.38837391, 1190742.52230196, 1222495.65623001, 1254248.79015807, 
    1286001.92408612, 1317755.05801417, 1349508.19194222, 1381261.32587028, 
    1413014.45979833, 1444767.59372638, 1476520.72765443, 1508273.86158249, 
    1540026.99551054, 1571780.12943859, 1603533.26336664, 1635286.39729469, 
    1667039.53122275, 1698792.6651508, 1730545.79907885,
  15820.7993152066, 47462.3979456197, 79103.9965760342, 110745.59520645, 
    142387.193836865, 174028.792467279, 205670.391097695, 237311.989728109, 
    268953.588358524, 300595.18698894, 332236.785619354, 363878.384249769, 
    395519.982880185, 427161.581510599, 458803.180141014, 490444.77877143, 
    522086.377401844, 553727.976032258, 585369.574662673, 617011.173293089, 
    648652.771923504, 680294.370553919, 711935.969184334, 743577.567814749, 
    775219.166445163, 806860.765075579, 838502.363705994, 870143.962336408, 
    901785.560966823, 933427.159597239, 965068.758227653, 996710.356858068, 
    1028351.95548848, 1059993.5541189, 1091635.15274931, 1123276.75137973, 
    1154918.35001014, 1186559.94864056, 1218201.54727097, 1249843.14590139, 
    1281484.7445318, 1313126.34316222, 1344767.94179263, 1376409.54042305, 
    1408051.13905346, 1439692.73768388, 1471334.33631429, 1502975.93494471, 
    1534617.53357512, 1566259.13220554, 1597900.73083595, 1629542.32946637, 
    1661183.92809678, 1692825.5267272, 1724467.12535761,
  15764.4961912364, 47293.4885737092, 78822.4809561833, 110351.473338659, 
    141880.465721133, 173409.458103607, 204938.450486082, 236467.442868557, 
    267996.435251031, 299525.427633506, 331054.42001598, 362583.412398455, 
    394112.40478093, 425641.397163404, 457170.389545878, 488699.381928354, 
    520228.374310828, 551757.366693301, 583286.359075776, 614815.351458251, 
    646344.343840726, 677873.3362232, 709402.328605675, 740931.32098815, 
    772460.313370624, 803989.305753099, 835518.298135574, 867047.290518048, 
    898576.282900523, 930105.275282998, 961634.267665472, 993163.260047947, 
    1024692.25243042, 1056221.2448129, 1087750.23719537, 1119279.22957785, 
    1150808.22196032, 1182337.21434279, 1213866.20672527, 1245395.19910774, 
    1276924.19149022, 1308453.18387269, 1339982.17625517, 1371511.16863764, 
    1403040.16102012, 1434569.15340259, 1466098.14578507, 1497627.13816754, 
    1529156.13055002, 1560685.12293249, 1592214.11531496, 1623743.10769744, 
    1655272.10007991, 1686801.09246239, 1718330.08484486,
  15707.659497797, 47122.9784933911, 78538.2974889865, 109953.616484583, 
    141368.935480179, 172784.254475774, 204199.573471371, 235614.892466966, 
    267030.211462562, 298445.530458159, 329860.849453754, 361276.168449349, 
    392691.487444946, 424106.806440542, 455522.125436137, 486937.444431734, 
    518352.763427329, 549768.082422924, 581183.40141852, 612598.720414117, 
    644014.039409713, 675429.358405308, 706844.677400904, 738259.996396501, 
    769675.315392096, 801090.634387692, 832505.953383288, 863921.272378884, 
    895336.59137448, 926751.910370076, 958167.229365671, 989582.548361267, 
    1020997.86735686, 1052413.18635246, 1083828.50534805, 1115243.82434365, 
    1146659.14333925, 1178074.46233484, 1209489.78133044, 1240905.10032603, 
    1272320.41932163, 1303735.73831723, 1335151.05731282, 1366566.37630842, 
    1397981.69530401, 1429397.01429961, 1460812.33329521, 1492227.6522908, 
    1523642.9712864, 1555058.29028199, 1586473.60927759, 1617888.92827318, 
    1649304.24726878, 1680719.56626438, 1712134.88525997,
  15650.2911586302, 46950.8734758905, 78251.4557931521, 109552.038110415, 
    140852.620427677, 172153.202744938, 203453.785062201, 234754.367379463, 
    266054.949696725, 297355.532013988, 328656.114331249, 359956.696648511, 
    391257.278965774, 422557.861283036, 453858.443600297, 485159.02591756, 
    516459.608234822, 547760.190552083, 579060.772869345, 610361.355186608, 
    641661.937503871, 672962.519821132, 704263.102138394, 735563.684455657, 
    766864.266772918, 798164.849090181, 829465.431407443, 860766.013724705, 
    892066.596041967, 923367.178359229, 954667.760676491, 985968.342993753, 
    1017268.92531102, 1048569.50762828, 1079870.08994554, 1111170.6722628, 
    1142471.25458006, 1173771.83689733, 1205072.41921459, 1236373.00153185, 
    1267673.58384911, 1298974.16616637, 1330274.74848364, 1361575.3308009, 
    1392875.91311816, 1424176.49543542, 1455477.07775268, 1486777.66006995, 
    1518078.24238721, 1549378.82470447, 1580679.40702173, 1611979.98933899, 
    1643280.57165626, 1674581.15397352, 1705881.73629078,
  15592.3931154715, 46777.1793464145, 77961.9655773589, 109146.751808305, 
    140331.538039249, 171516.324270193, 202701.110501139, 233885.896732083, 
    265070.682963028, 296255.469193973, 327440.255424918, 358625.041655862, 
    389809.827886808, 420994.614117752, 452179.400348696, 483364.186579642, 
    514548.972810586, 545733.75904153, 576918.545272475, 608103.331503421, 
    639288.117734366, 670472.90396531, 701657.690196255, 732842.4764272, 
    764027.262658145, 795212.04888909, 826396.835120035, 857581.621350979, 
    888766.407581924, 919951.193812869, 951135.980043813, 982320.766274758, 
    1013505.5525057, 1044690.33873665, 1075875.12496759, 1107059.91119854, 
    1138244.69742948, 1169429.48366043, 1200614.26989137, 1231799.05612232, 
    1262983.84235326, 1294168.62858421, 1325353.41481515, 1356538.2010461, 
    1387722.98727704, 1418907.77350799, 1450092.55973893, 1481277.34596988, 
    1512462.13220082, 1543646.91843176, 1574831.70466271, 1606016.49089365, 
    1637201.2771246, 1668386.06335554, 1699570.84958649,
  15533.9673279853, 46601.901983956, 77669.836639928, 108737.771295901, 
    139805.705951873, 170873.640607845, 201941.575263819, 233009.509919791, 
    264077.444575763, 295145.379231736, 326213.313887708, 357281.24854368, 
    388349.183199653, 419417.117855625, 450485.052511597, 481552.987167571, 
    512620.921823543, 543688.856479514, 574756.791135487, 605824.72579146, 
    636892.660447433, 667960.595103405, 699028.529759378, 730096.46441535, 
    761164.399071322, 792232.333727295, 823300.268383268, 854368.20303924, 
    885436.137695213, 916504.072351185, 947572.007007157, 978639.94166313, 
    1009707.8763191, 1040775.81097507, 1071843.74563105, 1102911.68028702, 
    1133979.61494299, 1165047.54959896, 1196115.48425494, 1227183.41891091, 
    1258251.35356688, 1289319.28822285, 1320387.22287883, 1351455.1575348, 
    1382523.09219077, 1413591.02684674, 1444658.96150272, 1475726.89615869, 
    1506794.83081466, 1537862.76547063, 1568930.70012661, 1599998.63478258, 
    1631066.56943855, 1662134.50409452, 1693202.4387505,
  15475.015773698, 46425.047321094, 77375.0788684913, 108325.11041589, 
    139275.141963287, 170225.173510685, 201175.205058083, 232125.236605481, 
    263075.268152878, 294025.299700277, 324975.331247674, 355925.362795071, 
    386875.39434247, 417825.425889867, 448775.457437265, 479725.488984663, 
    510675.520532061, 541625.552079457, 572575.583626855, 603525.615174254, 
    634475.646721652, 665425.678269049, 696375.709816447, 727325.741363845, 
    758275.772911243, 789225.804458641, 820175.836006039, 851125.867553436, 
    882075.899100834, 913025.930648232, 943975.962195629, 974925.993743028, 
    1005876.02529043, 1036826.05683782, 1067776.08838522, 1098726.11993262, 
    1129676.15148002, 1160626.18302741, 1191576.21457481, 1222526.24612221, 
    1253476.27766961, 1284426.30921701, 1315376.3407644, 1346326.3723118, 
    1377276.4038592, 1408226.4354066, 1439176.46695399, 1470126.49850139, 
    1501076.53004879, 1532026.56159619, 1562976.59314358, 1593926.62469098, 
    1624876.65623838, 1655826.68778578, 1686776.71933318,
  15415.540447931, 46246.6213437931, 77077.7022396564, 107908.783135521, 
    138739.864031384, 169570.944927248, 200402.025823112, 231233.106718976, 
    262064.187614839, 292895.268510704, 323726.349406567, 354557.430302431, 
    385388.511198295, 416219.592094159, 447050.672990022, 477881.753885887, 
    508712.83478175, 539543.915677613, 570374.996573476, 601206.077469341, 
    632037.158365205, 662868.239261068, 693699.320156932, 724530.401052797, 
    755361.48194866, 786192.562844524, 817023.643740388, 847854.724636251, 
    878685.805532115, 909516.886427979, 940347.967323842, 971179.048219707, 
    1002010.12911557, 1032841.21001143, 1063672.2909073, 1094503.37180316, 
    1125334.45269903, 1156165.53359489, 1186996.61449075, 1217827.69538662, 
    1248658.77628248, 1279489.85717834, 1310320.93807421, 1341152.01897007, 
    1371983.09986594, 1402814.1807618, 1433645.26165766, 1464476.34255353, 
    1495307.42344939, 1526138.50434525, 1556969.58524112, 1587800.66613698, 
    1618631.74703284, 1649462.82792871, 1680293.90882457,
  15355.5433637335, 46066.6300912005, 76777.7168186689, 107488.803546139, 
    138199.890273607, 168910.977001075, 199622.063728545, 230333.150456013, 
    261044.237183481, 291755.323910951, 322466.410638419, 353177.497365888, 
    383888.584093357, 414599.670820826, 445310.757548294, 476021.844275764, 
    506732.931003232, 537444.0177307, 568155.104458169, 598866.191185638, 
    629577.277913107, 660288.364640576, 690999.451368045, 721710.538095514, 
    752421.624822982, 783132.711550451, 813843.79827792, 844554.885005388, 
    875265.971732857, 905977.058460326, 936688.145187795, 967399.231915264, 
    998110.318642733, 1028821.4053702, 1059532.49209767, 1090243.57882514, 
    1120954.66555261, 1151665.75228008, 1182376.83900755, 1213087.92573501, 
    1243799.01246248, 1274510.09918995, 1305221.18591742, 1335932.27264489, 
    1366643.35937236, 1397354.44609983, 1428065.53282729, 1458776.61955476, 
    1489487.70628223, 1520198.7930097, 1550909.87973717, 1581620.96646464, 
    1612332.05319211, 1643043.13991958, 1673754.22664704,
  15295.0265518141, 45885.0796554423, 76475.1327590719, 107065.185862703, 
    137655.238966332, 168245.292069962, 198835.345173593, 229425.398277222, 
    260015.451380852, 290605.504484482, 321195.557588112, 351785.610691742, 
    382375.663795372, 412965.716899002, 443555.770002631, 474145.823106262, 
    504735.876209892, 535325.929313521, 565915.982417151, 596506.035520782, 
    627096.088624412, 657686.141728041, 688276.194831672, 718866.247935302, 
    749456.301038931, 780046.354142562, 810636.407246192, 841226.460349821, 
    871816.513453451, 902406.566557082, 932996.619660711, 963586.672764341, 
    994176.725867972, 1024766.7789716, 1055356.83207523, 1085946.88517886, 
    1116536.93828249, 1147126.99138612, 1177717.04448975, 1208307.09759338, 
    1238897.15069701, 1269487.20380064, 1300077.25690427, 1330667.3100079, 
    1361257.36311153, 1391847.41621516, 1422437.46931879, 1453027.52242242, 
    1483617.57552605, 1514207.62862968, 1544797.68173331, 1575387.73483694, 
    1605977.78794057, 1636567.8410442, 1667157.89414783,
  15233.9920604722, 45701.9761814166, 76169.9603023622, 106637.944423309, 
    137105.928544255, 167573.912665201, 198041.896786147, 228509.880907093, 
    258977.865028039, 289445.849148986, 319913.833269931, 350381.817390877, 
    380849.801511824, 411317.78563277, 441785.769753715, 472253.753874662, 
    502721.737995608, 533189.722116553, 563657.706237499, 594125.690358446, 
    624593.674479393, 655061.658600338, 685529.642721285, 715997.626842231, 
    746465.610963177, 776933.595084123, 807401.579205069, 837869.563326015, 
    868337.547446961, 898805.531567908, 929273.515688853, 959741.4998098, 
    990209.483930746, 1020677.46805169, 1051145.45217264, 1081613.43629358, 
    1112081.42041453, 1142549.40453548, 1173017.38865642, 1203485.37277737, 
    1233953.35689831, 1264421.34101926, 1294889.32514021, 1325357.30926115, 
    1355825.2933821, 1386293.27750305, 1416761.26162399, 1447229.24574494, 
    1477697.22986588, 1508165.21398683, 1538633.19810778, 1569101.18222872, 
    1599569.16634967, 1630037.15047061, 1660505.13459156,
  15172.4419555285, 45517.3258665855, 75862.2097776438, 106207.093688703, 
    136551.977599762, 166896.86151082, 197241.745421879, 227586.629332938, 
    257931.513243996, 288276.397155056, 318621.281066114, 348966.164977172, 
    379311.048888232, 409655.93279929, 440000.816710348, 470345.700621408, 
    500690.584532466, 531035.468443524, 561380.352354583, 591725.236265642, 
    622070.120176701, 652415.00408776, 682759.887998819, 713104.771909878, 
    743449.655820936, 773794.539731995, 804139.423643054, 834484.307554112, 
    864829.191465171, 895174.07537623, 925518.959287288, 955863.843198347, 
    986208.727109406, 1016553.61102046, 1046898.49493152, 1077243.37884258, 
    1107588.26275364, 1137933.1466647, 1168278.03057576, 1198622.91448682, 
    1228967.79839788, 1259312.68230893, 1289657.56621999, 1320002.45013105, 
    1350347.33404211, 1380692.21795317, 1411037.10186423, 1441381.98577529, 
    1471726.86968634, 1502071.7535974, 1532416.63750846, 1562761.52141952, 
    1593106.40533058, 1623451.28924164, 1653796.1731527,
  15110.3783202553, 45331.1349607658, 75551.8916012777, 105772.648241791, 
    135993.404882303, 166214.161522815, 196434.918163328, 226655.674803839, 
    256876.431444351, 287097.188084865, 317317.944725376, 347538.701365888, 
    377759.458006401, 407980.214646913, 438200.971287425, 468421.727927938, 
    498642.48456845, 528863.241208961, 559083.997849474, 589304.754489987, 
    619525.511130499, 649746.267771011, 679967.024411524, 710187.781052036, 
    740408.537692548, 770629.29433306, 800850.050973573, 831070.807614085, 
    861291.564254597, 891512.32089511, 921733.077535621, 951953.834176134, 
    982174.590816646, 1012395.34745716, 1042616.10409767, 1072836.86073818, 
    1103057.61737869, 1133278.37401921, 1163499.13065972, 1193719.88730023, 
    1223940.64394074, 1254161.40058126, 1284382.15722177, 1314602.91386228, 
    1344823.67050279, 1375044.42714331, 1405265.18378382, 1435485.94042433, 
    1465706.69706484, 1495927.45370535, 1526148.21034587, 1556368.96698638, 
    1586589.72362689, 1616810.4802674, 1647031.23690792,
  15047.8032553057, 45143.4097659172, 75239.01627653, 105334.622787144, 
    135430.229297757, 165525.83580837, 195621.442318983, 225717.048829596, 
    255812.655340209, 285908.261850823, 316003.868361436, 346099.474872049, 
    376195.081382663, 406290.687893275, 436386.294403888, 466481.900914502, 
    496577.507425115, 526673.113935727, 556768.720446341, 586864.326956955, 
    616959.933467568, 647055.539978181, 677151.146488794, 707246.752999407, 
    737342.35951002, 767437.966020634, 797533.572531247, 827629.17904186, 
    857724.785552473, 887820.392063087, 917915.9985737, 948011.605084313, 
    978107.211594926, 1008202.81810554, 1038298.42461615, 1068394.03112677, 
    1098489.63763738, 1128585.24414799, 1158680.85065861, 1188776.45716922, 
    1218872.06367983, 1248967.67019044, 1279063.27670106, 1309158.88321167, 
    1339254.48972228, 1369350.0962329, 1399445.70274351, 1429541.30925412, 
    1459636.91576474, 1489732.52227535, 1519828.12878596, 1549923.73529657, 
    1580019.34180719, 1610114.9483178, 1640210.55482841,
  14984.7188786429, 44954.1566359287, 74923.5943932158, 104893.032150504, 
    134862.469907791, 164831.907665078, 194801.345422367, 224770.783179654, 
    254740.220936941, 284709.658694229, 314679.096451516, 344648.534208803, 
    374617.971966092, 404587.409723379, 434556.847480666, 464526.285237954, 
    494495.722995241, 524465.160752527, 554434.598509815, 584404.036267104, 
    614373.474024391, 644342.911781678, 674312.349538966, 704281.787296254, 
    734251.225053541, 764220.662810828, 794190.100568116, 824159.538325403, 
    854128.976082691, 884098.413839979, 914067.851597266, 944037.289354553, 
    974006.727111841, 1003976.16486913, 1033945.60262642, 1063915.0403837, 
    1093884.47814099, 1123853.91589828, 1153823.35365557, 1183792.79141285, 
    1213762.22917014, 1243731.66692743, 1273701.10468472, 1303670.542442, 
    1333639.98019929, 1363609.41795658, 1393578.85571387, 1423548.29347115, 
    1453517.73122844, 1483487.16898573, 1513456.60674302, 1543426.0445003, 
    1573395.48225759, 1603364.92001488, 1633334.35777217,
  14921.127325468, 44763.3819764039, 74605.6366273411, 104447.89127828, 
    134290.145929217, 164132.400580154, 193974.655231093, 223816.90988203, 
    253659.164532967, 283501.419183905, 313343.673834843, 343185.92848578, 
    373028.183136718, 402870.437787656, 432712.692438593, 462554.947089531, 
    492397.201740469, 522239.456391405, 552081.711042343, 581923.965693281, 
    611766.220344219, 641608.474995156, 671450.729646094, 701292.984297032, 
    731135.238947969, 760977.493598907, 790819.748249845, 820662.002900782, 
    850504.25755172, 880346.512202658, 910188.766853595, 940031.021504533, 
    969873.276155471, 999715.530806408, 1029557.78545735, 1059400.04010828, 
    1089242.29475922, 1119084.54941016, 1148926.8040611, 1178769.05871203, 
    1208611.31336297, 1238453.56801391, 1268295.82266485, 1298138.07731578, 
    1327980.33196672, 1357822.58661766, 1387664.8412686, 1417507.09591954, 
    1447349.35057047, 1477191.60522141, 1507033.85987235, 1536876.11452328, 
    1566718.36917422, 1596560.62382516, 1626402.8784761,
  14857.030748148, 44571.0922444441, 74285.1537407413, 103999.21523704, 
    133713.276733337, 163427.338229635, 193141.399725933, 222855.46122223, 
    252569.522718528, 282283.584214826, 311997.645711123, 341711.707207421, 
    371425.768703719, 401139.830200017, 430853.891696314, 460567.953192613, 
    490282.01468891, 519996.076185207, 549710.137681504, 579424.199177803, 
    609138.260674101, 638852.322170398, 668566.383666696, 698280.445162994, 
    727994.506659291, 757708.568155589, 787422.629651887, 817136.691148184, 
    846850.752644482, 876564.81414078, 906278.875637077, 935992.937133375, 
    965706.998629673, 995421.06012597, 1025135.12162227, 1054849.18311857, 
    1084563.24461486, 1114277.30611116, 1143991.36760746, 1173705.42910376, 
    1203419.49060005, 1233133.55209635, 1262847.61359265, 1292561.67508895, 
    1322275.73658525, 1351989.79808154, 1381703.85957784, 1411417.92107414, 
    1441131.98257044, 1470846.04406673, 1500560.10556303, 1530274.16705933, 
    1559988.22855563, 1589702.29005192, 1619416.35154822,
  14792.4313161431, 44377.2939484293, 73962.1565807168, 103547.019213006, 
    133131.881845293, 162716.744477581, 192301.607109869, 221886.469742157, 
    251471.332374444, 281056.195006733, 310641.05763902, 340225.920271308, 
    369810.782903597, 399395.645535884, 428980.508168172, 458565.37080046, 
    488150.233432748, 517735.096065035, 547319.958697323, 576904.821329612, 
    606489.6839619, 636074.546594187, 665659.409226475, 695244.271858763, 
    724829.134491051, 754413.997123339, 783998.859755627, 813583.722387914, 
    843168.585020202, 872753.44765249, 902338.310284778, 931923.172917066, 
    961508.035549354, 991092.898181641, 1020677.76081393, 1050262.62344622, 
    1079847.4860785, 1109432.34871079, 1139017.21134308, 1168602.07397537, 
    1198186.93660766, 1227771.79923995, 1257356.66187223, 1286941.52450452, 
    1316526.38713681, 1346111.2497691, 1375696.11240138, 1405280.97503367, 
    1434865.83766596, 1464450.70029825, 1494035.56293054, 1523620.42556282, 
    1553205.28819511, 1582790.1508274, 1612375.01345969,
  14727.3312159329, 44181.9936477988, 73636.6560796658, 103091.318511534, 
    132545.980943401, 162000.643375268, 191455.305807137, 220909.968239004, 
    250364.630670871, 279819.293102739, 309273.955534606, 338728.617966473, 
    368183.280398342, 397637.942830209, 427092.605262076, 456547.267693944, 
    486001.930125811, 515456.592557678, 544911.254989545, 574365.917421414, 
    603820.579853281, 633275.242285149, 662729.904717016, 692184.567148884, 
    721639.229580751, 751093.892012619, 780548.554444487, 810003.216876354, 
    839457.879308221, 868912.541740089, 898367.204171956, 927821.866603824, 
    957276.529035692, 986731.191467559, 1016185.85389943, 1045640.51633129, 
    1075095.17876316, 1104549.84119503, 1134004.5036269, 1163459.16605876, 
    1192913.82849063, 1222368.4909225, 1251823.15335437, 1281277.81578623, 
    1310732.4782181, 1340187.14064997, 1369641.80308184, 1399096.4655137, 
    1428551.12794557, 1458005.79037744, 1487460.45280931, 1516915.11524117, 
    1546369.77767304, 1575824.44010491, 1605279.10253678,
  14661.7326509427, 43985.197952828, 73308.6632547146, 102632.128556602, 
    131955.593858489, 161279.059160376, 190602.524462263, 219925.98976415, 
    249249.455066037, 278572.920367924, 307896.385669811, 337219.850971698, 
    366543.316273585, 395866.781575472, 425190.246877359, 454513.712179246, 
    483837.177481133, 513160.642783019, 542484.108084906, 571807.573386794, 
    601131.038688681, 630454.503990568, 659777.969292455, 689101.434594342, 
    718424.899896229, 747748.365198116, 777071.830500003, 806395.29580189, 
    835718.761103777, 865042.226405664, 894365.691707551, 923689.157009438, 
    953012.622311325, 982336.087613211, 1011659.5529151, 1040983.01821699, 
    1070306.48351887, 1099629.94882076, 1128953.41412265, 1158276.87942453, 
    1187600.34472642, 1216923.81002831, 1246247.27533019, 1275570.74063208, 
    1304894.20593397, 1334217.67123586, 1363541.13653774, 1392864.60183963, 
    1422188.06714152, 1451511.5324434, 1480834.99774529, 1510158.46304718, 
    1539481.92834906, 1568805.39365095, 1598128.85895284,
  14595.6378414686, 43786.9135244057, 72978.189207344, 102169.464890284, 
    131360.740573222, 160552.01625616, 189743.2919391, 218934.567622038, 
    248125.843304977, 277317.118987916, 306508.394670855, 335699.670353793, 
    364890.946036733, 394082.221719671, 423273.497402609, 452464.773085549, 
    481656.048768487, 510847.324451425, 540038.600134364, 569229.875817304, 
    598421.151500243, 627612.427183181, 656803.70286612, 685994.978549059, 
    715186.254231997, 744377.529914936, 773568.805597875, 802760.081280814, 
    831951.356963753, 861142.632646692, 890333.90832963, 919525.184012569, 
    948716.459695508, 977907.735378447, 1007099.01106139, 1036290.28674432, 
    1065481.56242726, 1094672.8381102, 1123864.11379314, 1153055.38947608, 
    1182246.66515902, 1211437.94084196, 1240629.2165249, 1269820.49220783, 
    1299011.76789077, 1328203.04357371, 1357394.31925665, 1386585.59493959, 
    1415776.87062253, 1444968.14630547, 1474159.42198841, 1503350.69767134, 
    1532541.97335428, 1561733.24903722, 1590924.52472016,
  14529.0490246026, 43587.1470738079, 72645.2451230143, 101703.343172222, 
    130761.441221429, 159819.539270635, 188877.637319843, 217935.735369049, 
    246993.833418256, 276051.931467463, 305110.02951667, 334168.127565876, 
    363226.225615084, 392284.323664291, 421342.421713497, 450400.519762705, 
    479458.617811911, 508516.715861117, 537574.813910324, 566632.911959532, 
    595691.010008739, 624749.108057946, 653807.206107153, 682865.30415636, 
    711923.402205566, 740981.500254773, 770039.59830398, 799097.696353187, 
    828155.794402394, 857213.892451601, 886271.990500807, 915330.088550014, 
    944388.186599221, 973446.284648428, 1002504.38269763, 1031562.48074684, 
    1060620.57879605, 1089678.67684526, 1118736.77489446, 1147794.87294367, 
    1176852.97099288, 1205911.06904208, 1234969.16709129, 1264027.2651405, 
    1293085.3631897, 1322143.46123891, 1351201.55928812, 1380259.65733732, 
    1409317.75538653, 1438375.85343574, 1467433.95148494, 1496492.04953415, 
    1525550.14758336, 1554608.24563257, 1583666.34368177,
  14461.968454157, 43385.9053624709, 72309.8422707861, 101233.779179103, 
    130157.716087418, 159081.652995733, 188005.589904049, 216929.526812364, 
    245853.46372068, 274777.400628996, 303701.337537311, 332625.274445626, 
    361549.211353943, 390473.148262258, 419397.085170573, 448321.02207889, 
    477244.958987205, 506168.895895519, 535092.832803835, 564016.769712151, 
    592940.706620467, 621864.643528783, 650788.580437098, 679712.517345414, 
    708636.454253729, 737560.391162045, 766484.328070361, 795408.264978676, 
    824332.201886992, 853256.138795308, 882180.075703623, 911104.012611939, 
    940027.949520255, 968951.88642857, 997875.823336886, 1026799.7602452, 
    1055723.69715352, 1084647.63406183, 1113571.57097015, 1142495.50787846, 
    1171419.44478678, 1200343.38169509, 1229267.31860341, 1258191.25551173, 
    1287115.19242004, 1316039.12932836, 1344963.06623667, 1373887.00314499, 
    1402810.9400533, 1431734.87696162, 1460658.81386993, 1489582.75077825, 
    1518506.68768657, 1547430.62459488, 1576354.5615032,
  14394.3984005876, 43183.1952017627, 71971.992002939, 100760.788804117, 
    129549.585605293, 158338.382406469, 187127.179207647, 215915.976008823, 
    244704.772809999, 273493.569611177, 302282.366412353, 331071.16321353, 
    359859.960014707, 388648.756815884, 417437.55361706, 446226.350418237, 
    475015.147219414, 503803.944020589, 532592.740821766, 561381.537622944, 
    590170.334424121, 618959.131225297, 647747.928026474, 676536.724827651, 
    705325.521628827, 734114.318430004, 762903.115231181, 791691.912032357, 
    820480.708833534, 849269.505634711, 878058.302435888, 906847.099237064, 
    935635.896038241, 964424.692839418, 993213.489640594, 1022002.28644177, 
    1050791.08324295, 1079579.88004412, 1108368.6768453, 1137157.47364648, 
    1165946.27044766, 1194735.06724883, 1223523.86405001, 1252312.66085119, 
    1281101.45765236, 1309890.25445354, 1338679.05125472, 1367467.84805589, 
    1396256.64485707, 1425045.44165825, 1453834.23845942, 1482623.0352606, 
    1511411.83206178, 1540200.62886295, 1568989.42566413,
  14326.3411509172, 42979.0234527517, 71631.7057545873, 100284.388056424, 
    128937.07035826, 157589.752660096, 186242.434961932, 214895.117263768, 
    243547.799565604, 272200.481867441, 300853.164169276, 329505.846471112, 
    358158.528772949, 386811.211074785, 415463.89337662, 444116.575678457, 
    472769.257980293, 501421.940282128, 530074.622583964, 558727.304885801, 
    587379.987187637, 616032.669489473, 644685.351791309, 673338.034093145, 
    701990.716394981, 730643.398696817, 759296.080998654, 787948.763300489, 
    816601.445602325, 845254.127904162, 873906.810205997, 902559.492507834, 
    931212.17480967, 959864.857111505, 988517.539413342, 1017170.22171518, 
    1045822.90401701, 1074475.58631885, 1103128.26862069, 1131780.95092252, 
    1160433.63322436, 1189086.31552619, 1217738.99782803, 1246391.68012987, 
    1275044.3624317, 1303697.04473354, 1332349.72703537, 1361002.40933721, 
    1389655.09163905, 1418307.77394088, 1446960.45624272, 1475613.13854455, 
    1504265.82084639, 1532918.50314823, 1561571.18545006,
  14257.7990086584, 42773.3970259752, 71288.9950432932, 99804.5930606124, 
    128320.19107793, 156835.789095248, 185351.387112568, 213866.985129886, 
    242382.583147204, 270898.181164523, 299413.779181841, 327929.377199159, 
    356444.975216478, 384960.573233796, 413476.171251114, 441991.769268433, 
    470507.367285751, 499022.965303069, 527538.563320387, 556054.161337706, 
    584569.759355025, 613085.357372343, 641600.955389661, 670116.55340698, 
    698632.151424298, 727147.749441617, 755663.347458935, 784178.945476253, 
    812694.543493572, 841210.14151089, 869725.739528208, 898241.337545527, 
    926756.935562845, 955272.533580163, 983788.131597482, 1012303.7296148, 
    1040819.32763212, 1069334.92564944, 1097850.52366676, 1126366.12168407, 
    1154881.71970139, 1183397.31771871, 1211912.91573603, 1240428.51375335, 
    1268944.11177067, 1297459.70978798, 1325975.3078053, 1354490.90582262, 
    1383006.50383994, 1411522.10185726, 1440037.69987458, 1468553.29789189, 
    1497068.89590921, 1525584.49392653, 1554100.09194385,
  14188.774293735, 42566.3228812051, 70943.8714686764, 99321.4200561489, 
    127698.96864362, 156076.517231091, 184454.065818564, 212831.614406035, 
    241209.162993507, 269586.711580979, 297964.26016845, 326341.808755922, 
    354719.357343394, 383096.905930865, 411474.454518337, 439852.003105809, 
    468229.55169328, 496607.100280751, 524984.648868223, 553362.197455695, 
    581739.746043167, 610117.294630639, 638494.843218111, 666872.391805582, 
    695249.940393054, 723627.488980525, 752005.037567997, 780382.586155469, 
    808760.134742941, 837137.683330412, 865515.231917884, 893892.780505355, 
    922270.329092827, 950647.877680299, 979025.426267771, 1007402.97485524, 
    1035780.52344271, 1064158.07203019, 1092535.62061766, 1120913.16920513, 
    1149290.7177926, 1177668.26638007, 1206045.81496754, 1234423.36355502, 
    1262800.91214249, 1291178.46072996, 1319556.00931743, 1347933.5579049, 
    1376311.10649237, 1404688.65507984, 1433066.20366732, 1461443.75225479, 
    1489821.30084226, 1518198.84942973, 1546576.3980172,
  14119.2693424041, 42357.8080272124, 70596.3467120219, 98834.8853968326, 
    127073.424081642, 155311.962766452, 183550.501451262, 211789.040136072, 
    240027.578820881, 268266.117505692, 296504.656190501, 324743.194875311, 
    352981.733560122, 381220.272244931, 409458.810929741, 437697.349614551, 
    465935.888299361, 494174.42698417, 522412.96566898, 550651.504353791, 
    578890.043038601, 607128.58172341, 635367.12040822, 663605.65909303, 
    691844.19777784, 720082.73646265, 748321.27514746, 776559.81383227, 
    804798.35251708, 833036.89120189, 861275.429886699, 889513.968571509, 
    917752.507256319, 945991.045941129, 974229.584625939, 1002468.12331075, 
    1030706.66199556, 1058945.20068037, 1087183.73936518, 1115422.27804999, 
    1143660.8167348, 1171899.35541961, 1200137.89410442, 1228376.43278923, 
    1256614.97147404, 1284853.51015885, 1313092.04884366, 1341330.58752847, 
    1369569.12621328, 1397807.66489809, 1426046.2035829, 1454284.74226771, 
    1482523.28095252, 1510761.81963733, 1539000.35832214,
  14049.2865071767, 42147.85952153, 70246.4325358846, 98345.0055502403, 
    126443.578564595, 154542.151578949, 182640.724593305, 210739.29760766, 
    238837.870622014, 266936.44363637, 295035.016650725, 323133.589665079, 
    351232.162679435, 379330.735693789, 407429.308708144, 435527.8817225, 
    463626.454736854, 491725.027751208, 519823.600765563, 547922.173779919, 
    576020.746794274, 604119.319808629, 632217.892822984, 660316.465837339, 
    688415.038851694, 716513.611866049, 744612.184880404, 772710.757894758, 
    800809.330909114, 828907.903923469, 857006.476937823, 885105.049952178, 
    913203.622966534, 941302.195980888, 969400.768995243, 997499.342009599, 
    1025597.91502395, 1053696.48803831, 1081795.06105266, 1109893.63406702, 
    1137992.20708137, 1166090.78009573, 1194189.35311008, 1222287.92612444, 
    1250386.49913879, 1278485.07215315, 1306583.6451675, 1334682.21818186, 
    1362780.79119621, 1390879.36421057, 1418977.93722492, 1447076.51023928, 
    1475175.08325363, 1503273.65626799, 1531372.22928234,
  13978.8281567379, 41936.4844702137, 69894.1407836906, 97851.7970971688, 
    125809.453410646, 153767.109724123, 181724.766037601, 209682.422351078, 
    237640.078664555, 265597.734978033, 293555.39129151, 321513.047604987, 
    349470.703918465, 377428.360231942, 405386.016545419, 433343.672858897, 
    461301.329172374, 489258.98548585, 517216.641799328, 545174.298112806, 
    573131.954426284, 601089.610739761, 629047.267053238, 657004.923366716, 
    684962.579680193, 712920.23599367, 740877.892307148, 768835.548620625, 
    796793.204934102, 824750.86124758, 852708.517561057, 880666.173874534, 
    908623.830188012, 936581.486501489, 964539.142814966, 992496.799128444, 
    1020454.45544192, 1048412.1117554, 1076369.76806888, 1104327.42438235, 
    1132285.08069583, 1160242.73700931, 1188200.39332278, 1216158.04963626, 
    1244115.70594974, 1272073.36226322, 1300031.01857669, 1327988.67489017, 
    1355946.33120365, 1383903.98751713, 1411861.6438306, 1439819.30014408, 
    1467776.95645756, 1495734.61277104, 1523692.26908451,
  13907.8966758672, 41723.6900276015, 69539.4833793371, 97355.2767310738, 
    125171.070082809, 152986.863434545, 180802.656786282, 208618.450138017, 
    236434.243489753, 264250.036841489, 292065.830193225, 319881.623544961, 
    347697.416896697, 375513.210248433, 403329.003600168, 431144.796951905, 
    458960.590303641, 486776.383655376, 514592.177007112, 542407.970358848, 
    570223.763710584, 598039.55706232, 625855.350414056, 653671.143765792, 
    681486.937117528, 709302.730469264, 737118.523821, 764934.317172736, 
    792750.110524472, 820565.903876208, 848381.697227944, 876197.49057968, 
    904013.283931416, 931829.077283152, 959644.870634888, 987460.663986624, 
    1015276.45733836, 1043092.2506901, 1070908.04404183, 1098723.83739357, 
    1126539.6307453, 1154355.42409704, 1182171.21744877, 1209987.01080051, 
    1237802.80415225, 1265618.59750398, 1293434.39085572, 1321250.18420745, 
    1349065.97755919, 1376881.77091093, 1404697.56426266, 1432513.3576144, 
    1460329.15096613, 1488144.94431787, 1515960.7376696,
  13836.4944653574, 41509.4833960721, 69182.472326788, 96855.4612575051, 
    124528.450188221, 152201.439118937, 179874.428049654, 207547.41698037, 
    235220.405911086, 262893.394841803, 290566.383772519, 318239.372703235, 
    345912.361633952, 373585.350564668, 401258.339495384, 428931.328426101, 
    456604.317356817, 484277.306287532, 511950.295218249, 539623.284148966, 
    567296.273079682, 594969.262010398, 622642.250941115, 650315.239871831, 
    677988.228802547, 705661.217733264, 733334.20666398, 761007.195594696, 
    788680.184525413, 816353.173456129, 844026.162386845, 871699.151317562, 
    899372.140248278, 927045.129178994, 954718.118109711, 982391.107040427, 
    1010064.09597114, 1037737.08490186, 1065410.07383258, 1093083.06276329, 
    1120756.05169401, 1148429.04062473, 1176102.02955544, 1203775.01848616, 
    1231448.00741687, 1259120.99634759, 1286793.98527831, 1314466.97420902, 
    1342139.96313974, 1369812.95207046, 1397485.94100117, 1425158.92993189, 
    1452831.9188626, 1480504.90779332, 1508177.89672404,
  13764.6239419334, 41293.8718258003, 68823.1197096683, 96352.3675935375, 
    123881.615477406, 151410.863361274, 178940.111245143, 206469.359129011, 
    233998.607012879, 261527.854896748, 289057.102780616, 316586.350664484, 
    344115.598548353, 371644.846432221, 399174.094316089, 426703.342199959, 
    454232.590083827, 481761.837967694, 509291.085851563, 536820.333735432, 
    564349.5816193, 591878.829503169, 619408.077387037, 646937.325270906, 
    674466.573154774, 701995.821038642, 729525.068922511, 757054.316806379, 
    784583.564690248, 812112.812574117, 839642.060457984, 867171.308341853, 
    894700.556225722, 922229.80410959, 949759.051993459, 977288.299877327, 
    1004817.5477612, 1032346.79564506, 1059876.04352893, 1087405.2914128, 
    1114934.53929667, 1142463.78718054, 1169993.03506441, 1197522.28294827, 
    1225051.53083214, 1252580.77871601, 1280110.02659988, 1307639.27448375, 
    1335168.52236762, 1362697.77025148, 1390227.01813535, 1417756.26601922, 
    1445285.51390309, 1472814.76178696, 1500344.00967082,
  13692.2875381707, 41076.862614512, 68461.4376908544, 95846.0127671981, 
    123230.587843541, 150615.162919883, 177999.737996227, 205384.313072569, 
    232768.888148912, 260153.463225255, 287538.038301598, 314922.61337794, 
    342307.188454284, 369691.763530626, 397076.338606969, 424460.913683312, 
    451845.488759655, 479230.063835997, 506614.63891234, 533999.213988683, 
    561383.789065026, 588768.364141369, 616152.939217712, 643537.514294055, 
    670922.089370397, 698306.66444674, 725691.239523083, 753075.814599426, 
    780460.389675769, 807844.964752112, 835229.539828454, 862614.114904797, 
    889998.68998114, 917383.265057483, 944767.840133826, 972152.415210169, 
    999536.990286511, 1026921.56536285, 1054306.1404392, 1081690.71551554, 
    1109075.29059188, 1136459.86566823, 1163844.44074457, 1191229.01582091, 
    1218613.59089726, 1245998.1659736, 1273382.74104994, 1300767.31612628, 
    1328151.89120263, 1355536.46627897, 1382921.04135531, 1410305.61643165, 
    1437690.191508, 1465074.76658434, 1492459.34166068,
  13619.4877024124, 40858.4631072371, 68097.4385120629, 95336.41391689, 
    122575.389321716, 149814.364726542, 177053.340131369, 204292.315536195, 
    231531.290941021, 258770.266345848, 286009.241750673, 313248.217155499, 
    340487.192560326, 367726.167965152, 394965.143369978, 422204.118774805, 
    449443.094179631, 476682.069584456, 503921.044989283, 531160.02039411, 
    558398.995798936, 585637.971203762, 612876.946608589, 640115.922013415, 
    667354.897418241, 694593.872823067, 721832.848227894, 749071.82363272, 
    776310.799037546, 803549.774442373, 830788.749847198, 858027.725252025, 
    885266.700656851, 912505.676061677, 939744.651466504, 966983.62687133, 
    994222.602276156, 1021461.57768098, 1048700.55308581, 1075939.52849063, 
    1103178.50389546, 1130417.47930029, 1157656.45470511, 1184895.43010994, 
    1212134.40551477, 1239373.38091959, 1266612.35632442, 1293851.33172924, 
    1321090.30713407, 1348329.2825389, 1375568.25794372, 1402807.23334855, 
    1430046.20875337, 1457285.1841582, 1484524.15956303,
  13546.226898687, 40638.6806960609, 67731.134493436, 94823.5882908123, 
    121916.042088187, 149008.495885563, 176100.949682939, 203193.403480314, 
    230285.857277689, 257378.311075065, 284470.76487244, 311563.218669816, 
    338655.672467192, 365748.126264567, 392840.580061942, 419933.033859318, 
    447025.487656693, 474117.941454068, 501210.395251444, 528302.84904882, 
    555395.302846196, 582487.756643571, 609580.210440946, 636672.664238322, 
    663765.118035697, 690857.571833073, 717950.025630448, 745042.479427823, 
    772134.933225199, 799227.387022575, 826319.84081995, 853412.294617326, 
    880504.748414701, 907597.202212076, 934689.656009452, 961782.109806828, 
    988874.563604203, 1015967.01740158, 1043059.47119895, 1070151.92499633, 
    1097244.3787937, 1124336.83259108, 1151429.28638846, 1178521.74018583, 
    1205614.19398321, 1232706.64778058, 1259799.10157796, 1286891.55537533, 
    1313984.00917271, 1341076.46297008, 1368168.91676746, 1395261.37056483, 
    1422353.82436221, 1449446.27815959, 1476538.73195696,
  13472.5076066247, 40417.522819874, 67362.5380331245, 94307.5532463762, 
    121252.568459627, 148197.583672877, 175142.598886129, 202087.614099379, 
    229032.62931263, 255977.644525881, 282922.659739132, 309867.674952382, 
    336812.690165634, 363757.705378885, 390702.720592135, 417647.735805387, 
    444592.751018637, 471537.766231887, 498482.781445138, 525427.79665839, 
    552372.811871641, 579317.827084891, 606262.842298143, 633207.857511394, 
    660152.872724644, 687097.887937895, 714042.903151146, 740987.918364397, 
    767932.933577648, 794877.948790899, 821822.96400415, 848767.979217401, 
    875712.994430652, 902658.009643903, 929603.024857154, 956548.040070405, 
    983493.055283655, 1010438.07049691, 1037383.08571016, 1064328.10092341, 
    1091273.11613666, 1118218.13134991, 1145163.14656316, 1172108.16177641, 
    1199053.17698966, 1225998.19220291, 1252943.20741616, 1279888.22262941, 
    1306833.23784267, 1333778.25305592, 1360723.26826917, 1387668.28348242, 
    1414613.29869567, 1441558.31390892, 1468503.32912217,
  13398.3323213734, 40194.9969641202, 66991.6616068681, 93788.3262496171, 
    120584.990892365, 147381.655535113, 174178.320177862, 200974.98482061, 
    227771.649463358, 254568.314106107, 281364.978748855, 308161.643391603, 
    334958.308034352, 361754.9726771, 388551.637319848, 415348.301962597, 
    442144.966605345, 468941.631248092, 495738.29589084, 522534.96053359, 
    549331.625176338, 576128.289819086, 602924.954461834, 629721.619104583, 
    656518.283747331, 683314.948390079, 710111.613032828, 736908.277675576, 
    763704.942318324, 790501.606961073, 817298.271603821, 844094.936246569, 
    870891.600889318, 897688.265532066, 924484.930174814, 951281.594817563, 
    978078.259460311, 1004874.92410306, 1031671.58874581, 1058468.25338856, 
    1085264.9180313, 1112061.58267405, 1138858.2473168, 1165654.91195955, 
    1192451.5766023, 1219248.24124505, 1246044.90588779, 1272841.57053054, 
    1299638.23517329, 1326434.89981604, 1353231.56445879, 1380028.22910154, 
    1406824.89374428, 1433621.55838703, 1460418.22302978,
  13323.7035535144, 39971.1106605432, 66618.5177675731, 93265.9248746042, 
    119913.331981634, 146560.739088664, 173208.146195695, 199855.553302725, 
    226502.960409755, 253150.367516786, 279797.774623816, 306445.181730846, 
    333092.588837877, 359739.995944907, 386387.403051937, 413034.810158968, 
    439682.217265998, 466329.624373027, 492977.031480058, 519624.438587089, 
    546271.845694119, 572919.252801149, 599566.65990818, 626214.06701521, 
    652861.47412224, 679508.881229271, 706156.288336301, 732803.695443331, 
    759451.102550362, 786098.509657392, 812745.916764422, 839393.323871453, 
    866040.730978483, 892688.138085513, 919335.545192543, 945982.952299574, 
    972630.359406604, 999277.766513634, 1025925.17362066, 1052572.58072769, 
    1079219.98783473, 1105867.39494176, 1132514.80204879, 1159162.20915582, 
    1185809.61626285, 1212457.02336988, 1239104.43047691, 1265751.83758394, 
    1292399.24469097, 1319046.651798, 1345694.05890503, 1372341.46601206, 
    1398988.87311909, 1425636.28022612, 1452283.68733315,
  13248.6238289773, 39745.8714869319, 66243.1191448877, 92740.3668028446, 
    119237.6144608, 145734.862118756, 172232.109776713, 198729.357434669, 
    225226.605092625, 251723.852750581, 278221.100408537, 304718.348066493, 
    331215.59572445, 357712.843382406, 384210.091040361, 410707.338698318, 
    437204.586356274, 463701.834014229, 490199.081672186, 516696.329330143, 
    543193.576988099, 569690.824646055, 596188.072304011, 622685.319961967, 
    649182.567619923, 675679.815277879, 702177.062935836, 728674.310593791, 
    755171.558251748, 781668.805909704, 808166.05356766, 834663.301225616, 
    861160.548883572, 887657.796541528, 914155.044199484, 940652.291857441, 
    967149.539515397, 993646.787173353, 1020144.03483131, 1046641.28248926, 
    1073138.53014722, 1099635.77780518, 1126133.02546313, 1152630.27312109, 
    1179127.52077905, 1205624.768437, 1232122.01609496, 1258619.26375291, 
    1285116.51141087, 1311613.75906883, 1338111.00672678, 1364608.25438474, 
    1391105.50204269, 1417602.74970065, 1444099.99735861,
  13173.0956889546, 39519.2870668638, 65865.4784447742, 92211.6698226857, 
    118557.861200596, 144904.052578506, 171250.243956418, 197596.435334328, 
    223942.626712239, 250288.81809015, 276635.00946806, 302981.200845971, 
    329327.392223882, 355673.583601793, 382019.774979703, 408365.966357614, 
    434712.157735525, 461058.349113435, 487404.540491346, 513750.731869257, 
    540096.923247168, 566443.114625078, 592789.306002989, 619135.4973809, 
    645481.68875881, 671827.880136721, 698174.071514632, 724520.262892543, 
    750866.454270453, 777212.645648364, 803558.837026275, 829905.028404186, 
    856251.219782096, 882597.411160007, 908943.602537918, 935289.793915829, 
    961635.985293739, 987982.17667165, 1014328.36804956, 1040674.55942747, 
    1067020.75080538, 1093366.94218329, 1119713.1335612, 1146059.32493911, 
    1172405.51631703, 1198751.70769494, 1225097.89907285, 1251444.09045076, 
    1277790.28182867, 1304136.47320658, 1330482.66458449, 1356828.8559624, 
    1383175.04734031, 1409521.23871822, 1435867.43009613,
  13097.1216898156, 39291.3650694468, 65485.6084490792, 91679.8518287126, 
    117874.095208345, 144068.338587977, 170262.581967611, 196456.825347243, 
    222651.068726875, 248845.312106509, 275039.555486141, 301233.798865774, 
    327428.042245407, 353622.285625039, 379816.529004672, 406010.772384305, 
    432205.015763938, 458399.259143569, 484593.502523202, 510787.745902836, 
    536981.989282469, 563176.232662101, 589370.476041734, 615564.719421367, 
    641758.962800999, 667953.206180632, 694147.449560265, 720341.692939897, 
    746535.93631953, 772730.179699163, 798924.423078795, 825118.666458428, 
    851312.909838061, 877507.153217694, 903701.396597326, 929895.639976959, 
    956089.883356592, 982284.126736225, 1008478.37011586, 1034672.61349549, 
    1060866.85687512, 1087061.10025476, 1113255.34363439, 1139449.58701402, 
    1165643.83039365, 1191838.07377329, 1218032.31715292, 1244226.56053255, 
    1270420.80391218, 1296615.04729182, 1322809.29067145, 1349003.53405108, 
    1375197.77743071, 1401392.02081035, 1427586.26418998,
  13020.7044030199, 39062.1132090597, 65103.5220151006, 91144.9308211426, 
    117186.339627183, 143227.748433224, 169269.157239266, 195310.566045307, 
    221351.974851348, 247393.38365739, 273434.792463431, 299476.201269472, 
    325517.610075514, 351559.018881555, 377600.427687596, 403641.836493638, 
    429683.245299679, 455724.654105719, 481766.06291176, 507807.471717802, 
    533848.880523844, 559890.289329885, 585931.698135926, 611973.106941968, 
    638014.515748008, 664055.92455405, 690097.333360091, 716138.742166132, 
    742180.150972174, 768221.559778215, 794262.968584256, 820304.377390297, 
    846345.786196339, 872387.19500238, 898428.603808421, 924470.012614463, 
    950511.421420504, 976552.830226545, 1002594.23903259, 1028635.64783863, 
    1054677.05664467, 1080718.46545071, 1106759.87425675, 1132801.28306279, 
    1158842.69186883, 1184884.10067488, 1210925.50948092, 1236966.91828696, 
    1263008.327093, 1289049.73589904, 1315091.14470508, 1341132.55351112, 
    1367173.96231716, 1393215.3711232, 1419256.77992925,
  12943.8464150303, 38831.539245091, 64719.2320751527, 90606.9249052156, 
    116494.617735277, 142382.310565339, 168270.003395402, 194157.696225464, 
    220045.389055525, 245933.081885588, 271820.77471565, 297708.467545712, 
    323596.160375775, 349483.853205836, 375371.546035898, 401259.238865961, 
    427146.931696023, 453034.624526084, 478922.317356146, 504810.010186209, 
    530697.703016271, 556585.395846333, 582473.088676395, 608360.781506457, 
    634248.474336519, 660136.167166581, 686023.859996644, 711911.552826706, 
    737799.245656768, 763686.93848683, 789574.631316892, 815462.324146954, 
    841350.016977016, 867237.709807078, 893125.402637141, 919013.095467203, 
    944900.788297265, 970788.481127327, 996676.173957389, 1022563.86678745, 
    1048451.55961751, 1074339.25244758, 1100226.94527764, 1126114.6381077, 
    1152002.33093776, 1177890.02376782, 1203777.71659789, 1229665.40942795, 
    1255553.10225801, 1281440.79508807, 1307328.48791813, 1333216.1807482, 
    1359103.87357826, 1384991.56640832, 1410879.25923838,
  12866.5503272255, 38599.6509816764, 64332.7516361284, 90065.8522905816, 
    115798.952945034, 141532.053599486, 167265.154253939, 192998.254908391, 
    218731.355562843, 244464.456217296, 270197.556871748, 295930.6575262, 
    321663.758180653, 347396.858835105, 373129.959489557, 398863.06014401, 
    424596.160798462, 450329.261452914, 476062.362107367, 501795.46276182, 
    527528.563416272, 553261.664070724, 578994.764725177, 604727.865379629, 
    630460.966034082, 656194.066688534, 681927.167342987, 707660.267997439, 
    733393.368651891, 759126.469306344, 784859.569960796, 810592.670615248, 
    836325.771269701, 862058.871924153, 887791.972578605, 913525.073233058, 
    939258.17388751, 964991.274541963, 990724.375196415, 1016457.47585087, 
    1042190.57650532, 1067923.67715977, 1093656.77781422, 1119389.87846868, 
    1145122.97912313, 1170856.07977758, 1196589.18043203, 1222322.28108649, 
    1248055.38174094, 1273788.48239539, 1299521.58304984, 1325254.6837043, 
    1350987.78435875, 1376720.8850132, 1402453.98566765,
  12788.8187558116, 38366.4562674347, 63944.0937790589, 89521.7312906842, 
    115099.368802308, 140677.006313933, 166254.643825558, 191832.281337182, 
    217409.918848806, 242987.556360432, 268565.193872056, 294142.83138368, 
    319720.468895305, 345298.10640693, 370875.743918554, 396453.381430179, 
    422031.018941803, 447608.656453427, 473186.293965052, 498763.931476677, 
    524341.568988302, 549919.206499926, 575496.844011551, 601074.481523175, 
    626652.1190348, 652229.756546424, 677807.394058049, 703385.031569674, 
    728962.669081298, 754540.306592923, 780117.944104547, 805695.581616172, 
    831273.219127797, 856850.856639421, 882428.494151046, 908006.131662671, 
    933583.769174295, 959161.40668592, 984739.044197545, 1010316.68170917, 
    1035894.31922079, 1061471.95673242, 1087049.59424404, 1112627.23175567, 
    1138204.86926729, 1163782.50677892, 1189360.14429054, 1214937.78180217, 
    1240515.41931379, 1266093.05682542, 1291670.69433704, 1317248.33184866, 
    1342825.96936029, 1368403.60687191, 1393981.24438354,
  12710.6543317339, 38131.9629952018, 63553.2716586707, 88974.5803221407, 
    114395.88898561, 139817.197649079, 165238.506312549, 190659.814976018, 
    216081.123639486, 241502.432302956, 266923.740966425, 292345.049629894, 
    317766.358293364, 343187.666956833, 368608.975620302, 394030.284283772, 
    419451.592947241, 444872.90161071, 470294.210274179, 495715.518937649, 
    521136.827601119, 546558.136264588, 571979.444928057, 597400.753591527, 
    622822.062254995, 648243.370918465, 673664.679581934, 699085.988245403, 
    724507.296908873, 749928.605572342, 775349.914235811, 800771.22289928, 
    826192.53156275, 851613.840226219, 877035.148889688, 902456.457553158, 
    927877.766216627, 953299.074880096, 978720.383543566, 1004141.69220703, 
    1029563.0008705, 1054984.30953397, 1080405.61819744, 1105826.92686091, 
    1131248.23552438, 1156669.54418785, 1182090.85285132, 1207512.16151479, 
    1232933.47017826, 1258354.77884173, 1283776.0875052, 1309197.39616867, 
    1334618.70483214, 1360040.0134956, 1385461.32215907,
  12632.0597005879, 37896.1791017638, 63160.2985029408, 88424.4179041188, 
    113688.537305296, 138952.656706473, 164216.776107651, 189480.895508828, 
    214745.014910005, 240009.134311183, 265273.25371236, 290537.373113537, 
    315801.492514715, 341065.611915892, 366329.731317069, 391593.850718247, 
    416857.970119424, 442122.0895206, 467386.208921778, 492650.328322956, 
    517914.447724133, 543178.56712531, 568442.686526487, 593706.805927665, 
    618970.925328842, 644235.044730019, 669499.164131197, 694763.283532374, 
    720027.402933551, 745291.522334729, 770555.641735906, 795819.761137083, 
    821083.880538261, 846347.999939438, 871612.119340615, 896876.238741793, 
    922140.35814297, 947404.477544147, 972668.596945325, 997932.716346502, 
    1023196.83574768, 1048460.95514886, 1073725.07455003, 1098989.19395121, 
    1124253.31335239, 1149517.43275357, 1174781.55215474, 1200045.67155592, 
    1225309.7909571, 1250573.91035827, 1275838.02975945, 1301102.14916063, 
    1326366.26856181, 1351630.38796298, 1376894.50736416,
  12553.0375225295, 37659.1125675885, 62765.1876126486, 87871.2626577097, 
    112977.33770277, 138083.41274783, 163189.487792891, 188295.562837951, 
    213401.637883011, 238507.712928072, 263613.787973132, 288719.863018192, 
    313825.938063253, 338932.013108313, 364038.088153374, 389144.163198435, 
    414250.238243495, 439356.313288554, 464462.388333615, 489568.463378676, 
    514674.538423737, 539780.613468796, 564886.688513857, 589992.763558918, 
    615098.838603978, 640204.913649038, 665310.988694099, 690417.063739159, 
    715523.13878422, 740629.21382928, 765735.28887434, 790841.363919401, 
    815947.438964461, 841053.514009521, 866159.589054582, 891265.664099643, 
    916371.739144703, 941477.814189763, 966583.889234824, 991689.964279884, 
    1016796.03932494, 1041902.11437001, 1067008.18941507, 1092114.26446013, 
    1117220.33950519, 1142326.41455025, 1167432.48959531, 1192538.56464037, 
    1217644.63968543, 1242750.71473049, 1267856.78977555, 1292962.86482061, 
    1318068.93986567, 1343175.01491073, 1368281.08995579,
  12473.5904721849, 37420.7714165547, 62367.9523609256, 87315.1333052975, 
    112262.314249668, 137209.495194039, 162156.676138411, 187103.857082782, 
    212051.038027153, 236998.218971525, 261945.399915896, 286892.580860267, 
    311839.761804639, 336786.94274901, 361734.12369338, 386681.304637752, 
    411628.485582123, 436575.666526494, 461522.847470865, 486470.028415237, 
    511417.209359608, 536364.390303979, 561311.571248351, 586258.752192722, 
    611205.933137093, 636153.114081464, 661100.295025836, 686047.475970207, 
    710994.656914578, 735941.83785895, 760889.018803321, 785836.199747692, 
    810783.380692064, 835730.561636434, 860677.742580806, 885624.923525177, 
    910572.104469548, 935519.28541392, 960466.466358291, 985413.647302662, 
    1010360.82824703, 1035308.00919141, 1060255.19013578, 1085202.37108015, 
    1110149.55202452, 1135096.73296889, 1160043.91391326, 1184991.09485763, 
    1209938.275802, 1234885.45674637, 1259832.63769075, 1284779.81863512, 
    1309726.99957949, 1334674.18052386, 1359621.36146823,
  12393.7212385604, 37181.1637156813, 61968.6061928033, 86756.0486699263, 
    111543.491147048, 136330.93362417, 161118.376101293, 185905.818578415, 
    210693.261055537, 235480.70353266, 260268.146009782, 285055.588486904, 
    309843.030964027, 334630.473441149, 359417.915918271, 384205.358395394, 
    408992.800872516, 433780.243349637, 458567.68582676, 483355.128303883, 
    508142.570781005, 532930.013258127, 557717.455735249, 582504.898212372, 
    607292.340689494, 632079.783166616, 656867.225643739, 681654.668120861, 
    706442.110597983, 731229.553075106, 756016.995552228, 780804.43802935, 
    805591.880506473, 830379.322983595, 855166.765460717, 879954.20793784, 
    904741.650414962, 929529.092892084, 954316.535369206, 979103.977846328, 
    1003891.42032345, 1028678.86280057, 1053466.3052777, 1078253.74775482, 
    1103041.19023194, 1127828.63270906, 1152616.07518618, 1177403.51766331, 
    1202190.96014043, 1226978.40261755, 1251765.84509467, 1276553.2875718, 
    1301340.73004892, 1326128.17252604, 1350915.61500316 ;

 x_v =
  0, 32027.1265791512, 64054.2531583023, 96081.3797374562, 128108.50631661, 
    160135.632895761, 192162.759474915, 224189.886054069, 256217.01263322, 
    288244.139212374, 320271.265791528, 352298.392370679, 384325.518949833, 
    416352.645528987, 448379.772108138, 480406.898687292, 512434.025266446, 
    544461.151845597, 576488.27842475, 608515.405003903, 640542.531583057, 
    672569.65816221, 704596.784741362, 736623.911320516, 768651.037899669, 
    800678.164478821, 832705.291057975, 864732.417637128, 896759.54421628, 
    928786.670795434, 960813.797374587, 992840.923953739, 1024868.05053289, 
    1056895.17711205, 1088922.3036912, 1120949.43027035, 1152976.5568495, 
    1185003.68342866, 1217030.81000781, 1249057.93658696, 1281085.06316612, 
    1313112.18974527, 1345139.31632442, 1377166.44290358, 1409193.56948273, 
    1441220.69606188, 1473247.82264103, 1505274.94922019, 1537302.07579934, 
    1569329.20237849, 1601356.32895765, 1633383.4555368, 1665410.58211595, 
    1697437.70869511, 1729464.83527426, 1761491.96185341,
  0, 31918.2855542959, 63836.5711085918, 95754.8566628905, 127673.142217189, 
    159591.427771485, 191509.713325784, 223427.998880082, 255346.284434378, 
    287264.569988677, 319182.855542976, 351101.141097272, 383019.42665157, 
    414937.712205869, 446855.997760165, 478774.283314463, 510692.568868762, 
    542610.854423058, 574529.139977355, 606447.425531654, 638365.711085953, 
    670283.99664025, 702202.282194547, 734120.567748846, 766038.853303143, 
    797957.138857441, 829875.424411739, 861793.709966036, 893711.995520334, 
    925630.281074632, 957548.56662893, 989466.852183227, 1021385.13773753, 
    1053303.42329182, 1085221.70884612, 1117139.99440042, 1149058.27995472, 
    1180976.56550901, 1212894.85106331, 1244813.13661761, 1276731.42217191, 
    1308649.70772621, 1340567.9932805, 1372486.2788348, 1404404.5643891, 
    1436322.8499434, 1468241.13549769, 1500159.42105199, 1532077.70660629, 
    1563995.99216059, 1595914.27771488, 1627832.56326918, 1659750.84882348, 
    1691669.13437778, 1723587.41993207, 1755505.70548637,
  0, 31808.3642141593, 63616.7284283186, 95425.0926424806, 127233.456856643, 
    159041.821070802, 190850.185284964, 222658.549499126, 254466.913713285, 
    286275.277927447, 318083.642141609, 349892.006355768, 381700.37056993, 
    413508.734784092, 445317.098998252, 477125.463212414, 508933.827426576, 
    540742.191640735, 572550.555854896, 604358.920069058, 636167.28428322, 
    667975.64849738, 699784.012711541, 731592.376925703, 763400.741139864, 
    795209.105354024, 827017.469568186, 858825.833782347, 890634.197996508, 
    922442.56221067, 954250.92642483, 986059.290638991, 1017867.65485315, 
    1049676.01906731, 1081484.38328147, 1113292.74749564, 1145101.1117098, 
    1176909.47592396, 1208717.84013812, 1240526.20435228, 1272334.56856644, 
    1304142.9327806, 1335951.29699476, 1367759.66120892, 1399568.02542309, 
    1431376.38963725, 1463184.75385141, 1494993.11806557, 1526801.48227973, 
    1558609.84649389, 1590418.21070805, 1622226.57492221, 1654034.93913637, 
    1685843.30335053, 1717651.6675647, 1749460.03177886,
  0, 31697.3662792319, 63394.7325584637, 95092.0988376983, 126789.465116933, 
    158486.831396165, 190184.197675399, 221881.563954634, 253578.930233866, 
    285276.2965131, 316973.662792335, 348671.029071567, 380368.395350801, 
    412065.761630036, 443763.127909268, 475460.494188502, 507157.860467737, 
    538855.226746969, 570552.593026202, 602249.959305436, 633947.325584671, 
    665644.691863904, 697342.058143137, 729039.424422372, 760736.790701605, 
    792434.156980838, 824131.523260073, 855828.889539306, 887526.255818539, 
    919223.622097774, 950920.988377007, 982618.35465624, 1014315.72093547, 
    1046013.08721471, 1077710.45349394, 1109407.81977318, 1141105.18605241, 
    1172802.55233164, 1204499.91861088, 1236197.28489011, 1267894.65116934, 
    1299592.01744858, 1331289.38372781, 1362986.75000704, 1394684.11628628, 
    1426381.48256551, 1458078.84884475, 1489776.21512398, 1521473.58140321, 
    1553170.94768245, 1584868.31396168, 1616565.68024091, 1648263.04652015, 
    1679960.41279938, 1711657.77907861, 1743355.14535785,
  0, 31585.295506443, 63170.5910128859, 94755.8865193316, 126341.182025777, 
    157926.47753222, 189511.773038666, 221097.068545112, 252682.364051555, 
    284267.659558, 315852.955064446, 347438.250570889, 379023.546077334, 
    410608.84158378, 442194.137090223, 473779.432596669, 505364.728103114, 
    536950.023609557, 568535.319116002, 600120.614622447, 631705.910128893, 
    663291.205635337, 694876.501141782, 726461.796648227, 758047.092154672, 
    789632.387661116, 821217.683167562, 852802.978674006, 884388.27418045, 
    915973.569686896, 947558.86519334, 979144.160699785, 1010729.45620623, 
    1042314.75171267, 1073900.04721912, 1105485.34272556, 1137070.63823201, 
    1168655.93373845, 1200241.2292449, 1231826.52475134, 1263411.82025779, 
    1294997.11576423, 1326582.41127068, 1358167.70677712, 1389753.00228357, 
    1421338.29779001, 1452923.59329646, 1484508.8888029, 1516094.18430935, 
    1547679.47981579, 1579264.77532224, 1610850.07082868, 1642435.36633513, 
    1674020.66184157, 1705605.95734801, 1737191.25285446,
  0, 31472.1556890334, 62944.3113780669, 94416.467067103, 125888.622756139, 
    157360.778445173, 188832.934134209, 220305.089823245, 251777.245512278, 
    283249.401201314, 314721.55689035, 346193.712579384, 377665.86826842, 
    409138.023957456, 440610.17964649, 472082.335335526, 503554.491024562, 
    535026.646713595, 566498.80240263, 597970.958091666, 629443.113780702, 
    660915.269469737, 692387.425158772, 723859.580847808, 755331.736536843, 
    786803.892225878, 818276.047914914, 849748.203603948, 881220.359292983, 
    912692.514982019, 944164.670671054, 975636.826360089, 1007108.98204913, 
    1038581.13773816, 1070053.29342719, 1101525.44911623, 1132997.60480527, 
    1164469.7604943, 1195941.91618334, 1227414.07187237, 1258886.22756141, 
    1290358.38325044, 1321830.53893948, 1353302.69462851, 1384774.85031755, 
    1416247.00600658, 1447719.16169562, 1479191.31738465, 1510663.47307369, 
    1542135.62876272, 1573607.78445176, 1605079.94014079, 1636552.09582983, 
    1668024.25151886, 1699496.4072079, 1730968.56289693,
  0, 31357.9506564272, 62715.9013128544, 94073.8519692843, 125431.802625714, 
    156789.753282141, 188147.703938571, 219505.654595001, 250863.605251428, 
    282221.555907858, 313579.506564288, 344937.457220715, 376295.407877145, 
    407653.358533575, 439011.309190002, 470369.259846432, 501727.210502862, 
    533085.161159289, 564443.111815718, 595801.062472148, 627159.013128577, 
    658516.963785006, 689874.914441435, 721232.865097864, 752590.815754293, 
    783948.766410721, 815306.717067151, 846664.66772358, 878022.618380008, 
    909380.569036438, 940738.519692867, 972096.470349295, 1003454.42100573, 
    1034812.37166215, 1066170.32231858, 1097528.27297501, 1128886.22363144, 
    1160244.17428787, 1191602.1249443, 1222960.07560073, 1254318.02625716, 
    1285675.97691359, 1317033.92757001, 1348391.87822644, 1379749.82888287, 
    1411107.7795393, 1442465.73019573, 1473823.68085216, 1505181.63150859, 
    1536539.58216502, 1567897.53282145, 1599255.48347788, 1630613.4341343, 
    1661971.38479073, 1693329.33544716, 1724687.28610359,
  0, 31242.6842741017, 62485.3685482033, 93728.0528223077, 124970.737096412, 
    156213.421370514, 187456.105644618, 218698.789918722, 249941.474192824, 
    281184.158466928, 312426.842741033, 343669.527015134, 374912.211289239, 
    406154.895563343, 437397.579837445, 468640.264111549, 499882.948385653, 
    531125.632659755, 562368.316933858, 593611.001207962, 624853.685482067, 
    656096.36975617, 687339.054030273, 718581.738304377, 749824.42257848, 
    781067.106852583, 812309.791126687, 843552.47540079, 874795.159674893, 
    906037.843948998, 937280.528223101, 968523.212497204, 999765.896771308, 
    1031008.58104541, 1062251.26531951, 1093493.94959362, 1124736.63386772, 
    1155979.31814182, 1187222.00241593, 1218464.68669003, 1249707.37096413, 
    1280950.05523824, 1312192.73951234, 1343435.42378645, 1374678.10806055, 
    1405920.79233465, 1437163.47660876, 1468406.16088286, 1499648.84515696, 
    1530891.52943107, 1562134.21370517, 1593376.89797927, 1624619.58225338, 
    1655862.26652748, 1687104.95080158, 1718347.63507569,
  0, 31126.3604434569, 62252.7208869137, 93379.0813303732, 124505.441773833, 
    155631.80221729, 186758.162660749, 217884.523104209, 249010.883547665, 
    280137.243991125, 311263.604434585, 342389.964878041, 373516.325321501, 
    404642.68576496, 435769.046208417, 466895.406651877, 498021.767095336, 
    529148.127538793, 560274.487982251, 591400.848425711, 622527.20886917, 
    653653.569312628, 684779.929756087, 715906.290199546, 747032.650643004, 
    778159.011086463, 809285.371529922, 840411.73197338, 871538.092416839, 
    902664.452860298, 933790.813303756, 964917.173747214, 996043.534190674, 
    1027169.89463413, 1058296.25507759, 1089422.61552105, 1120548.97596451, 
    1151675.33640797, 1182801.69685143, 1213928.05729488, 1245054.41773834, 
    1276180.7781818, 1307307.13862526, 1338433.49906872, 1369559.85951218, 
    1400686.21995564, 1431812.58039909, 1462938.94084255, 1494065.30128601, 
    1525191.66172947, 1556318.02217293, 1587444.38261639, 1618570.74305985, 
    1649697.1035033, 1680823.46394676, 1711949.82439022,
  0, 31008.9831016833, 62017.9662033667, 93026.9493050527, 124035.932406739, 
    155044.915508422, 186053.898610108, 217062.881711794, 248071.864813477, 
    279080.847915163, 310089.831016849, 341098.814118533, 372107.797220219, 
    403116.780321905, 434125.763423588, 465134.746525274, 496143.72962696, 
    527152.712728643, 558161.695830328, 589170.678932014, 620179.6620337, 
    651188.645135385, 682197.628237069, 713206.611338755, 744215.59444044, 
    775224.577542125, 806233.560643811, 837242.543745496, 868251.52684718, 
    899260.509948866, 930269.493050551, 961278.476152236, 992287.459253922, 
    1023296.44235561, 1054305.42545729, 1085314.40855898, 1116323.39166066, 
    1147332.37476235, 1178341.35786403, 1209350.34096572, 1240359.3240674, 
    1271368.30716909, 1302377.29027077, 1333386.27337246, 1364395.25647414, 
    1395404.23957583, 1426413.22267751, 1457422.2057792, 1488431.18888088, 
    1519440.17198257, 1550449.15508425, 1581458.13818594, 1612467.12128762, 
    1643476.10438931, 1674485.08749099, 1705494.07059268,
  0, 30890.556221629, 61781.112443258, 92671.6686648897, 123562.224886521, 
    154452.78110815, 185343.337329782, 216233.893551414, 247124.449773043, 
    278015.005994674, 308905.562216306, 339796.118437935, 370686.674659567, 
    401577.230881198, 432467.787102827, 463358.343324459, 494248.899546091, 
    525139.45576772, 556030.01198935, 586920.568210982, 617811.124432613, 
    648701.680654244, 679592.236875874, 710482.793097506, 741373.349319136, 
    772263.905540766, 803154.461762398, 834045.017984028, 864935.574205659, 
    895826.13042729, 926716.686648921, 957607.242870551, 988497.799092183, 
    1019388.35531381, 1050278.91153544, 1081169.46775708, 1112060.02397871, 
    1142950.58020034, 1173841.13642197, 1204731.6926436, 1235622.24886523, 
    1266512.80508686, 1297403.36130849, 1328293.91753012, 1359184.47375175, 
    1390075.02997338, 1420965.58619501, 1451856.14241664, 1482746.69863827, 
    1513637.2548599, 1544527.81108154, 1575418.36730317, 1606308.9235248, 
    1637199.47974643, 1668090.03596806, 1698980.59218969,
  0, 30771.0838116645, 61542.1676233291, 92313.2514349962, 123084.335246663, 
    153855.419058328, 184626.502869995, 215397.586681662, 246168.670493327, 
    276939.754304994, 307710.838116661, 338481.921928326, 369253.005739993, 
    400024.08955166, 430795.173363324, 461566.257174992, 492337.340986659, 
    523108.424798323, 553879.508609989, 584650.592421656, 615421.676233323, 
    646192.760044989, 676963.843856655, 707734.927668322, 738506.011479988, 
    769277.095291654, 800048.179103321, 830819.262914987, 861590.346726653, 
    892361.43053832, 923132.514349986, 953903.598161652, 984674.681973319, 
    1015445.76578498, 1046216.84959665, 1076987.93340832, 1107759.01721998, 
    1138530.10103165, 1169301.18484332, 1200072.26865498, 1230843.35246665, 
    1261614.43627831, 1292385.52008998, 1323156.60390165, 1353927.68771331, 
    1384698.77152498, 1415469.85533665, 1446240.93914831, 1477012.02295998, 
    1507783.10677164, 1538554.19058331, 1569325.27439498, 1600096.35820664, 
    1630867.44201831, 1661638.52582997, 1692409.60964164,
  0, 30650.5699155476, 61301.1398310952, 91951.7097466455, 122602.279662196, 
    153252.849577743, 183903.419493294, 214553.989408844, 245204.559324391, 
    275855.129239942, 306505.699155492, 337156.26907104, 367806.83898659, 
    398457.40890214, 429107.978817688, 459758.548733238, 490409.118648788, 
    521059.688564336, 551710.258479885, 582360.828395435, 613011.398310985, 
    643661.968226534, 674312.538142083, 704963.108057633, 735613.677973182, 
    766264.247888731, 796914.817804281, 827565.38771983, 858215.957635379, 
    888866.527550929, 919517.097466478, 950167.667382027, 980818.237297578, 
    1011468.80721313, 1042119.37712868, 1072769.94704423, 1103420.51695977, 
    1134071.08687532, 1164721.65679087, 1195372.22670642, 1226022.79662197, 
    1256673.36653752, 1287323.93645307, 1317974.50636862, 1348625.07628417, 
    1379275.64619972, 1409926.21611527, 1440576.78603082, 1471227.35594637, 
    1501877.92586192, 1532528.49577747, 1563179.06569301, 1593829.63560856, 
    1624480.20552411, 1655130.77543966, 1685781.34535521,
  0, 30529.0186122863, 61058.0372245726, 91587.0558368615, 122116.07444915, 
    152645.093061437, 183174.111673726, 213703.130286014, 244232.148898301, 
    274761.16751059, 305290.186122879, 335819.204735165, 366348.223347454, 
    396877.241959743, 427406.260572029, 457935.279184318, 488464.297796607, 
    518993.316408893, 549522.335021181, 580051.35363347, 610580.372245759, 
    641109.390858046, 671638.409470334, 702167.428082623, 732696.44669491, 
    763225.465307198, 793754.483919487, 824283.502531774, 854812.521144062, 
    885341.539756351, 915870.558368638, 946399.576980926, 976928.595593215, 
    1007457.6142055, 1037986.63281779, 1068515.65143008, 1099044.67004237, 
    1129573.68865465, 1160102.70726694, 1190631.72587923, 1221160.74449152, 
    1251689.76310381, 1282218.7817161, 1312747.80032838, 1343276.81894067, 
    1373805.83755296, 1404334.85616525, 1434863.87477754, 1465392.89338982, 
    1495921.91200211, 1526450.9306144, 1556979.94922669, 1587508.96783898, 
    1618037.98645126, 1648567.00506355, 1679096.02367584,
  0, 30406.4340160007, 60812.8680320014, 91219.3020480046, 121625.736064008, 
    152032.170080009, 182438.604096012, 212845.038112015, 243251.472128016, 
    273657.906144019, 304064.340160022, 334470.774176023, 364877.208192026, 
    395283.64220803, 425690.07622403, 456096.510240034, 486502.944256037, 
    516909.378272037, 547315.812288039, 577722.246304043, 608128.680320046, 
    638535.114336048, 668941.54835205, 699347.982368053, 729754.416384055, 
    760160.850400057, 790567.284416061, 820973.718432063, 851380.152448065, 
    881786.586464068, 912193.02048007, 942599.454496072, 973005.888512075, 
    1003412.32252808, 1033818.75654408, 1064225.19056008, 1094631.62457608, 
    1125038.05859209, 1155444.49260809, 1185850.92662409, 1216257.36064009, 
    1246663.7946561, 1277070.2286721, 1307476.6626881, 1337883.0967041, 
    1368289.53072011, 1398695.96473611, 1429102.39875211, 1459508.83276811, 
    1489915.26678412, 1520321.70080012, 1550728.13481612, 1581134.56883212, 
    1611541.00284813, 1641947.43686413, 1672353.87088013,
  0, 30282.8202757838, 60565.6405515675, 90848.4608273539, 121131.28110314, 
    151414.101378924, 181696.92165471, 211979.741930497, 242262.562206281, 
    272545.382482067, 302828.202757853, 333111.023033637, 363393.843309423, 
    393676.66358521, 423959.483860994, 454242.30413678, 484525.124412566, 
    514807.94468835, 545090.764964135, 575373.585239921, 605656.405515708, 
    635939.225791493, 666222.046067278, 696504.866343064, 726787.686618849, 
    757070.506894634, 787353.327170421, 817636.147446206, 847918.967721991, 
    878201.787997777, 908484.608273562, 938767.428549347, 969050.248825134, 
    999333.069100919, 1029615.8893767, 1059898.70965249, 1090181.52992828, 
    1120464.35020406, 1150747.17047985, 1181029.99075563, 1211312.81103142, 
    1241595.6313072, 1271878.45158299, 1302161.27185877, 1332444.09213456, 
    1362726.91241034, 1393009.73268613, 1423292.55296192, 1453575.3732377, 
    1483858.19351349, 1514141.01378927, 1544423.83406506, 1574706.65434084, 
    1604989.47461663, 1635272.29489241, 1665555.1151682,
  0, 30158.181575561, 60316.363151122, 90474.5447266856, 120632.726302249, 
    150790.90787781, 180949.089453374, 211107.271028937, 241265.452604498, 
    271423.634180062, 301581.815755626, 331739.997331187, 361898.17890675, 
    392056.360482314, 422214.542057875, 452372.723633438, 482530.905209002, 
    512689.086784563, 542847.268360125, 573005.449935689, 603163.631511252, 
    633321.813086815, 663479.994662377, 693638.176237941, 723796.357813503, 
    753954.539389065, 784112.720964629, 814270.902540191, 844429.084115753, 
    874587.265691317, 904745.447266879, 934903.628842442, 965061.810418005, 
    995219.991993567, 1025378.17356913, 1055536.35514469, 1085694.53672026, 
    1115852.71829582, 1146010.89987138, 1176169.08144694, 1206327.26302251, 
    1236485.44459807, 1266643.62617363, 1296801.80774919, 1326959.98932476, 
    1357118.17090032, 1387276.35247588, 1417434.53405145, 1447592.71562701, 
    1477750.89720257, 1507909.07877813, 1538067.2603537, 1568225.44192926, 
    1598383.62350482, 1628541.80508038, 1658699.98665595,
  0, 30032.5221339486, 60065.0442678973, 90097.5664018485, 120130.0885358, 
    150162.610669748, 180195.132803699, 210227.654937651, 240260.177071599, 
    270292.69920555, 300325.221339502, 330357.74347345, 360390.265607401, 
    390422.787741353, 420455.309875301, 450487.832009253, 480520.354143204, 
    510552.876277152, 540585.398411102, 570617.920545053, 600650.442679005, 
    630682.964812955, 660715.486946904, 690748.009080856, 720780.531214806, 
    750813.053348755, 780845.575482707, 810878.097616657, 840910.619750606, 
    870943.141884558, 900975.664018508, 931008.186152457, 961040.708286409, 
    991073.230420359, 1021105.75255431, 1051138.27468826, 1081170.79682221, 
    1111203.31895616, 1141235.84109011, 1171268.36322406, 1201300.88535801, 
    1231333.40749196, 1261365.92962591, 1291398.45175986, 1321430.97389381, 
    1351463.49602776, 1381496.01816171, 1411528.54029566, 1441561.06242961, 
    1471593.58456356, 1501626.10669751, 1531658.62883146, 1561691.15096541, 
    1591723.67309937, 1621756.19523331, 1651788.71736726,
  0, 29905.8462041109, 59811.6924082217, 89717.5386123352, 119623.384816449, 
    149529.231020559, 179435.077224673, 209340.923428786, 239246.769632897, 
    269152.615837011, 299058.462041124, 328964.308245235, 358870.154449348, 
    388776.000653462, 418681.846857573, 448587.693061686, 478493.539265799, 
    508399.38546991, 538305.231674022, 568211.077878136, 598116.924082249, 
    628022.770286361, 657928.616490473, 687834.462694587, 717740.308898699, 
    747646.155102811, 777552.001306925, 807457.847511037, 837363.693715149, 
    867269.539919262, 897175.386123374, 927081.232327486, 956987.0785316, 
    986892.924735712, 1016798.77093982, 1046704.61714394, 1076610.46334805, 
    1106516.30955216, 1136422.15575628, 1166328.00196039, 1196233.8481645, 
    1226139.69436861, 1256045.54057273, 1285951.38677684, 1315857.23298095, 
    1345763.07918506, 1375668.92538918, 1405574.77159329, 1435480.6177974, 
    1465386.46400151, 1495292.31020563, 1525198.15640974, 1555104.00261385, 
    1585009.84881796, 1614915.69502208, 1644821.54122619,
  0, 29778.158073616, 59556.316147232, 89334.4742208505, 119112.632294469, 
    148890.790368085, 178668.948441704, 208447.106515322, 238225.264588938, 
    268003.422662557, 297781.580736175, 327559.738809791, 357337.89688341, 
    387116.054957028, 416894.213030644, 446672.371104263, 476450.529177881, 
    506228.687251497, 536006.845325114, 565785.003398733, 595563.161472352, 
    625341.319545969, 655119.477619586, 684897.635693204, 714675.793766822, 
    744453.951840439, 774232.109914057, 804010.267987675, 833788.426061292, 
    863566.58413491, 893344.742208528, 923122.900282145, 952901.058355763, 
    982679.21642938, 1012457.374503, 1042235.53257662, 1072013.69065023, 
    1101791.84872385, 1131570.00679747, 1161348.16487109, 1191126.3229447, 
    1220904.48101832, 1250682.63909194, 1280460.79716556, 1310238.95523918, 
    1340017.11331279, 1369795.27138641, 1399573.42946003, 1429351.58753365, 
    1459129.74560726, 1488907.90368088, 1518686.0617545, 1548464.21982812, 
    1578242.37790173, 1608020.53597535, 1637798.69404897,
  0, 29649.4620642911, 59298.9241285822, 88948.3861928759, 118597.84825717, 
    148247.310321461, 177896.772385754, 207546.234450048, 237195.696514339, 
    266845.158578633, 296494.620642926, 326144.082707218, 355793.544771511, 
    385443.006835805, 415092.468900096, 444741.93096439, 474391.393028683, 
    504040.855092974, 533690.317157267, 563339.779221561, 592989.241285854, 
    622638.703350147, 652288.165414439, 681937.627478732, 711587.089543025, 
    741236.551607317, 770886.013671611, 800535.475735903, 830184.937800195, 
    859834.399864489, 889483.861928781, 919133.323993074, 948782.786057367, 
    978432.24812166, 1008081.71018595, 1037731.17225025, 1067380.63431454, 
    1097030.09637883, 1126679.55844312, 1156329.02050742, 1185978.48257171, 
    1215627.944636, 1245277.40670029, 1274926.86876459, 1304576.33082888, 
    1334225.79289317, 1363875.25495747, 1393524.71702176, 1423174.17908605, 
    1452823.64115034, 1482473.10321464, 1512122.56527893, 1541772.02734322, 
    1571421.48940752, 1601070.95147181, 1630720.4135361,
  0, 29519.762532076, 59039.5250641521, 88559.2875962306, 118079.050128309, 
    147598.812660385, 177118.575192464, 206638.337724542, 236158.100256618, 
    265677.862788697, 295197.625320775, 324717.387852851, 354237.15038493, 
    383756.912917009, 413276.675449084, 442796.437981163, 472316.200513242, 
    501835.963045318, 531355.725577395, 560875.488109473, 590395.250641552, 
    619915.013173629, 649434.775705707, 678954.538237785, 708474.300769862, 
    737994.06330194, 767513.825834018, 797033.588366095, 826553.350898173, 
    856073.113430251, 885592.875962328, 915112.638494406, 944632.401026484, 
    974152.163558562, 1003671.92609064, 1033191.68862272, 1062711.45115479, 
    1092231.21368687, 1121750.97621895, 1151270.73875103, 1180790.5012831, 
    1210310.26381518, 1239830.02634726, 1269349.78887934, 1298869.55141142, 
    1328389.31394349, 1357909.07647557, 1387428.83900765, 1416948.60153973, 
    1446468.3640718, 1475988.12660388, 1505507.88913596, 1535027.65166804, 
    1564547.41420012, 1594067.17673219, 1623586.93926427,
  0, 29389.0638668756, 58778.1277337512, 88167.1916006292, 117556.255467507, 
    146945.319334383, 176334.383201261, 205723.447068139, 235112.510935015, 
    264501.574801893, 293890.638668771, 323279.702535646, 352668.766402524, 
    382057.830269403, 411446.894136278, 440835.958003156, 470225.021870034, 
    499614.08573691, 529003.149603787, 558392.213470665, 587781.277337543, 
    617170.34120442, 646559.405071296, 675948.468938175, 705337.532805051, 
    734726.596671928, 764115.660538806, 793504.724405683, 822893.78827256, 
    852282.852139438, 881671.916006315, 911060.979873192, 940450.04374007, 
    969839.107606947, 999228.171473823, 1028617.2353407, 1058006.29920758, 
    1087395.36307446, 1116784.42694133, 1146173.49080821, 1175562.55467509, 
    1204951.61854197, 1234340.68240884, 1263729.74627572, 1293118.8101426, 
    1322507.87400947, 1351896.93787635, 1381286.00174323, 1410675.06561011, 
    1440064.12947698, 1469453.19334386, 1498842.25721074, 1528231.32107761, 
    1557620.38494449, 1587009.44881137, 1616398.51267825,
  0, 29257.3704924112, 58514.7409848224, 87772.1114772361, 117029.48196965, 
    146286.852462061, 175544.222954475, 204801.593446888, 234058.9639393, 
    263316.334431713, 292573.704924127, 321831.075416538, 351088.445908952, 
    380345.816401366, 409603.186893777, 438860.557386191, 468117.927878605, 
    497375.298371016, 526632.668863428, 555890.039355842, 585147.409848256, 
    614404.780340668, 643662.150833081, 672919.521325494, 702176.891817907, 
    731434.262310319, 760691.632802733, 789949.003295145, 819206.373787558, 
    848463.744279972, 877721.114772384, 906978.485264797, 936235.85575721, 
    965493.226249623, 994750.596742035, 1024007.96723445, 1053265.33772686, 
    1082522.70821927, 1111780.07871169, 1141037.4492041, 1170294.81969651, 
    1199552.19018893, 1228809.56068134, 1258066.93117375, 1287324.30166617, 
    1316581.67215858, 1345839.04265099, 1375096.4131434, 1404353.78363582, 
    1433611.15412823, 1462868.52462064, 1492125.89511305, 1521383.26560547, 
    1550640.63609788, 1579898.00659029, 1609155.37708271,
  0, 29124.6868660712, 58249.3737321424, 87374.060598216, 116498.74746429, 
    145623.434330361, 174748.121196435, 203872.808062508, 232997.494928579, 
    262122.181794653, 291246.868660727, 320371.555526798, 349496.242392872, 
    378620.929258945, 407745.616125016, 436870.30299109, 465994.989857164, 
    495119.676723235, 524244.363589307, 553369.050455381, 582493.737321455, 
    611618.424187527, 640743.1110536, 669867.797919673, 698992.484785746, 
    728117.171651818, 757241.858517891, 786366.545383964, 815491.232250036, 
    844615.91911611, 873740.605982182, 902865.292848255, 931989.979714328, 
    961114.666580401, 990239.353446473, 1019364.04031255, 1048488.72717862, 
    1077613.41404469, 1106738.10091077, 1135862.78777684, 1164987.47464291, 
    1194112.16150898, 1223236.84837506, 1252361.53524113, 1281486.2221072, 
    1310610.90897327, 1339735.59583935, 1368860.28270542, 1397984.96957149, 
    1427109.65643757, 1456234.34330364, 1485359.03016971, 1514483.71703578, 
    1543608.40390186, 1572733.09076793, 1601857.777634,
  0, 28991.0174787596, 57982.0349575192, 86973.0524362813, 115964.069915043, 
    144955.087393803, 173946.104872565, 202937.122351327, 231928.139830087, 
    260919.157308849, 289910.174787611, 318901.19226637, 347892.209745132, 
    376883.227223895, 405874.244702654, 434865.262181416, 463856.279660178, 
    492847.297138938, 521838.314617699, 550829.332096461, 579820.349575223, 
    608811.367053984, 637802.384532744, 666793.402011506, 695784.419490267, 
    724775.436969028, 753766.45444779, 782757.471926551, 811748.489405312, 
    840739.506884074, 869730.524362835, 898721.541841595, 927712.559320358, 
    956703.576799118, 985694.594277879, 1014685.61175664, 1043676.6292354, 
    1072667.64671416, 1101658.66419292, 1130649.68167169, 1159640.69915045, 
    1188631.71662921, 1217622.73410797, 1246613.75158673, 1275604.76906549, 
    1304595.78654425, 1333586.80402301, 1362577.82150178, 1391568.83898054, 
    1420559.8564593, 1449550.87393806, 1478541.89141682, 1507532.90889558, 
    1536523.92637434, 1565514.9438531, 1594505.96133186,
  0, 28856.3668547445, 57712.7337094891, 86569.100564236, 115425.467418983, 
    144281.834273728, 173138.201128475, 201994.567983222, 230850.934837966, 
    259707.301692713, 288563.66854746, 317420.035402205, 346276.402256952, 
    375132.769111698, 403989.135966443, 432845.50282119, 461701.869675937, 
    490558.236530681, 519414.603385427, 548270.970240174, 577127.337094921, 
    605983.703949667, 634840.070804413, 663696.43765916, 692552.804513905, 
    721409.171368651, 750265.538223398, 779121.905078144, 807978.27193289, 
    836834.638787637, 865691.005642382, 894547.372497128, 923403.739351875, 
    952260.106206621, 981116.473061366, 1009972.83991611, 1038829.20677086, 
    1067685.57362561, 1096541.94048035, 1125398.3073351, 1154254.67418984, 
    1183111.04104459, 1211967.40789934, 1240823.77475408, 1269680.14160883, 
    1298536.50846357, 1327392.87531832, 1356249.24217307, 1385105.60902781, 
    1413961.97588256, 1442818.34273731, 1471674.70959205, 1500531.0764468, 
    1529387.44330154, 1558243.81015629, 1587100.17701104,
  0, 28720.7395515048, 57441.4791030095, 86162.2186545168, 114882.958206024, 
    143603.697757529, 172324.437309036, 201045.176860543, 229765.916412048, 
    258486.655963555, 287207.395515062, 315928.135066567, 344648.874618074, 
    373369.614169582, 402090.353721086, 430811.093272594, 459531.832824101, 
    488252.572375606, 516973.311927112, 545694.051478619, 574414.791030126, 
    603135.530581632, 631856.270133138, 660577.009684645, 689297.749236151, 
    718018.488787657, 746739.228339164, 775459.96789067, 804180.707442176, 
    832901.446993683, 861622.186545189, 890342.926096695, 919063.665648203, 
    947784.405199709, 976505.144751214, 1005225.88430272, 1033946.62385423, 
    1062667.36340573, 1091388.10295724, 1120108.84250875, 1148829.58206025, 
    1177550.32161176, 1206271.06116327, 1234991.80071477, 1263712.54026628, 
    1292433.27981779, 1321154.01936929, 1349874.7589208, 1378595.4984723, 
    1407316.23802381, 1436036.97757532, 1464757.71712682, 1493478.45667833, 
    1522199.19622984, 1550919.93578134, 1579640.67533285,
  0, 28584.1401595756, 57168.2803191512, 85752.4204787293, 114336.560638307, 
    142920.700797883, 171504.840957461, 200088.981117039, 228673.121276615, 
    257257.261436193, 285841.401595771, 314425.541755346, 343009.681914924, 
    371593.822074502, 400177.962234078, 428762.102393656, 457346.242553234, 
    485930.38271281, 514514.522872387, 543098.663031965, 571682.803191543, 
    600266.94335112, 628851.083510696, 657435.223670274, 686019.363829851, 
    714603.503989428, 743187.644149006, 771771.784308583, 800355.92446816, 
    828940.064627738, 857524.204787314, 886108.344946891, 914692.485106469, 
    943276.625266046, 971860.765425623, 1000444.9055852, 1029029.04574478, 
    1057613.18590435, 1086197.32606393, 1114781.46622351, 1143365.60638309, 
    1171949.74654266, 1200533.88670224, 1229118.02686182, 1257702.1670214, 
    1286286.30718097, 1314870.44734055, 1343454.58750013, 1372038.7276597, 
    1400622.86781928, 1429207.00797886, 1457791.14813843, 1486375.28829801, 
    1514959.42845759, 1543543.56861717, 1572127.70877674,
  0, 28446.5733023934, 56893.1466047868, 85339.7199071827, 113786.293209579, 
    142232.866511972, 170679.439814368, 199126.013116764, 227572.586419157, 
    256019.159721553, 284465.733023949, 312912.306326342, 341358.879628738, 
    369805.452931134, 398252.026233527, 426698.599535923, 455145.172838319, 
    483591.746140713, 512038.319443107, 540484.892745503, 568931.466047899, 
    597378.039350293, 625824.612652688, 654271.185955084, 682717.759257479, 
    711164.332559873, 739610.905862269, 768057.479164664, 796504.052467058, 
    824950.625769454, 853397.199071849, 881843.772374243, 910290.345676639, 
    938736.918979034, 967183.492281428, 995630.065583824, 1024076.63888622, 
    1052523.21218861, 1080969.78549101, 1109416.3587934, 1137862.9320958, 
    1166309.50539819, 1194756.07870059, 1223202.65200298, 1251649.22530538, 
    1280095.79860777, 1308542.37191017, 1336988.94521256, 1365435.51851496, 
    1393882.09181735, 1422328.66511975, 1450775.23842214, 1479221.81172454, 
    1507668.38502693, 1536114.95832933, 1564561.53163172,
  0, 28308.0436361392, 56616.0872722784, 84924.13090842, 113232.174544562, 
    141540.218180701, 169848.261816842, 198156.305452984, 226464.349089123, 
    254772.392725265, 283080.436361406, 311388.479997545, 339696.523633687, 
    368004.567269829, 396312.610905968, 424620.654542109, 452928.698178251, 
    481236.74181439, 509544.785450531, 537852.829086672, 566160.872722814, 
    594468.916358954, 622776.959995094, 651085.003631236, 679393.047267376, 
    707701.090903517, 736009.134539658, 764317.178175799, 792625.221811939, 
    820933.265448081, 849241.309084221, 877549.352720362, 905857.396356503, 
    934165.439992644, 962473.483628784, 990781.527264926, 1019089.57090107, 
    1047397.61453721, 1075705.65817335, 1104013.70180949, 1132321.74544563, 
    1160629.78908177, 1188937.83271791, 1217245.87635405, 1245553.91999019, 
    1273861.96362633, 1302170.00726247, 1330478.05089862, 1358786.09453476, 
    1387094.1381709, 1415402.18180704, 1443710.22544318, 1472018.26907932, 
    1500326.31271546, 1528634.3563516, 1556942.39998774,
  0, 28168.5558495808, 56337.1116991616, 84505.6675487449, 112674.223398328, 
    140842.779247909, 169011.335097492, 197179.890947075, 225348.446796656, 
    253517.002646239, 281685.558495823, 309854.114345403, 338022.670194987, 
    366191.22604457, 394359.781894151, 422528.337743734, 450696.893593317, 
    478865.449442898, 507034.00529248, 535202.561142063, 563371.116991646, 
    591539.672841228, 619708.228690811, 647876.784540394, 676045.340389976, 
    704213.896239558, 732382.452089141, 760551.007938723, 788719.563788305, 
    816888.119637888, 845056.67548747, 873225.231337052, 901393.787186635, 
    929562.343036217, 957730.8988858, 985899.454735383, 1014068.01058496, 
    1042236.56643455, 1070405.12228413, 1098573.67813371, 1126742.23398329, 
    1154910.78983288, 1183079.34568246, 1211247.90153204, 1239416.45738162, 
    1267585.01323121, 1295753.56908079, 1323922.12493037, 1352090.68077995, 
    1380259.23662954, 1408427.79247912, 1436596.3483287, 1464764.90417828, 
    1492933.46002787, 1521102.01587745, 1549270.57172703,
  0, 28028.1146639146, 56056.2293278291, 84084.3439917461, 112112.458655663, 
    140140.573319578, 168168.687983495, 196196.802647412, 224224.917311326, 
    252253.031975243, 280281.14663916, 308309.261303075, 336337.375966991, 
    364365.490630908, 392393.605294823, 420421.71995874, 448449.834622657, 
    476477.949286571, 504506.063950487, 532534.178614404, 560562.293278321, 
    588590.407942237, 616618.522606153, 644646.637270069, 672674.751933985, 
    700702.866597901, 728730.981261818, 756759.095925734, 784787.21058965, 
    812815.325253566, 840843.439917482, 868871.554581398, 896899.669245315, 
    924927.783909231, 952955.898573146, 980984.013237063, 1009012.12790098, 
    1037040.24256489, 1065068.35722881, 1093096.47189273, 1121124.58655664, 
    1149152.70122056, 1177180.81588448, 1205208.93054839, 1233237.04521231, 
    1261265.15987622, 1289293.27454014, 1317321.38920406, 1345349.50386797, 
    1373377.61853189, 1401405.7331958, 1429433.84785972, 1457461.96252364, 
    1485490.07718755, 1513518.19185147, 1541546.30651538,
  0, 27886.7248326051, 55773.4496652101, 83660.1744978176, 111546.899330425, 
    139433.62416303, 167320.348995637, 195207.073828245, 223093.79866085, 
    250980.523493457, 278867.248326065, 306753.97315867, 334640.697991277, 
    362527.422823885, 390414.14765649, 418300.872489097, 446187.597321705, 
    474074.32215431, 501961.046986916, 529847.771819524, 557734.496652131, 
    585621.221484737, 613507.946317344, 641394.671149951, 669281.395982557, 
    697168.120815163, 725054.845647771, 752941.570480377, 780828.295312983, 
    808715.020145591, 836601.744978197, 864488.469810803, 892375.194643411, 
    920261.919476017, 948148.644308623, 976035.369141231, 1003922.09397384, 
    1031808.81880644, 1059695.54363905, 1087582.26847166, 1115468.99330426, 
    1143355.71813687, 1171242.44296948, 1199129.16780208, 1227015.89263469, 
    1254902.6174673, 1282789.3422999, 1310676.06713251, 1338562.79196512, 
    1366449.51679772, 1394336.24163033, 1422222.96646294, 1450109.69129554, 
    1477996.41612815, 1505883.14096076, 1533769.86579336,
  0, 27744.3911412245, 55488.7822824491, 83233.173423676, 110977.564564903, 
    138721.955706127, 166466.346847354, 194210.737988581, 221955.129129806, 
    249699.520271033, 277443.91141226, 305188.302553484, 332932.693694711, 
    360677.084835938, 388421.475977163, 416165.86711839, 443910.258259616, 
    471654.649400841, 499399.040542067, 527143.431683294, 554887.822824521, 
    582632.213965746, 610376.605106972, 638120.996248199, 665865.387389425, 
    693609.778530651, 721354.169671877, 749098.560813103, 776842.951954329, 
    804587.343095556, 832331.734236782, 860076.125378007, 887820.516519234, 
    915564.90766046, 943309.298801686, 971053.689942913, 998798.081084138, 
    1026542.47222536, 1054286.86336659, 1082031.25450782, 1109775.64564904, 
    1137520.03679027, 1165264.4279315, 1193008.81907272, 1220753.21021395, 
    1248497.60135517, 1276241.9924964, 1303986.38363763, 1331730.77477885, 
    1359475.16592008, 1387219.5570613, 1414963.94820253, 1442708.33934376, 
    1470452.73048498, 1498197.12162621, 1525941.51276743,
  0, 27601.1184072908, 55202.2368145816, 82803.3552218747, 110404.473629168, 
    138005.592036459, 165606.710443752, 193207.828851045, 220808.947258336, 
    248410.065665629, 276011.184072922, 303612.302480213, 331213.420887506, 
    358814.539294799, 386415.65770209, 414016.776109383, 441617.894516676, 
    469219.012923967, 496820.131331259, 524421.249738552, 552022.368145845, 
    579623.486553137, 607224.604960429, 634825.723367722, 662426.841775015, 
    690027.960182307, 717629.0785896, 745230.196996892, 772831.315404184, 
    800432.433811477, 828033.552218769, 855634.670626061, 883235.789033354, 
    910836.907440646, 938438.025847938, 966039.144255231, 993640.262662523, 
    1021241.38106982, 1048842.49947711, 1076443.6178844, 1104044.73629169, 
    1131645.85469899, 1159246.97310628, 1186848.09151357, 1214449.20992086, 
    1242050.32832815, 1269651.44673545, 1297252.56514274, 1324853.68355003, 
    1352454.80195732, 1380055.92036462, 1407657.03877191, 1435258.1571792, 
    1462859.27558649, 1490460.39399378, 1518061.51240108,
  0, 27456.9114801041, 54913.8229602082, 82370.7344403146, 109827.645920421, 
    137284.557400525, 164741.468880631, 192198.380360738, 219655.291840842, 
    247112.203320948, 274569.114801055, 302026.026281159, 329482.937761265, 
    356939.849241372, 384396.760721476, 411853.672201582, 439310.583681689, 
    466767.495161793, 494224.406641898, 521681.318122004, 549138.229602111, 
    576595.141082216, 604052.052562321, 631508.964042428, 658965.875522533, 
    686422.787002638, 713879.698482745, 741336.60996285, 768793.521442955, 
    796250.432923062, 823707.344403167, 851164.255883272, 878621.167363378, 
    906078.078843484, 933534.990323589, 960991.901803695, 988448.813283801, 
    1015905.72476391, 1043362.63624401, 1070819.54772412, 1098276.45920422, 
    1125733.37068433, 1153190.28216443, 1180647.19364454, 1208104.10512465, 
    1235561.01660475, 1263017.92808486, 1290474.83956496, 1317931.75104507, 
    1345388.66252517, 1372845.57400528, 1400302.48548538, 1427759.39696549, 
    1455216.3084456, 1482673.2199257, 1510130.13140581,
  0, 27311.775240583, 54623.550481166, 81935.3257217513, 109247.100962337, 
    136558.87620292, 163870.651443505, 191182.42668409, 218494.201924673, 
    245805.977165259, 273117.752405844, 300429.527646427, 327741.302887012, 
    355053.078127598, 382364.853368181, 409676.628608766, 436988.403849351, 
    464300.179089934, 491611.954330518, 518923.729571104, 546235.504811689, 
    573547.280052273, 600859.055292858, 628170.830533443, 655482.605774027, 
    682794.381014611, 710106.156255197, 737417.931495781, 764729.706736365, 
    792041.48197695, 819353.257217534, 846665.032458118, 873976.807698704, 
    901288.582939288, 928600.358179872, 955912.133420457, 983223.908661042, 
    1010535.68390163, 1037847.45914221, 1065159.2343828, 1092471.00962338, 
    1119782.78486396, 1147094.56010455, 1174406.33534513, 1201718.11058572, 
    1229029.8858263, 1256341.66106689, 1283653.43630747, 1310965.21154806, 
    1338276.98678864, 1365588.76202923, 1392900.53726981, 1420212.31251039, 
    1447524.08775098, 1474835.86299156, 1502147.63823215,
  0, 27165.7146010993, 54331.4292021987, 81497.1438033003, 108662.858404402, 
    135828.573005501, 162994.287606603, 190160.002207705, 217325.716808804, 
    244491.431409906, 271657.146011007, 298822.860612107, 325988.575213208, 
    353154.28981431, 380320.004415409, 407485.719016511, 434651.433617612, 
    461817.148218712, 488982.862819812, 516148.577420914, 543314.292022016, 
    570480.006623116, 597645.721224217, 624811.435825318, 651977.150426419, 
    679142.865027519, 706308.579628621, 733474.294229721, 760640.008830822, 
    787805.723431923, 814971.438033024, 842137.152634124, 869302.867235226, 
    896468.581836327, 923634.296437427, 950800.011038529, 977965.725639629, 
    1005131.44024073, 1032297.15484183, 1059462.86944293, 1086628.58404403, 
    1113794.29864513, 1140960.01324623, 1168125.72784733, 1195291.44244844, 
    1222457.15704954, 1249622.87165064, 1276788.58625174, 1303954.30085284, 
    1331120.01545394, 1358285.73005504, 1385451.44465614, 1412617.15925724, 
    1439782.87385834, 1466948.58845944, 1494114.30306054,
  0, 27018.7345053117, 54037.4690106233, 81056.2035159373, 108074.938021251, 
    135093.672526563, 162112.407031877, 189131.141537191, 216149.876042502, 
    243168.610547816, 270187.34505313, 297206.079558442, 324224.814063756, 
    351243.54856907, 378262.283074382, 405281.017579696, 432299.752085009, 
    459318.486590321, 486337.221095634, 513355.955600948, 540374.690106262, 
    567393.424611575, 594412.159116887, 621430.893622201, 648449.628127514, 
    675468.362632827, 702487.097138141, 729505.831643454, 756524.566148767, 
    783543.300654081, 810562.035159393, 837580.769664706, 864599.50417002, 
    891618.238675333, 918636.973180646, 945655.70768596, 972674.442191273, 
    999693.176696585, 1026711.9112019, 1053730.64570721, 1080749.38021252, 
    1107768.11471784, 1134786.84922315, 1161805.58372846, 1188824.31823378, 
    1215843.05273909, 1242861.7872444, 1269880.52174972, 1296899.25625503, 
    1323917.99076034, 1350936.72526566, 1377955.45977097, 1404974.19427628, 
    1431992.9287816, 1459011.66328691, 1486030.39779222,
  0, 26870.8399279981, 53741.6798559961, 80612.5197839965, 107483.359711997, 
    134354.199639995, 161225.039567995, 188095.879495996, 214966.719423994, 
    241837.559351994, 268708.399279994, 295579.239207992, 322450.079135993, 
    349320.919063993, 376191.758991991, 403062.598919992, 429933.438847992, 
    456804.27877599, 483675.118703989, 510545.95863199, 537416.79855999, 
    564287.638487989, 591158.478415988, 618029.318343989, 644900.158271988, 
    671770.998199987, 698641.838127987, 725512.678055987, 752383.517983986, 
    779254.357911986, 806125.197839986, 832996.037767985, 859866.877695985, 
    886737.717623984, 913608.557551984, 940479.397479984, 967350.237407983, 
    994221.077335983, 1021091.91726398, 1047962.75719198, 1074833.59711998, 
    1101704.43704798, 1128575.27697598, 1155446.11690398, 1182316.95683198, 
    1209187.79675998, 1236058.63668798, 1262929.47661598, 1289800.31654398, 
    1316671.15647198, 1343541.99639998, 1370412.83632798, 1397283.67625598, 
    1424154.51618398, 1451025.35611198, 1477896.19603997,
  0, 26722.0358748878, 53444.0717497756, 80166.1076246656, 106888.143499556, 
    133610.179374443, 160332.215249334, 187054.251124224, 213776.286999111, 
    240498.322874001, 267220.358748892, 293942.394623779, 320664.430498669, 
    347386.466373559, 374108.502248447, 400830.538123337, 427552.573998227, 
    454274.609873115, 480996.645748004, 507718.681622894, 534440.717497784, 
    561162.753372673, 587884.789247562, 614606.825122452, 641328.860997341, 
    668050.89687223, 694772.93274712, 721494.968622009, 748217.004496898, 
    774939.040371788, 801661.076246677, 828383.112121566, 855105.147996456, 
    881827.183871345, 908549.219746234, 935271.255621124, 961993.291496013, 
    988715.327370902, 1015437.36324579, 1042159.39912068, 1068881.43499557, 
    1095603.47087046, 1122325.50674535, 1149047.54262024, 1175769.57849513, 
    1202491.61437002, 1229213.65024491, 1255935.6861198, 1282657.72199468, 
    1309379.75786957, 1336101.79374446, 1362823.82961935, 1389545.86549424, 
    1416267.90136913, 1442989.93724402, 1469711.97311891,
  0, 26572.3273824917, 53144.6547649834, 79716.9821474774, 106289.309529971, 
    132861.636912463, 159433.964294957, 186006.291677451, 212578.619059943, 
    239150.946442437, 265723.273824931, 292295.601207422, 318867.928589916, 
    345440.25597241, 372012.583354902, 398584.910737396, 425157.23811989, 
    451729.565502382, 478301.892884875, 504874.220267369, 531446.547649863, 
    558018.875032356, 584591.202414848, 611163.529797342, 637735.857179835, 
    664308.184562328, 690880.511944822, 717452.839327315, 744025.166709808, 
    770597.494092302, 797169.821474795, 823742.148857287, 850314.476239781, 
    876886.803622274, 903459.131004767, 930031.458387261, 956603.785769754, 
    983176.113152247, 1009748.44053474, 1036320.76791723, 1062893.09529973, 
    1089465.42268222, 1116037.75006471, 1142610.07744721, 1169182.4048297, 
    1195754.73221219, 1222327.05959469, 1248899.38697718, 1275471.71435967, 
    1302044.04174217, 1328616.36912466, 1355188.69650715, 1381761.02388965, 
    1408333.35127214, 1434905.67865463, 1461478.00603712,
  0, 26421.7195179319, 52843.4390358639, 79265.158553798, 105686.878071732, 
    132108.597589664, 158530.317107598, 184952.036625533, 211373.756143464, 
    237795.475661399, 264217.195179333, 290638.914697265, 317060.634215199, 
    343482.353733133, 369904.073251065, 396325.792768999, 422747.512286933, 
    449169.231804865, 475590.951322799, 502012.670840733, 528434.390358667, 
    554856.1098766, 581277.829394533, 607699.548912467, 634121.2684304, 
    660542.987948333, 686964.707466267, 713386.4269842, 739808.146502133, 
    766229.866020068, 792651.585538001, 819073.305055934, 845495.024573868, 
    871916.744091801, 898338.463609734, 924760.183127668, 951181.902645601, 
    977603.622163534, 1004025.34168147, 1030447.0611994, 1056868.78071733, 
    1083290.50023527, 1109712.2197532, 1136133.93927113, 1162555.65878907, 
    1188977.378307, 1215399.09782494, 1241820.81734287, 1268242.5368608, 
    1294664.25637874, 1321085.97589667, 1347507.6954146, 1373929.41493254, 
    1400351.13445047, 1426772.8539684, 1453194.57348634,
  0, 26270.2173787702, 52540.4347575405, 78810.6521363129, 105080.869515085, 
    131351.086893856, 157621.304272628, 183891.521651401, 210161.739030171, 
    236431.956408943, 262702.173787716, 288972.391166486, 315242.608545258, 
    341512.825924031, 367783.043302801, 394053.260681574, 420323.478060346, 
    446593.695439116, 472863.912817888, 499134.13019666, 525404.347575433, 
    551674.564954204, 577944.782332975, 604214.999711748, 630485.217090519, 
    656755.43446929, 683025.651848063, 709295.869226834, 735566.086605606, 
    761836.303984378, 788106.521363149, 814376.738741921, 840646.956120693, 
    866917.173499465, 893187.390878236, 919457.608257008, 945727.82563578, 
    971998.043014551, 998268.260393323, 1024538.47777209, 1050808.69515087, 
    1077078.91252964, 1103349.12990841, 1129619.34728718, 1155889.56466595, 
    1182159.78204473, 1208429.9994235, 1234700.21680227, 1260970.43418104, 
    1287240.65155981, 1313510.86893858, 1339781.08631735, 1366051.30369613, 
    1392321.5210749, 1418591.73845367, 1444861.95583244,
  0, 26117.8260928355, 52235.652185671, 78353.4782785087, 104471.304371346, 
    130589.130464182, 156706.95655702, 182824.782649857, 208942.608742693, 
    235060.434835531, 261178.260928368, 287296.087021204, 313413.913114042, 
    339531.739206879, 365649.565299715, 391767.391392553, 417885.21748539, 
    444003.043578226, 470120.869671062, 496238.6957639, 522356.521856738, 
    548474.347949574, 574592.174042411, 600710.000135249, 626827.826228085, 
    652945.652320922, 679063.47841376, 705181.304506596, 731299.130599433, 
    757416.956692271, 783534.782785107, 809652.608877944, 835770.434970782, 
    861888.261063618, 888006.087156455, 914123.913249293, 940241.739342129, 
    966359.565434966, 992477.391527804, 1018595.21762064, 1044713.04371348, 
    1070830.86980631, 1096948.69589915, 1123066.52199199, 1149184.34808483, 
    1175302.17417766, 1201420.0002705, 1227537.82636334, 1253655.65245617, 
    1279773.47854901, 1305891.30464185, 1332009.13073468, 1358126.95682752, 
    1384244.78292036, 1410362.60901319, 1436480.43510603,
  0, 25964.5508180502, 51929.1016361004, 77893.6524541528, 103858.203272205, 
    129822.754090255, 155787.304908308, 181751.85572636, 207716.406544411, 
    233680.957362463, 259645.508180515, 285610.058998566, 311574.609816618, 
    337539.16063467, 363503.711452721, 389468.262270773, 415432.813088825, 
    441397.363906876, 467361.914724927, 493326.465542979, 519291.016361032, 
    545255.567179083, 571220.117997134, 597184.668815187, 623149.219633238, 
    649113.770451289, 675078.321269342, 701042.872087393, 727007.422905445, 
    752971.973723497, 778936.524541548, 804901.0753596, 830865.626177652, 
    856830.176995703, 882794.727813755, 908759.278631807, 934723.829449859, 
    960688.38026791, 986652.931085962, 1012617.48190401, 1038582.03272206, 
    1064546.58354012, 1090511.13435817, 1116475.68517622, 1142440.23599427, 
    1168404.78681232, 1194369.33763038, 1220333.88844843, 1246298.43926648, 
    1272262.99008453, 1298227.54090258, 1324192.09172063, 1350156.64253869, 
    1376121.19335674, 1402085.74417479, 1428050.29499284,
  0, 25810.3967422558, 51620.7934845116, 77431.1902267696, 103241.586969028, 
    129051.983711283, 154862.380453541, 180672.777195799, 206483.173938055, 
    232293.570680313, 258103.967422571, 283914.364164827, 309724.760907085, 
    335535.157649343, 361345.554391599, 387155.951133857, 412966.347876115, 
    438776.74461837, 464587.141360627, 490397.538102885, 516207.934845143, 
    542018.3315874, 567828.728329657, 593639.125071915, 619449.521814172, 
    645259.918556429, 671070.315298687, 696880.712040944, 722691.1087832, 
    748501.505525458, 774311.902267715, 800122.299009972, 825932.69575223, 
    851743.092494487, 877553.489236744, 903363.885979002, 929174.282721259, 
    954984.679463516, 980795.076205774, 1006605.47294803, 1032415.86969029, 
    1058226.26643255, 1084036.6631748, 1109847.05991706, 1135657.45665932, 
    1161467.85340157, 1187278.25014383, 1213088.64688609, 1238899.04362835, 
    1264709.4403706, 1290519.83711286, 1316330.23385512, 1342140.63059737, 
    1367951.02733963, 1393761.42408189, 1419571.82082415,
  0, 25655.369083037, 51310.7381660741, 76966.1072491133, 102621.476332152, 
    128276.845415189, 153932.214498229, 179587.583581268, 205242.952664305, 
    230898.321747344, 256553.690830383, 282209.05991342, 307864.42899646, 
    333519.798079499, 359175.167162536, 384830.536245575, 410485.905328614, 
    436141.274411651, 461796.643494689, 487452.012577729, 513107.381660768, 
    538762.750743806, 564418.119826844, 590073.488909883, 615728.857992921, 
    641384.22707596, 667039.596158999, 692694.965242037, 718350.334325075, 
    744005.703408114, 769661.072491152, 795316.441574191, 820971.81065723, 
    846627.179740268, 872282.548823306, 897937.917906345, 923593.286989383, 
    949248.656072422, 974904.025155461, 1000559.3942385, 1026214.76332154, 
    1051870.13240458, 1077525.50148761, 1103180.87057065, 1128836.23965369, 
    1154491.60873673, 1180146.97781977, 1205802.34690281, 1231457.71598585, 
    1257113.08506888, 1282768.45415192, 1308423.82323496, 1334079.192318, 
    1359734.56140104, 1385389.93048408, 1411045.29956711,
  0, 25499.4730875455, 50998.946175091, 76498.4192626386, 101997.892350186, 
    127497.365437732, 152996.838525279, 178496.311612827, 203995.784700373, 
    229495.25778792, 254994.730875468, 280494.203963013, 305993.677050561, 
    331493.150138109, 356992.623225654, 382492.096313202, 407991.56940075, 
    433491.042488295, 458990.515575842, 484489.988663389, 509989.461750937, 
    535488.934838483, 560988.40792603, 586487.881013578, 611987.354101124, 
    637486.827188671, 662986.300276218, 688485.773363765, 713985.246451312, 
    739484.719538859, 764984.192626406, 790483.665713953, 815983.1388015, 
    841482.611889047, 866982.084976593, 892481.558064141, 917981.031151687, 
    943480.504239234, 968979.977326782, 994479.450414328, 1019978.92350188, 
    1045478.39658942, 1070977.86967697, 1096477.34276452, 1121976.81585206, 
    1147476.28893961, 1172975.76202716, 1198475.2351147, 1223974.70820225, 
    1249474.1812898, 1274973.65437734, 1300473.12746489, 1325972.60055244, 
    1351472.07363999, 1376971.54672753, 1402471.01981508,
  0, 25342.7140323219, 50685.4280646437, 76028.1420969678, 101370.856129292, 
    126713.570161614, 152056.284193938, 177398.998226262, 202741.712258584, 
    228084.426290908, 253427.140323232, 278769.854355554, 304112.568387878, 
    329455.282420202, 354797.996452523, 380140.710484847, 405483.424517171, 
    430826.138549493, 456168.852581816, 481511.56661414, 506854.280646464, 
    532196.994678787, 557539.70871111, 582882.422743434, 608225.136775757, 
    633567.85080808, 658910.564840404, 684253.278872727, 709595.99290505, 
    734938.706937374, 760281.420969697, 785624.13500202, 810966.849034344, 
    836309.563066667, 861652.27709899, 886994.991131314, 912337.705163637, 
    937680.41919596, 963023.133228284, 988365.847260607, 1013708.56129293, 
    1039051.27532525, 1064393.98935758, 1089736.7033899, 1115079.41742222, 
    1140422.13145455, 1165764.84548687, 1191107.55951919, 1216450.27355152, 
    1241792.98758384, 1267135.70161616, 1292478.41564849, 1317821.12968081, 
    1343163.84371313, 1368506.55774546, 1393849.27177778,
  0, 25185.0972231174, 50370.1944462349, 75555.2916693545, 100740.388892474, 
    125925.486115592, 151110.583338711, 176295.680561831, 201480.777784948, 
    226665.875008068, 251850.972231187, 277036.069454305, 302221.166677424, 
    327406.263900544, 352591.361123661, 377776.458346781, 402961.5555699, 
    428146.652793018, 453331.750016136, 478516.847239256, 503701.944462376, 
    528887.041685494, 554072.138908613, 579257.236131732, 604442.333354851, 
    629627.430577969, 654812.527801089, 679997.625024207, 705182.722247326, 
    730367.819470445, 755552.916693564, 780738.013916682, 805923.111139802, 
    831108.20836292, 856293.305586039, 881478.402809158, 906663.500032277, 
    931848.597255395, 957033.694478515, 982218.791701633, 1007403.88892475, 
    1032588.98614787, 1057774.08337099, 1082959.18059411, 1108144.27781723, 
    1133329.37504035, 1158514.47226347, 1183699.56948658, 1208884.6667097, 
    1234069.76393282, 1259254.86115594, 1284439.95837906, 1309625.05560218, 
    1334810.1528253, 1359995.25004842, 1385180.34727153,
  0, 25026.6279947144, 50053.2559894288, 75079.8839841453, 100106.511978862, 
    125133.139973576, 150159.767968293, 175186.395963009, 200213.023957724, 
    225239.65195244, 250266.279947157, 275292.907941871, 300319.535936588, 
    325346.163931304, 350372.791926019, 375399.419920735, 400426.047915452, 
    425452.675910166, 450479.303904882, 475505.931899598, 500532.559894315, 
    525559.18788903, 550585.815883746, 575612.443878462, 600639.071873178, 
    625665.699867893, 650692.32786261, 675718.955857325, 700745.583852041, 
    725772.211846757, 750798.839841473, 775825.467836188, 800852.095830905, 
    825878.72382562, 850905.351820336, 875931.979815052, 900958.607809768, 
    925985.235804483, 951011.8637992, 976038.491793915, 1001065.11978863, 
    1026091.74778335, 1051118.37577806, 1076145.00377278, 1101171.63176749, 
    1126198.25976221, 1151224.88775693, 1176251.51575164, 1201278.14374636, 
    1226304.77174107, 1251331.39973579, 1276358.0277305, 1301384.65572522, 
    1326411.28371994, 1351437.91171465, 1376464.53970937,
  0, 24867.3117107454, 49734.6234214907, 74601.9351322382, 99469.2468429856, 
    124336.558553731, 149203.870264478, 174071.181975226, 198938.493685971, 
    223805.805396719, 248673.117107466, 273540.428818212, 298407.740528959, 
    323275.052239707, 348142.363950452, 373009.675661199, 397876.987371947, 
    422744.299082692, 447611.610793439, 472478.922504186, 497346.234214934, 
    522213.54592568, 547080.857636426, 571948.169347174, 596815.48105792, 
    621682.792768667, 646550.104479414, 671417.416190161, 696284.727900907, 
    721152.039611655, 746019.351322401, 770886.663033147, 795753.974743895, 
    820621.286454641, 845488.598165388, 870355.909876135, 895223.221586882, 
    920090.533297628, 944957.845008376, 969825.156719122, 994692.468429868, 
    1019559.78014062, 1044427.09185136, 1069294.40356211, 1094161.71527286, 
    1119029.0269836, 1143896.33869435, 1168763.6504051, 1193630.96211584, 
    1218498.27382659, 1243365.58553734, 1268232.89724808, 1293100.20895883, 
    1317967.52066958, 1342834.83238032, 1367702.14409107 ;

 x_psi =
  16013.5632895756, 48040.6898687267, 80067.8164478792, 112094.943027033, 
    144122.069606186, 176149.196185338, 208176.322764492, 240203.449343645, 
    272230.575922797, 304257.702501951, 336284.829081103, 368311.955660256, 
    400339.08223941, 432366.208818562, 464393.335397715, 496420.461976869, 
    528447.588556021, 560474.715135173, 592501.841714326, 624528.96829348, 
    656556.094872633, 688583.221451786, 720610.348030939, 752637.474610092, 
    784664.601189245, 816691.727768398, 848718.854347551, 880745.980926704, 
    912773.107505857, 944800.23408501, 976827.360664163, 1008854.48724332, 
    1040881.61382247, 1072908.74040162, 1104935.86698078, 1136962.99355993, 
    1168990.12013908, 1201017.24671823, 1233044.37329739, 1265071.49987654, 
    1297098.62645569, 1329125.75303485, 1361152.879614, 1393180.00619315, 
    1425207.13277231, 1457234.25935146, 1489261.38593061, 1521288.51250976, 
    1553315.63908892, 1585342.76566807, 1617369.89224722, 1649397.01882638, 
    1681424.14540553, 1713451.27198468, 1745478.39856383,
  15959.142777148, 47877.4283314439, 79795.7138857412, 111713.99944004, 
    143632.284994337, 175550.570548634, 207468.856102933, 239387.14165723, 
    271305.427211528, 303223.712765826, 335141.998320124, 367060.283874421, 
    398978.56942872, 430896.854983017, 462815.140537314, 494733.426091613, 
    526651.71164591, 558569.997200207, 590488.282754505, 622406.568308803, 
    654324.853863101, 686243.139417398, 718161.424971696, 750079.710525995, 
    781997.996080292, 813916.28163459, 845834.567188888, 877752.852743185, 
    909671.138297483, 941589.423851781, 973507.709406078, 1005425.99496038, 
    1037344.28051467, 1069262.56606897, 1101180.85162327, 1133099.13717757, 
    1165017.42273186, 1196935.70828616, 1228853.99384046, 1260772.27939476, 
    1292690.56494906, 1324608.85050335, 1356527.13605765, 1388445.42161195, 
    1420363.70716625, 1452281.99272054, 1484200.27827484, 1516118.56382914, 
    1548036.84938344, 1579955.13493774, 1611873.42049203, 1643791.70604633, 
    1675709.99160063, 1707628.27715493, 1739546.56270922,
  15904.1821070796, 47712.5463212389, 79520.9105353996, 111329.274749562, 
    143137.638963722, 174946.003177883, 206754.367392045, 238562.731606206, 
    270371.095820366, 302179.460034528, 333987.824248689, 365796.188462849, 
    397604.552677011, 429412.916891172, 461221.281105333, 493029.645319495, 
    524838.009533655, 556646.373747815, 588454.737961977, 620263.102176139, 
    652071.4663903, 683879.830604461, 715688.194818622, 747496.559032783, 
    779304.923246944, 811113.287461105, 842921.651675267, 874730.015889427, 
    906538.380103589, 938346.74431775, 970155.10853191, 1001963.47274607, 
    1033771.83696023, 1065580.20117439, 1097388.56538856, 1129196.92960272, 
    1161005.29381688, 1192813.65803104, 1224622.0222452, 1256430.38645936, 
    1288238.75067352, 1320047.11488768, 1351855.47910184, 1383663.843316, 
    1415472.20753017, 1447280.57174433, 1479088.93595849, 1510897.30017265, 
    1542705.66438681, 1574514.02860097, 1606322.39281513, 1638130.75702929, 
    1669939.12124345, 1701747.48545761, 1733555.84967178,
  15848.6831396159, 47546.0494188478, 79243.415698081, 110940.781977316, 
    142638.148256549, 174335.514535782, 206032.880815017, 237730.24709425, 
    269427.613373483, 301124.979652718, 332822.345931951, 364519.712211184, 
    396217.078490419, 427914.444769652, 459611.811048885, 491309.17732812, 
    523006.543607353, 554703.909886585, 586401.276165819, 618098.642445054, 
    649796.008724288, 681493.375003521, 713190.741282755, 744888.107561989, 
    776585.473841222, 808282.840120456, 839980.20639969, 871677.572678923, 
    903374.938958157, 935072.305237391, 966769.671516624, 998467.037795858, 
    1030164.40407509, 1061861.77035432, 1093559.13663356, 1125256.50291279, 
    1156953.86919203, 1188651.23547126, 1220348.60175049, 1252045.96802973, 
    1283743.33430896, 1315440.70058819, 1347138.06686743, 1378835.43314666, 
    1410532.7994259, 1442230.16570513, 1473927.53198436, 1505624.8982636, 
    1537322.26454283, 1569019.63082206, 1600716.9971013, 1632414.36338053, 
    1664111.72965976, 1695809.095939, 1727506.46221823,
  15792.6477532215, 47377.9432596645, 78963.2387661088, 110548.534272554, 
    142133.829778999, 173719.125285443, 205304.420791889, 236889.716298333, 
    268475.011804777, 300060.307311223, 331645.602817667, 363230.898324112, 
    394816.193830557, 426401.489337002, 457986.784843446, 489572.080349892, 
    521157.375856336, 552742.67136278, 584327.966869225, 615913.26237567, 
    647498.557882115, 679083.85338856, 710669.148895005, 742254.44440145, 
    773839.739907894, 805425.035414339, 837010.330920784, 868595.626427228, 
    900180.921933673, 931766.217440118, 963351.512946562, 994936.808453007, 
    1026522.10395945, 1058107.3994659, 1089692.69497234, 1121277.99047879, 
    1152863.28598523, 1184448.58149168, 1216033.87699812, 1247619.17250457, 
    1279204.46801101, 1310789.76351746, 1342375.0590239, 1373960.35453034, 
    1405545.65003679, 1437130.94554323, 1468716.24104968, 1500301.53655612, 
    1531886.83206257, 1563472.12756901, 1595057.42307546, 1626642.7185819, 
    1658228.01408835, 1689813.30959479, 1721398.60510124,
  15736.0778445167, 47208.2335335502, 78680.3892225849, 110152.544911621, 
    141624.700600656, 173096.856289691, 204569.011978727, 236041.167667762, 
    267513.323356796, 298985.479045832, 330457.634734867, 361929.790423902, 
    393401.946112938, 424874.101801973, 456346.257491008, 487818.413180044, 
    519290.568869079, 550762.724558113, 582234.880247148, 613707.035936184, 
    645179.19162522, 676651.347314254, 708123.50300329, 739595.658692325, 
    771067.81438136, 802539.970070396, 834012.125759431, 865484.281448466, 
    896956.437137501, 928428.592826537, 959900.748515572, 991372.904204607, 
    1022845.05989364, 1054317.21558268, 1085789.37127171, 1117261.52696075, 
    1148733.68264978, 1180205.83833882, 1211677.99402785, 1243150.14971689, 
    1274622.30540592, 1306094.46109496, 1337566.61678399, 1369038.77247303, 
    1400510.92816207, 1431983.0838511, 1463455.23954014, 1494927.39522917, 
    1526399.55091821, 1557871.70660724, 1589343.86229628, 1620816.01798531, 
    1652288.17367435, 1683760.32936338, 1715232.48505242,
  15678.9753282136, 47036.9259846408, 78394.8766410693, 109752.827297499, 
    141110.777953928, 172468.728610356, 203826.679266786, 235184.629923215, 
    266542.580579643, 297900.531236073, 329258.481892502, 360616.43254893, 
    391974.38320536, 423332.333861789, 454690.284518217, 486048.235174647, 
    517406.185831076, 548764.136487504, 580122.087143933, 611480.037800363, 
    642837.988456792, 674195.93911322, 705553.889769649, 736911.840426079, 
    768269.791082507, 799627.741738936, 830985.692395366, 862343.643051794, 
    893701.593708223, 925059.544364652, 956417.495021081, 987775.44567751, 
    1019133.39633394, 1050491.34699037, 1081849.2976468, 1113207.24830323, 
    1144565.19895965, 1175923.14961608, 1207281.10027251, 1238639.05092894, 
    1269997.00158537, 1301354.9522418, 1332712.90289823, 1364070.85355466, 
    1395428.80421109, 1426786.75486752, 1458144.70552395, 1489502.65618037, 
    1520860.6068368, 1552218.55749323, 1583576.50814966, 1614934.45880609, 
    1646292.40946252, 1677650.36011895, 1709008.31077538,
  15621.3421370508, 46864.0264111525, 78106.7106852555, 109349.39495936, 
    140592.079233463, 171834.763507566, 203077.44778167, 234320.132055773, 
    265562.816329876, 296805.500603981, 328048.184878083, 359290.869152186, 
    390533.553426291, 421776.237700394, 453018.921974497, 484261.606248601, 
    515504.290522704, 546746.974796806, 577989.65907091, 609232.343345014, 
    640475.027619118, 671717.711893221, 702960.396167325, 734203.080441428, 
    765445.764715531, 796688.448989635, 827931.133263739, 859173.817537842, 
    890416.501811945, 921659.186086049, 952901.870360152, 984144.554634256, 
    1015387.23890836, 1046629.92318246, 1077872.60745657, 1109115.29173067, 
    1140357.97600477, 1171600.66027888, 1202843.34455298, 1234086.02882708, 
    1265328.71310119, 1296571.39737529, 1327814.08164939, 1359056.7659235, 
    1390299.4501976, 1421542.1344717, 1452784.81874581, 1484027.50301991, 
    1515270.18729401, 1546512.87156812, 1577755.55584222, 1608998.24011632, 
    1640240.92439043, 1671483.60866453, 1702726.29293863,
  15563.1802217284, 46689.5406651853, 77815.9011086435, 108942.261552103, 
    140068.621995561, 171194.982439019, 202321.342882479, 233447.703325937, 
    264574.063769395, 295700.424212855, 326826.784656313, 357953.145099771, 
    389079.505543231, 420205.865986689, 451332.226430147, 482458.586873606, 
    513584.947317065, 544711.307760522, 575837.668203981, 606964.02864744, 
    638090.389090899, 669216.749534358, 700343.109977816, 731469.470421275, 
    762595.830864734, 793722.191308192, 824848.551751651, 855974.912195109, 
    887101.272638568, 918227.633082027, 949353.993525485, 980480.353968944, 
    1011606.7144124, 1042733.07485586, 1073859.43529932, 1104985.79574278, 
    1136112.15618624, 1167238.5166297, 1198364.87707315, 1229491.23751661, 
    1260617.59796007, 1291743.95840353, 1322870.31884699, 1353996.67929045, 
    1385123.03973391, 1416249.40017736, 1447375.76062082, 1478502.12106428, 
    1509628.48150774, 1540754.8419512, 1571881.20239466, 1603007.56283812, 
    1634133.92328158, 1665260.28372503, 1696386.64416849,
  15504.4915508417, 46513.474652525, 77522.4577542097, 108531.440855896, 
    139540.42395758, 170549.407059265, 201558.390160951, 232567.373262636, 
    263576.35636432, 294585.339466006, 325594.322567691, 356603.305669376, 
    387612.288771062, 418621.271872746, 449630.254974431, 480639.238076117, 
    511648.221177802, 542657.204279486, 573666.187381171, 604675.170482857, 
    635684.153584542, 666693.136686227, 697702.119787912, 728711.102889598, 
    759720.085991282, 790729.069092968, 821738.052194653, 852747.035296338, 
    883756.018398023, 914765.001499709, 945773.984601393, 976782.967703079, 
    1007791.95080476, 1038800.93390645, 1069809.91700813, 1100818.90010982, 
    1131827.8832115, 1162836.86631319, 1193845.84941487, 1224854.83251656, 
    1255863.81561824, 1286872.79871993, 1317881.78182161, 1348890.7649233, 
    1379899.74802499, 1410908.73112667, 1441917.71422836, 1472926.69733004, 
    1503935.68043173, 1534944.66353341, 1565953.6466351, 1596962.62973678, 
    1627971.61283847, 1658980.59594015, 1689989.57904184,
  15445.2781108145, 46335.8343324435, 77226.3905540739, 108116.946775706, 
    139007.502997336, 169898.059218966, 200788.615440598, 231679.171662228, 
    262569.727883859, 293460.28410549, 324350.840327121, 355241.396548751, 
    386131.952770383, 417022.508992013, 447913.065213643, 478803.621435275, 
    509694.177656905, 540584.733878535, 571475.290100166, 602365.846321797, 
    633256.402543429, 664146.958765059, 695037.51498669, 725928.071208321, 
    756818.627429951, 787709.183651582, 818599.739873213, 849490.296094844, 
    880380.852316475, 911271.408538106, 942161.964759736, 973052.520981367, 
    1003943.077203, 1034833.63342463, 1065724.18964626, 1096614.74586789, 
    1127505.30208952, 1158395.85831115, 1189286.41453278, 1220176.97075441, 
    1251067.52697604, 1281958.08319767, 1312848.63941931, 1343739.19564094, 
    1374629.75186257, 1405520.3080842, 1436410.86430583, 1467301.42052746, 
    1498191.97674909, 1529082.53297072, 1559973.08919235, 1590863.64541398, 
    1621754.20163561, 1652644.75785724, 1683535.31407887,
  15385.5419058323, 46156.6257174968, 76927.7095291626, 107698.79334083, 
    138469.877152496, 169240.960964161, 200012.044775829, 230783.128587494, 
    261554.21239916, 292325.296210827, 323096.380022493, 353867.463834159, 
    384638.547645826, 415409.631457492, 446180.715269158, 476951.799080825, 
    507722.882892491, 538493.966704156, 569265.050515823, 600036.13432749, 
    630807.218139156, 661578.301950822, 692349.385762489, 723120.469574155, 
    753891.553385821, 784662.637197487, 815433.721009154, 846204.80482082, 
    876975.888632486, 907746.972444153, 938518.056255819, 969289.140067485, 
    1000060.22387915, 1030831.30769082, 1061602.39150248, 1092373.47531415, 
    1123144.55912582, 1153915.64293748, 1184686.72674915, 1215457.81056081, 
    1246228.89437248, 1276999.97818415, 1307771.06199581, 1338542.14580748, 
    1369313.22961915, 1400084.31343081, 1430855.39724248, 1461626.48105414, 
    1492397.56486581, 1523168.64867748, 1553939.73248914, 1584710.81630081, 
    1615481.90011248, 1646252.98392414, 1677024.06773581,
  15325.2849577738, 45975.8548733214, 76626.4247888704, 107276.994704421, 
    137927.56461997, 168578.134535518, 199228.704451069, 229879.274366618, 
    260529.844282167, 291180.414197717, 321830.984113266, 352481.554028815, 
    383132.123944365, 413782.693859914, 444433.263775463, 475083.833691013, 
    505734.403606562, 536384.97352211, 567035.54343766, 597686.11335321, 
    628336.68326876, 658987.253184309, 689637.823099858, 720288.393015408, 
    750938.962930957, 781589.532846506, 812240.102762056, 842890.672677605, 
    873541.242593154, 904191.812508704, 934842.382424253, 965492.952339802, 
    996143.522255352, 1026794.0921709, 1057444.66208645, 1088095.232002, 
    1118745.80191755, 1149396.3718331, 1180046.94174865, 1210697.5116642, 
    1241348.08157975, 1271998.6514953, 1302649.22141085, 1333299.79132639, 
    1363950.36124194, 1394600.93115749, 1425251.50107304, 1455902.07098859, 
    1486552.64090414, 1517203.21081969, 1547853.78073524, 1578504.35065079, 
    1609154.92056634, 1639805.49048189, 1670456.06039744,
  15264.5093061431, 45793.5279184294, 76322.546530717, 106851.565143006, 
    137380.583755294, 167909.602367581, 198438.62097987, 228967.639592158, 
    259496.658204445, 290025.676816734, 320554.695429022, 351083.714041309, 
    381612.732653598, 412141.751265886, 442670.769878173, 473199.788490462, 
    503728.80710275, 534257.825715037, 564786.844327325, 595315.862939614, 
    625844.881551902, 656373.90016419, 686902.918776478, 717431.937388766, 
    747960.956001054, 778489.974613342, 809018.993225631, 839548.011837918, 
    870077.030450206, 900606.049062495, 931135.067674782, 961664.086287071, 
    992193.104899359, 1022722.12351165, 1053251.14212393, 1083780.16073622, 
    1114309.17934851, 1144838.1979608, 1175367.21657309, 1205896.23518537, 
    1236425.25379766, 1266954.27240995, 1297483.29102224, 1328012.30963453, 
    1358541.32824682, 1389070.3468591, 1419599.36547139, 1450128.38408368, 
    1480657.40269597, 1511186.42130826, 1541715.43992054, 1572244.45853283, 
    1602773.47714512, 1633302.49575741, 1663831.51436969,
  15203.2170080003, 45609.651024001, 76016.085040003, 106422.519056006, 
    136828.953072008, 167235.38708801, 197641.821104013, 228048.255120015, 
    258454.689136017, 288861.123152021, 319267.557168023, 349673.991184025, 
    380080.425200028, 410486.85921603, 440893.293232032, 471299.727248035, 
    501706.161264037, 532112.595280038, 562519.029296041, 592925.463312044, 
    623331.897328047, 653738.331344049, 684144.765360052, 714551.199376054, 
    744957.633392056, 775364.067408059, 805770.501424062, 836176.935440063, 
    866583.369456066, 896989.803472069, 927396.237488071, 957802.671504073, 
    988209.105520076, 1018615.53953608, 1049021.97355208, 1079428.40756808, 
    1109834.84158409, 1140241.27560009, 1170647.70961609, 1201054.14363209, 
    1231460.5776481, 1261867.0116641, 1292273.4456801, 1322679.8796961, 
    1353086.31371211, 1383492.74772811, 1413899.18174411, 1444305.61576011, 
    1474712.04977611, 1505118.48379212, 1535524.91780812, 1565931.35182412, 
    1596337.78584012, 1626744.21985613, 1657150.65387213,
  15141.4101378919, 45424.2304136757, 75707.0506894607, 105989.870965247, 
    136272.691241032, 166555.511516817, 196838.331792604, 227121.152068389, 
    257403.972344174, 287686.79261996, 317969.612895745, 348252.43317153, 
    378535.253447317, 408818.073723102, 439100.893998887, 469383.714274673, 
    499666.534550458, 529949.354826243, 560232.175102028, 590514.995377815, 
    620797.8156536, 651080.635929385, 681363.456205171, 711646.276480957, 
    741929.096756742, 772211.917032528, 802494.737308313, 832777.557584098, 
    863060.377859884, 893343.19813567, 923626.018411455, 953908.838687241, 
    984191.658963026, 1014474.47923881, 1044757.2995146, 1075040.11979038, 
    1105322.94006617, 1135605.76034195, 1165888.58061774, 1196171.40089352, 
    1226454.22116931, 1256737.0414451, 1287019.86172088, 1317302.68199667, 
    1347585.50227245, 1377868.32254824, 1408151.14282402, 1438433.96309981, 
    1468716.78337559, 1498999.60365138, 1529282.42392716, 1559565.24420295, 
    1589848.06447874, 1620130.88475452, 1650413.70503031,
  15079.0907877805, 45237.2723633415, 75395.4539389038, 105553.635514467, 
    135711.81709003, 165869.998665592, 196028.180241156, 226186.361816718, 
    256344.54339228, 286502.724967844, 316660.906543406, 346819.088118968, 
    376977.269694532, 407135.451270094, 437293.632845657, 467451.81442122, 
    497609.995996782, 527768.177572344, 557926.359147907, 588084.540723471, 
    618242.722299034, 648400.903874596, 678559.085450159, 708717.267025722, 
    738875.448601284, 769033.630176847, 799191.81175241, 829349.993327972, 
    859508.174903535, 889666.356479098, 919824.53805466, 949982.719630223, 
    980140.901205786, 1010299.08278135, 1040457.26435691, 1070615.44593247, 
    1100773.62750804, 1130931.8090836, 1161089.99065916, 1191248.17223472, 
    1221406.35381029, 1251564.53538585, 1281722.71696141, 1311880.89853698, 
    1342039.08011254, 1372197.2616881, 1402355.44326366, 1432513.62483923, 
    1462671.80641479, 1492829.98799035, 1522988.16956591, 1553146.35114148, 
    1583304.53271704, 1613462.7142926, 1643620.89586816,
  15016.2610669743, 45048.7832009229, 75081.3053348729, 105113.827468824, 
    135146.349602774, 165178.871736724, 195211.393870675, 225243.916004625, 
    255276.438138575, 285308.960272526, 315341.482406476, 345374.004540426, 
    375406.526674377, 405439.048808327, 435471.570942277, 465504.093076228, 
    495536.615210178, 525569.137344127, 555601.659478078, 585634.181612029, 
    615666.70374598, 645699.225879929, 675731.74801388, 705764.270147831, 
    735796.792281781, 765829.314415731, 795861.836549682, 825894.358683632, 
    855926.880817582, 885959.402951533, 915991.925085483, 946024.447219433, 
    976056.969353384, 1006089.49148733, 1036122.01362128, 1066154.53575523, 
    1096187.05788918, 1126219.58002314, 1156252.10215709, 1186284.62429104, 
    1216317.14642499, 1246349.66855894, 1276382.19069289, 1306414.71282684, 
    1336447.23496079, 1366479.75709474, 1396512.27922869, 1426544.80136264, 
    1456577.32349659, 1486609.84563054, 1516642.36776449, 1546674.88989844, 
    1576707.41203239, 1606739.93416634, 1636772.45630029,
  14952.9231020554, 44858.7693061663, 74764.6155102784, 104670.461714392, 
    134576.307918504, 164482.154122616, 194388.00032673, 224293.846530842, 
    254199.692734954, 284105.538939067, 314011.385143179, 343917.231347292, 
    373823.077551405, 403728.923755517, 433634.769959629, 463540.616163743, 
    493446.462367855, 523352.308571966, 553258.154776079, 583164.000980193, 
    613069.847184305, 642975.693388417, 672881.53959253, 702787.385796643, 
    732693.232000755, 762599.078204868, 792504.924408981, 822410.770613093, 
    852316.616817205, 882222.463021318, 912128.30922543, 942034.155429543, 
    971940.001633656, 1001845.84783777, 1031751.69404188, 1061657.54024599, 
    1091563.38645011, 1121469.23265422, 1151375.07885833, 1181280.92506244, 
    1211186.77126656, 1241092.61747067, 1270998.46367478, 1300904.30987889, 
    1330810.15608301, 1360716.00228712, 1390621.84849123, 1420527.69469534, 
    1450433.54089946, 1480339.38710357, 1510245.23330768, 1540151.07951179, 
    1570056.92571591, 1599962.77192002, 1629868.61812413,
  14889.079036808, 44667.237110424, 74445.3951840412, 104223.55325766, 
    134001.711331277, 163779.869404894, 193558.027478513, 223336.18555213, 
    253114.343625747, 282892.501699366, 312670.659772983, 342448.8178466, 
    372226.975920219, 402005.133993836, 431783.292067453, 461561.450141072, 
    491339.608214689, 521117.766288306, 550895.924361924, 580674.082435542, 
    610452.24050916, 640230.398582777, 670008.556656395, 699786.714730013, 
    729564.87280363, 759343.030877248, 789121.188950866, 818899.347024483, 
    848677.505098101, 878455.663171719, 908233.821245336, 938011.979318954, 
    967790.137392572, 997568.295466189, 1027346.45353981, 1057124.61161342, 
    1086902.76968704, 1116680.92776066, 1146459.08583428, 1176237.24390789, 
    1206015.40198151, 1235793.56005513, 1265571.71812875, 1295349.87620237, 
    1325128.03427598, 1354906.1923496, 1384684.35042322, 1414462.50849684, 
    1444240.66657045, 1474018.82464407, 1503796.98271769, 1533575.14079131, 
    1563353.29886492, 1593131.45693854, 1622909.61501216,
  14824.7310321456, 44474.1930964367, 74123.6551607291, 103773.117225023, 
    133422.579289315, 163072.041353608, 192721.503417901, 222370.965482194, 
    252020.427546486, 281669.88961078, 311319.351675072, 340968.813739364, 
    370618.275803658, 400267.73786795, 429917.199932243, 459566.661996537, 
    489216.124060829, 518865.586125121, 548515.048189414, 578164.510253707, 
    607813.972318, 637463.434382293, 667112.896446586, 696762.358510879, 
    726411.820575171, 756061.282639464, 785710.744703757, 815360.206768049, 
    845009.668832342, 874659.130896635, 904308.592960928, 933958.05502522, 
    963607.517089513, 993256.979153806, 1022906.4412181, 1052555.90328239, 
    1082205.36534668, 1111854.82741098, 1141504.28947527, 1171153.75153956, 
    1200803.21360386, 1230452.67566815, 1260102.13773244, 1289751.59979673, 
    1319401.06186103, 1349050.52392532, 1378699.98598961, 1408349.44805391, 
    1437998.9101182, 1467648.37218249, 1497297.83424678, 1526947.29631108, 
    1556596.75837537, 1586246.22043966, 1615895.68250395,
  14759.881266038, 44279.643798114, 73799.4063301913, 103319.16886227, 
    132838.931394347, 162358.693926424, 191878.456458503, 221398.21899058, 
    250917.981522658, 280437.744054736, 309957.506586813, 339477.269118891, 
    368997.031650969, 398516.794183046, 428036.556715124, 457556.319247202, 
    487076.08177928, 516595.844311356, 546115.606843434, 575635.369375513, 
    605155.131907591, 634674.894439668, 664194.656971746, 693714.419503824, 
    723234.182035901, 752753.944567979, 782273.707100057, 811793.469632134, 
    841313.232164212, 870832.99469629, 900352.757228367, 929872.519760445, 
    959392.282292523, 988912.0448246, 1018431.80735668, 1047951.56988876, 
    1077471.33242083, 1106991.09495291, 1136510.85748499, 1166030.62001707, 
    1195550.38254914, 1225070.14508122, 1254589.9076133, 1284109.67014538, 
    1313629.43267746, 1343149.19520953, 1372668.95774161, 1402188.72027369, 
    1431708.48280577, 1461228.24533784, 1490748.00786992, 1520267.770402, 
    1549787.53293408, 1579307.29546615, 1608827.05799823,
  14694.5319334378, 44083.5958003134, 73472.6596671902, 102861.723534068, 
    132250.787400945, 161639.851267822, 191028.9151347, 220417.979001577, 
    249807.042868454, 279196.106735332, 308585.170602209, 337974.234469085, 
    367363.298335964, 396752.36220284, 426141.426069717, 455530.489936595, 
    484919.553803472, 514308.617670348, 543697.681537226, 573086.745404104, 
    602475.809270981, 631864.873137858, 661253.937004736, 690643.000871613, 
    720032.06473849, 749421.128605367, 778810.192472245, 808199.256339122, 
    837588.320205999, 866977.384072877, 896366.447939753, 925755.511806631, 
    955144.575673508, 984533.639540385, 1013922.70340726, 1043311.76727414, 
    1072700.83114102, 1102089.89500789, 1131478.95887477, 1160868.02274165, 
    1190257.08660853, 1219646.1504754, 1249035.21434228, 1278424.27820916, 
    1307813.34207604, 1337202.40594291, 1366591.46980979, 1395980.53367667, 
    1425369.59754354, 1454758.66141042, 1484147.7252773, 1513536.78914418, 
    1542925.85301105, 1572314.91687793, 1601703.98074481,
  14628.6852462056, 43886.0557386168, 73143.4262310293, 102400.796723443, 
    131658.167215855, 160915.537708268, 190172.908200682, 219430.278693094, 
    248687.649185507, 277945.01967792, 307202.390170333, 336459.760662745, 
    365717.131155159, 394974.501647571, 424231.872139984, 453489.242632398, 
    482746.61312481, 512003.983617222, 541261.354109635, 570518.724602049, 
    599776.095094462, 629033.465586874, 658290.836079287, 687548.206571701, 
    716805.577064113, 746062.947556526, 775320.318048939, 804577.688541352, 
    833835.059033765, 863092.429526178, 892349.80001859, 921607.170511003, 
    950864.541003416, 980121.911495829, 1009379.28198824, 1038636.65248066, 
    1067894.02297307, 1097151.39346548, 1126408.76395789, 1155666.13445031, 
    1184923.50494272, 1214180.87543513, 1243438.24592755, 1272695.61641996, 
    1301952.98691237, 1331210.35740478, 1360467.7278972, 1389725.09838961, 
    1418982.46888202, 1448239.83937444, 1477497.20986685, 1506754.58035926, 
    1536011.95085167, 1565269.32134409, 1594526.6918365,
  14562.3434330356, 43687.0302991068, 72811.7171651792, 101936.404031253, 
    131061.090897325, 160185.777763398, 189310.464629471, 218435.151495544, 
    247559.838361616, 276684.52522769, 305809.212093762, 334933.898959835, 
    364058.585825908, 393183.272691981, 422307.959558053, 451432.646424127, 
    480557.333290199, 509682.020156271, 538806.707022344, 567931.393888418, 
    597056.080754491, 626180.767620563, 655305.454486636, 684430.141352709, 
    713554.828218782, 742679.515084855, 771804.201950928, 800928.888817, 
    830053.575683073, 859178.262549146, 888302.949415219, 917427.636281292, 
    946552.323147365, 975677.010013437, 1004801.69687951, 1033926.38374558, 
    1063051.07061166, 1092175.75747773, 1121300.4443438, 1150425.13120987, 
    1179549.81807595, 1208674.50494202, 1237799.19180809, 1266923.87867417, 
    1296048.56554024, 1325173.25240631, 1354297.93927238, 1383422.62613846, 
    1412547.31300453, 1441671.9998706, 1470796.68673667, 1499921.37360275, 
    1529046.06046882, 1558170.74733489, 1587295.43420097,
  14495.5087393798, 43486.5262181394, 72477.5436969002, 101468.561175662, 
    130459.578654423, 159450.596133184, 188441.613611946, 217432.631090707, 
    246423.648569468, 275414.66604823, 304405.683526991, 333396.701005751, 
    362387.718484513, 391378.735963274, 420369.753442035, 449360.770920797, 
    478351.788399558, 507342.805878318, 536333.82335708, 565324.840835842, 
    594315.858314603, 623306.875793364, 652297.893272126, 681288.910750887, 
    710279.928229648, 739270.945708409, 768261.963187171, 797252.980665931, 
    826243.998144693, 855235.015623454, 884226.033102215, 913217.050580976, 
    942208.068059738, 971199.085538499, 1000190.10301726, 1029181.12049602, 
    1058172.13797478, 1087163.15545354, 1116154.17293231, 1145145.19041107, 
    1174136.20788983, 1203127.22536859, 1232118.24284735, 1261109.26032611, 
    1290100.27780487, 1319091.29528363, 1348082.3127624, 1377073.33024116, 
    1406064.34771992, 1435055.36519868, 1464046.38267744, 1493037.4001562, 
    1522028.41763496, 1551019.43511372, 1580010.45259248,
  14428.1834273723, 43284.5502821168, 72140.9171368626, 100997.28399161, 
    129853.650846355, 158710.017701101, 187566.384555848, 216422.751410594, 
    245279.11826534, 274135.485120087, 302991.851974832, 331848.218829578, 
    360704.585684325, 389560.952539071, 418417.319393817, 447273.686248563, 
    476130.053103309, 504986.419958054, 533842.786812801, 562699.153667548, 
    591555.520522294, 620411.88737704, 649268.254231786, 678124.621086532, 
    706980.987941278, 735837.354796025, 764693.721650771, 793550.088505517, 
    822406.455360263, 851262.822215009, 880119.189069755, 908975.555924502, 
    937831.922779248, 966688.289633994, 995544.65648874, 1024401.02334349, 
    1053257.39019823, 1082113.75705298, 1110970.12390772, 1139826.49076247, 
    1168682.85761722, 1197539.22447196, 1226395.59132671, 1255251.95818146, 
    1284108.3250362, 1312964.69189095, 1341821.05874569, 1370677.42560044, 
    1399533.79245519, 1428390.15930993, 1457246.52616468, 1486102.89301942, 
    1514959.25987417, 1543815.62672892, 1572671.99358366,
  14360.3697757524, 43081.1093272572, 71801.8488787632, 100522.58843027, 
    129243.327981776, 157964.067533282, 186684.80708479, 215405.546636296, 
    244126.286187802, 272847.025739309, 301567.765290815, 330288.504842321, 
    359009.244393828, 387729.983945334, 416450.72349684, 445171.463048347, 
    473892.202599853, 502612.942151359, 531333.681702865, 560054.421254372, 
    588775.160805879, 617495.900357385, 646216.639908892, 674937.379460398, 
    703658.119011904, 732378.858563411, 761099.598114917, 789820.337666423, 
    818541.07721793, 847261.816769436, 875982.556320942, 904703.295872449, 
    933424.035423956, 962144.774975462, 990865.514526968, 1019586.25407847, 
    1048306.99362998, 1077027.73318149, 1105748.47273299, 1134469.2122845, 
    1163189.95183601, 1191910.69138751, 1220631.43093902, 1249352.17049053, 
    1278072.91004203, 1306793.64959354, 1335514.38914504, 1364235.12869655, 
    1392955.86824806, 1421676.60779956, 1450397.34735107, 1479118.08690258, 
    1507838.82645408, 1536559.56600559, 1565280.3055571,
  14292.0700797878, 42876.2102393634, 71460.3503989402, 100044.490558518, 
    128628.630718095, 157212.770877672, 185796.91103725, 214381.051196827, 
    242965.191356404, 271549.331515982, 300133.471675558, 328717.611835135, 
    357301.751994713, 385885.89215429, 414470.032313867, 443054.172473445, 
    471638.312633022, 500222.452792598, 528806.592952176, 557390.733111754, 
    585974.873271331, 614559.013430908, 643143.153590485, 671727.293750063, 
    700311.433909639, 728895.574069217, 757479.714228794, 786063.854388371, 
    814647.994547949, 843232.134707526, 871816.274867103, 900400.41502668, 
    928984.555186258, 957568.695345834, 986152.835505412, 1014736.97566499, 
    1043321.11582457, 1071905.25598414, 1100489.39614372, 1129073.5363033, 
    1157657.67646287, 1186241.81662245, 1214825.95678203, 1243410.09694161, 
    1271994.23710118, 1300578.37726076, 1329162.51742034, 1357746.65757992, 
    1386330.79773949, 1414914.93789907, 1443499.07805865, 1472083.21821822, 
    1500667.3583778, 1529251.49853738, 1557835.63869696,
  14223.2866511967, 42669.8599535901, 71116.4332559848, 99563.0065583806, 
    128009.579860775, 156456.15316317, 184902.726465566, 213349.29976796, 
    241795.873070355, 270242.446372751, 298689.019675146, 327135.59297754, 
    355582.166279936, 384028.739582331, 412475.312884725, 440921.886187121, 
    469368.459489516, 497815.03279191, 526261.606094305, 554708.179396701, 
    583154.752699096, 611601.326001491, 640047.899303886, 668494.472606281, 
    696941.045908676, 725387.619211071, 753834.192513466, 782280.765815861, 
    810727.339118256, 839173.912420651, 867620.485723046, 896067.059025441, 
    924513.632327836, 952960.205630231, 981406.778932626, 1009853.35223502, 
    1038299.92553742, 1066746.49883981, 1095193.07214221, 1123639.6454446, 
    1152086.218747, 1180532.79204939, 1208979.36535179, 1237425.93865418, 
    1265872.51195658, 1294319.08525897, 1322765.65856137, 1351212.23186376, 
    1379658.80516616, 1408105.37846855, 1436551.95177095, 1464998.52507334, 
    1493445.09837574, 1521891.67167813, 1550338.24498053,
  14154.0218180696, 42462.0654542088, 70770.1090903492, 99078.1527264907, 
    127386.196362631, 155694.239998772, 184002.283634913, 212310.327271054, 
    240618.370907194, 268926.414543335, 297234.458179476, 325542.501815616, 
    353850.545451758, 382158.589087898, 410466.632724039, 438774.67636018, 
    467082.719996321, 495390.76363246, 523698.807268601, 552006.850904743, 
    580314.894540884, 608622.938177024, 636930.981813165, 665239.025449306, 
    693547.069085447, 721855.112721588, 750163.156357729, 778471.199993869, 
    806779.24363001, 835087.287266151, 863395.330902291, 891703.374538432, 
    920011.418174573, 948319.461810714, 976627.505446855, 1004935.549083, 
    1033243.59271914, 1061551.63635528, 1089859.67999142, 1118167.72362756, 
    1146475.7672637, 1174783.81089984, 1203091.85453598, 1231399.89817212, 
    1259707.94180826, 1288015.9854444, 1316324.02908054, 1344632.07271669, 
    1372940.11635283, 1401248.15998897, 1429556.20362511, 1457864.24726125, 
    1486172.29089739, 1514480.33453353, 1542788.37816967,
  14084.2779247904, 42252.8337743712, 70421.3896239533, 98589.9454735365, 
    126758.501323119, 154927.057172701, 183095.613022284, 211264.168871866, 
    239432.724721448, 267601.280571031, 295769.836420613, 323938.392270195, 
    352106.948119778, 380275.50396936, 408444.059818942, 436612.615668525, 
    464781.171518108, 492949.727367689, 521118.283217272, 549286.839066855, 
    577455.394916437, 605623.95076602, 633792.506615602, 661961.062465185, 
    690129.618314767, 718298.174164349, 746466.730013932, 774635.285863514, 
    802803.841713097, 830972.397562679, 859140.953412261, 887309.509261844, 
    915478.065111426, 943646.620961009, 971815.176810591, 999983.732660174, 
    1028152.28850976, 1056320.84435934, 1084489.40020892, 1112657.9560585, 
    1140826.51190809, 1168995.06775767, 1197163.62360725, 1225332.17945683, 
    1253500.73530642, 1281669.291156, 1309837.84700558, 1338006.40285516, 
    1366174.95870475, 1394343.51455433, 1422512.07040391, 1450680.62625349, 
    1478849.18210307, 1507017.73795266, 1535186.29380224,
  14014.0573319573, 42042.1719958718, 70070.2866597876, 98098.4013237046, 
    126126.51598762, 154154.630651536, 182182.745315453, 210210.859979369, 
    238238.974643285, 266267.089307202, 294295.203971117, 322323.318635033, 
    350351.43329895, 378379.547962866, 406407.662626781, 434435.777290698, 
    462463.891954614, 490492.006618529, 518520.121282446, 546548.235946363, 
    574576.350610279, 602604.465274195, 630632.579938111, 658660.694602027, 
    686688.809265943, 714716.92392986, 742745.038593776, 770773.153257692, 
    798801.267921608, 826829.382585524, 854857.49724944, 882885.611913356, 
    910913.726577273, 938941.841241189, 966969.955905105, 994998.070569021, 
    1023026.18523294, 1051054.29989685, 1079082.41456077, 1107110.52922469, 
    1135138.6438886, 1163166.75855252, 1191194.87321643, 1219222.98788035, 
    1247251.10254427, 1275279.21720818, 1303307.3318721, 1331335.44653601, 
    1359363.56119993, 1387391.67586385, 1415419.79052776, 1443447.90519168, 
    1471476.01985559, 1499504.13451951, 1527532.24918343,
  13943.3624163025, 41830.0872489076, 69716.8120815138, 97603.5369141213, 
    125490.261746728, 153376.986579334, 181263.711411941, 209150.436244547, 
    237037.161077154, 264923.885909761, 292810.610742367, 320697.335574974, 
    348584.060407581, 376470.785240187, 404357.510072794, 432244.234905401, 
    460130.959738007, 488017.684570613, 515904.40940322, 543791.134235827, 
    571677.859068434, 599564.58390104, 627451.308733647, 655338.033566254, 
    683224.75839886, 711111.483231467, 738998.208064074, 766884.93289668, 
    794771.657729287, 822658.382561894, 850545.1073945, 878431.832227107, 
    906318.557059714, 934205.28189232, 962092.006724927, 989978.731557534, 
    1017865.45639014, 1045752.18122275, 1073638.90605535, 1101525.63088796, 
    1129412.35572057, 1157299.08055317, 1185185.80538578, 1213072.53021839, 
    1240959.25505099, 1268845.9798836, 1296732.70471621, 1324619.42954881, 
    1352506.15438142, 1380392.87921403, 1408279.60404663, 1436166.32887924, 
    1464053.05371185, 1491939.77854445, 1519826.50337706,
  13872.1955706123, 41616.5867118368, 69360.9778530625, 97105.3689942895, 
    124849.760135515, 152594.151276741, 180338.542417968, 208082.933559194, 
    235827.324700419, 263571.715841646, 291316.106982872, 319060.498124098, 
    346804.889265325, 374549.28040655, 402293.671547776, 430038.062689003, 
    457782.453830229, 485526.844971454, 513271.23611268, 541015.627253907, 
    568760.018395133, 596504.409536359, 624248.800677586, 651993.191818812, 
    679737.582960038, 707481.974101264, 735226.36524249, 762970.756383716, 
    790715.147524942, 818459.538666169, 846203.929807395, 873948.320948621, 
    901692.712089847, 929437.103231073, 957181.494372299, 984925.885513526, 
    1012670.27665475, 1040414.66779598, 1068159.0589372, 1095903.45007843, 
    1123647.84121966, 1151392.23236088, 1179136.62350211, 1206881.01464333, 
    1234625.40578456, 1262369.79692579, 1290114.18806701, 1317858.57920824, 
    1345602.97034946, 1373347.36149069, 1401091.75263192, 1428836.14377314, 
    1456580.53491437, 1484324.92605559, 1512069.31719682,
  13800.5592036454, 41401.6776109362, 69002.7960182282, 96603.9144255213, 
    124205.032832813, 151806.151240105, 179407.269647398, 207008.38805469, 
    234609.506461982, 262210.624869275, 289811.743276567, 317412.861683859, 
    345013.980091153, 372615.098498445, 400216.216905737, 427817.33531303, 
    455418.453720322, 483019.572127613, 510620.690534906, 538221.808942199, 
    565822.927349491, 593424.045756783, 621025.164164076, 648626.282571369, 
    676227.40097866, 703828.519385953, 731429.637793246, 759030.756200538, 
    786631.87460783, 814232.993015123, 841834.111422415, 869435.229829707, 
    897036.348237, 924637.466644292, 952238.585051585, 979839.703458877, 
    1007440.82186617, 1035041.94027346, 1062643.05868075, 1090244.17708805, 
    1117845.29549534, 1145446.41390263, 1173047.53230992, 1200648.65071722, 
    1228249.76912451, 1255850.8875318, 1283452.00593909, 1311053.12434639, 
    1338654.24275368, 1366255.36116097, 1393856.47956826, 1421457.59797555, 
    1449058.71638285, 1476659.83479014, 1504260.95319743,
  13728.455740052, 41185.3672201561, 68642.2787002614, 96099.1901803678, 
    123556.101660473, 151013.013140578, 178469.924620685, 205926.83610079, 
    233383.747580895, 260840.659061002, 288297.570541107, 315754.482021212, 
    343211.393501319, 370668.304981424, 398125.216461529, 425582.127941635, 
    453039.039421741, 480495.950901845, 507952.862381951, 535409.773862058, 
    562866.685342163, 590323.596822269, 617780.508302375, 645237.41978248, 
    672694.331262586, 700151.242742691, 727608.154222797, 755065.065702903, 
    782521.977183008, 809978.888663114, 837435.800143219, 864892.711623325, 
    892349.623103431, 919806.534583536, 947263.446063642, 974720.357543748, 
    1002177.26902385, 1029634.18050396, 1057091.09198406, 1084548.00346417, 
    1112004.91494428, 1139461.82642438, 1166918.73790449, 1194375.64938459, 
    1221832.5608647, 1249289.4723448, 1276746.38382491, 1304203.29530502, 
    1331660.20678512, 1359117.11826523, 1386574.02974533, 1414030.94122544, 
    1441487.85270554, 1468944.76418565, 1496401.67566575,
  13655.8876202915, 40967.6628608745, 68279.4381014587, 95591.213342044, 
    122902.988582628, 150214.763823212, 177526.539063798, 204838.314304382, 
    232150.089544966, 259461.864785551, 286773.640026136, 314085.41526672, 
    341397.190507305, 368708.965747889, 396020.740988473, 423332.516229059, 
    450644.291469643, 477956.066710226, 505267.841950811, 532579.617191397, 
    559891.392431981, 587203.167672565, 614514.94291315, 641826.718153735, 
    669138.493394319, 696450.268634904, 723762.043875489, 751073.819116073, 
    778385.594356657, 805697.369597242, 833009.144837826, 860320.920078411, 
    887632.695318996, 914944.47055958, 942256.245800165, 969568.02104075, 
    996879.796281334, 1024191.57152192, 1051503.3467625, 1078815.12200309, 
    1106126.89724367, 1133438.67248426, 1160750.44772484, 1188062.22296543, 
    1215373.99820601, 1242685.77344659, 1269997.54868718, 1297309.32392776, 
    1324621.09916835, 1351932.87440893, 1379244.64964952, 1406556.4248901, 
    1433868.20013069, 1461179.97537127, 1488491.75061186,
  13582.8573005497, 40748.571901649, 67914.2865027495, 95080.0011038511, 
    122245.715704952, 149411.430306052, 176577.144907154, 203742.859508254, 
    230908.574109355, 258074.288710456, 285240.003311557, 312405.717912657, 
    339571.432513759, 366737.14711486, 393902.86171596, 421068.576317062, 
    448234.290918162, 475400.005519262, 502565.720120363, 529731.434721465, 
    556897.149322566, 584062.863923666, 611228.578524767, 638394.293125869, 
    665560.007726969, 692725.72232807, 719891.436929171, 747057.151530272, 
    774222.866131373, 801388.580732474, 828554.295333574, 855720.009934675, 
    882885.724535776, 910051.439136877, 937217.153737978, 964382.868339079, 
    991548.582940179, 1018714.29754128, 1045880.01214238, 1073045.72674348, 
    1100211.44134458, 1127377.15594568, 1154542.87054678, 1181708.58514789, 
    1208874.29974899, 1236040.01435009, 1263205.72895119, 1290371.44355229, 
    1317537.15815339, 1344702.87275449, 1371868.58735559, 1399034.30195669, 
    1426200.01655779, 1453365.73115889, 1480531.44575999,
  13509.3672526558, 40528.1017579675, 67546.8362632803, 94565.5707685942, 
    121584.305273907, 148603.03977922, 175621.774284534, 202640.508789847, 
    229659.243295159, 256677.977800473, 283696.712305786, 310715.446811099, 
    337734.181316413, 364752.915821726, 391771.650327039, 418790.384832352, 
    445809.119337665, 472827.853842978, 499846.588348291, 526865.322853605, 
    553884.057358918, 580902.791864231, 607921.526369544, 634940.260874858, 
    661958.995380171, 688977.729885484, 715996.464390797, 743015.19889611, 
    770033.933401424, 797052.667906737, 824071.40241205, 851090.136917363, 
    878108.871422677, 905127.605927989, 932146.340433303, 959165.074938616, 
    986183.809443929, 1013202.54394924, 1040221.27845456, 1067240.01295987, 
    1094258.74746518, 1121277.4819705, 1148296.21647581, 1175314.95098112, 
    1202333.68548643, 1229352.41999175, 1256371.15449706, 1283389.88900237, 
    1310408.62350769, 1337427.358013, 1364446.09251831, 1391464.82702363, 
    1418483.56152894, 1445502.29603425, 1472521.03053957,
  13435.419963999, 40306.2598919971, 67177.0998199963, 94047.9397479966, 
    120918.779675996, 147789.619603995, 174660.459531995, 201531.299459995, 
    228402.139387994, 255272.979315994, 282143.819243993, 309014.659171993, 
    335885.499099993, 362756.339027992, 389627.178955991, 416498.018883992, 
    443368.858811991, 470239.69873999, 497110.538667989, 523981.37859599, 
    550852.218523989, 577723.058451989, 604593.898379989, 631464.738307988, 
    658335.578235988, 685206.418163987, 712077.258091987, 738948.098019986, 
    765818.937947986, 792689.777875986, 819560.617803985, 846431.457731985, 
    873302.297659985, 900173.137587984, 927043.977515984, 953914.817443984, 
    980785.657371983, 1007656.49729998, 1034527.33722798, 1061398.17715598, 
    1088269.01708398, 1115139.85701198, 1142010.69693998, 1168881.53686798, 
    1195752.37679598, 1222623.21672398, 1249494.05665198, 1276364.89657998, 
    1303235.73650798, 1330106.57643598, 1356977.41636398, 1383848.25629198, 
    1410719.09621998, 1437589.93614798, 1464460.77607597,
  13361.0179374439, 40083.0538123317, 66805.0896872206, 93527.1255621107, 
    120249.161437, 146971.197311888, 173693.233186779, 200415.269061667, 
    227137.304936556, 253859.340811446, 280581.376686335, 307303.412561224, 
    334025.448436114, 360747.484311003, 387469.520185892, 414191.556060782, 
    440913.591935671, 467635.62781056, 494357.663685449, 521079.699560339, 
    547801.735435229, 574523.771310118, 601245.807185007, 627967.843059896, 
    654689.878934785, 681411.914809675, 708133.950684565, 734855.986559453, 
    761578.022434343, 788300.058309232, 815022.094184121, 841744.130059011, 
    868466.1659339, 895188.201808789, 921910.237683679, 948632.273558568, 
    975354.309433457, 1002076.34530835, 1028798.38118324, 1055520.41705813, 
    1082242.45293301, 1108964.4888079, 1135686.52468279, 1162408.56055768, 
    1189130.59643257, 1215852.63230746, 1242574.66818235, 1269296.70405724, 
    1296018.73993213, 1322740.77580702, 1349462.81168191, 1376184.8475568, 
    1402906.88343169, 1429628.91930658, 1456350.95518146,
  13286.1636912459, 39858.4910737376, 66430.8184562304, 93003.1458387244, 
    119575.473221217, 146147.80060371, 172720.127986204, 199292.455368697, 
    225864.78275119, 252437.110133684, 279009.437516177, 305581.764898669, 
    332154.092281163, 358726.419663656, 385298.747046149, 411871.074428643, 
    438443.401811136, 465015.729193628, 491588.056576122, 518160.383958616, 
    544732.711341109, 571305.038723602, 597877.366106095, 624449.693488589, 
    651022.020871082, 677594.348253575, 704166.675636068, 730739.003018561, 
    757311.330401055, 783883.657783548, 810455.985166041, 837028.312548534, 
    863600.639931028, 890172.96731352, 916745.294696014, 943317.622078507, 
    969889.949461, 996462.276843494, 1023034.60422599, 1049606.93160848, 
    1076179.25899097, 1102751.58637347, 1129323.91375596, 1155896.24113845, 
    1182468.56852095, 1209040.89590344, 1235613.22328593, 1262185.55066843, 
    1288757.87805092, 1315330.20543341, 1341902.53281591, 1368474.8601984, 
    1395047.18758089, 1421619.51496338, 1448191.84234588,
  13210.859758966, 39632.5792768979, 66054.298794831, 92476.0183127651, 
    118897.737830698, 145319.457348631, 171741.176866565, 198162.896384499, 
    224584.615902432, 251006.335420366, 277428.054938299, 303849.774456232, 
    330271.493974166, 356693.213492099, 383114.933010032, 409536.652527966, 
    435958.372045899, 462380.091563832, 488801.811081766, 515223.5305997, 
    541645.250117633, 568066.969635566, 594488.6891535, 620910.408671434, 
    647332.128189367, 673753.8477073, 700175.567225234, 726597.286743167, 
    753019.006261101, 779440.725779034, 805862.445296967, 832284.164814901, 
    858705.884332835, 885127.603850767, 911549.323368701, 937971.042886635, 
    964392.762404568, 990814.481922501, 1017236.20144043, 1043657.92095837, 
    1070079.6404763, 1096501.35999424, 1122923.07951217, 1149344.7990301, 
    1175766.51854804, 1202188.23806597, 1228609.9575839, 1255031.67710184, 
    1281453.39661977, 1307875.1161377, 1334296.83565564, 1360718.55517357, 
    1387140.2746915, 1413561.99420944, 1439983.71372737,
  13135.1086893851, 39405.3260681553, 65675.5434469267, 91945.7608256992, 
    118215.978204471, 144486.195583242, 170756.412962014, 197026.630340786, 
    223296.847719557, 249567.06509833, 275837.282477101, 302107.499855872, 
    328377.717234645, 354647.934613416, 380918.151992187, 407188.36937096, 
    433458.586749731, 459728.804128502, 485999.021507274, 512269.238886046, 
    538539.456264818, 564809.67364359, 591079.891022362, 617350.108401133, 
    643620.325779905, 669890.543158677, 696160.760537449, 722430.97791622, 
    748701.195294992, 774971.412673764, 801241.630052535, 827511.847431307, 
    853782.064810079, 880052.28218885, 906322.499567622, 932592.716946394, 
    958862.934325165, 985133.151703937, 1011403.36908271, 1037673.58646148, 
    1063943.80384025, 1090214.02121902, 1116484.2385978, 1142754.45597657, 
    1169024.67335534, 1195294.89073411, 1221565.10811288, 1247835.32549165, 
    1274105.54287043, 1300375.7602492, 1326645.97762797, 1352916.19500674, 
    1379186.41238551, 1405456.62976428, 1431726.84714306,
  13058.9130464178, 39176.7391392533, 65294.5652320899, 91412.3913249276, 
    117530.217417764, 143648.043510601, 169765.869603439, 195883.695696275, 
    222001.521789112, 248119.34788195, 274237.173974786, 300355.000067623, 
    326472.82616046, 352590.652253297, 378708.478346134, 404826.304438971, 
    430944.130531808, 457061.956624644, 483179.782717481, 509297.608810319, 
    535415.434903156, 561533.260995993, 587651.08708883, 613768.913181667, 
    639886.739274504, 666004.565367341, 692122.391460178, 718240.217553015, 
    744358.043645852, 770475.869738689, 796593.695831526, 822711.521924363, 
    848829.3480172, 874947.174110037, 901065.000202874, 927182.826295711, 
    953300.652388548, 979418.478481385, 1005536.30457422, 1031654.13066706, 
    1057771.9567599, 1083889.78285273, 1110007.60894557, 1136125.43503841, 
    1162243.26113124, 1188361.08722408, 1214478.91331692, 1240596.73940975, 
    1266714.56550259, 1292832.39159543, 1318950.21768826, 1345068.0437811, 
    1371185.86987394, 1397303.69596678, 1423421.52205961,
  12982.2754090251, 38946.8262270753, 64911.3770451266, 90875.9278631791, 
    116840.47868123, 142805.029499282, 168769.580317334, 194734.131135385, 
    220698.681953437, 246663.232771489, 272627.783589541, 298592.334407592, 
    324556.885225644, 350521.436043695, 376485.986861747, 402450.537679799, 
    428415.088497851, 454379.639315901, 480344.190133953, 506308.740952005, 
    532273.291770057, 558237.842588109, 584202.393406161, 610166.944224212, 
    636131.495042264, 662096.045860316, 688060.596678368, 714025.147496419, 
    739989.698314471, 765954.249132523, 791918.799950574, 817883.350768626, 
    843847.901586678, 869812.452404729, 895777.003222781, 921741.554040833, 
    947706.104858884, 973670.655676936, 999635.206494988, 1025599.75731304, 
    1051564.30813109, 1077528.85894914, 1103493.40976719, 1129457.96058525, 
    1155422.5114033, 1181387.06222135, 1207351.6130394, 1233316.16385745, 
    1259280.7146755, 1285245.26549356, 1311209.81631161, 1337174.36712966, 
    1363138.91794771, 1389103.46876576, 1415068.01958381,
  12905.1983711279, 38715.5951133837, 64525.9918556406, 90336.3885978986, 
    116146.785340155, 141957.182082412, 167767.57882467, 193577.975566927, 
    219388.372309184, 245198.769051442, 271009.165793699, 296819.562535956, 
    322629.959278214, 348440.356020471, 374250.752762728, 400061.149504986, 
    425871.546247242, 451681.942989499, 477492.339731756, 503302.736474014, 
    529113.133216272, 554923.529958528, 580733.926700786, 606544.323443043, 
    632354.7201853, 658165.116927558, 683975.513669815, 709785.910412072, 
    735596.307154329, 761406.703896587, 787217.100638844, 813027.497381101, 
    838837.894123359, 864648.290865615, 890458.687607873, 916269.08435013, 
    942079.481092387, 967889.877834645, 993700.274576902, 1019510.67131916, 
    1045321.06806142, 1071131.46480367, 1096941.86154593, 1122752.25828819, 
    1148562.65503045, 1174373.0517727, 1200183.44851496, 1225993.84525722, 
    1251804.24199947, 1277614.63874173, 1303425.03548399, 1329235.43222625, 
    1355045.8289685, 1380856.22571076, 1406666.62245302,
  12827.6845415185, 38483.0536245555, 64138.4227075937, 89793.7917906329, 
    115449.160873671, 141104.529956709, 166759.899039748, 192415.268122786, 
    218070.637205825, 243726.006288864, 269381.375371902, 295036.74445494, 
    320692.113537979, 346347.482621017, 372002.851704056, 397658.220787095, 
    423313.589870133, 448968.95895317, 474624.328036209, 500279.697119248, 
    525935.066202287, 551590.435285325, 577245.804368364, 602901.173451402, 
    628556.542534441, 654211.911617479, 679867.280700518, 705522.649783556, 
    731178.018866595, 756833.387949633, 782488.757032672, 808144.12611571, 
    833799.495198749, 859454.864281787, 885110.233364826, 910765.602447864, 
    936420.971530903, 962076.340613941, 987731.70969698, 1013387.07878002, 
    1039042.44786306, 1064697.8169461, 1090353.18602913, 1116008.55511217, 
    1141663.92419521, 1167319.29327825, 1192974.66236129, 1218630.03144433, 
    1244285.40052736, 1269940.7696104, 1295596.13869344, 1321251.50777648, 
    1346906.87685952, 1372562.24594256, 1398217.6150256,
  12749.7365437727, 38249.2096313182, 63748.6827188648, 89248.1558064124, 
    114747.628893959, 140247.101981506, 165746.575069053, 191246.0481566, 
    216745.521244146, 242244.994331694, 267744.467419241, 293243.940506787, 
    318743.413594335, 344242.886681881, 369742.359769428, 395241.832856976, 
    420741.305944522, 446240.779032068, 471740.252119615, 497239.725207163, 
    522739.19829471, 548238.671382257, 573738.144469804, 599237.617557351, 
    624737.090644898, 650236.563732445, 675736.036819992, 701235.509907538, 
    726734.982995086, 752234.456082633, 777733.929170179, 803233.402257726, 
    828732.875345273, 854232.34843282, 879731.821520367, 905231.294607914, 
    930730.767695461, 956230.240783008, 981729.713870555, 1007229.1869581, 
    1032728.66004565, 1058228.1331332, 1083727.60622074, 1109227.07930829, 
    1134726.55239584, 1160226.02548338, 1185725.49857093, 1211224.97165848, 
    1236724.44474602, 1262223.91783357, 1287723.39092112, 1313222.86400867, 
    1338722.33709621, 1364221.81018376, 1389721.28327131,
  12671.3570161609, 38014.0710484828, 63356.7850808058, 88699.4991131298, 
    114042.213145453, 139384.927177776, 164727.6412101, 190070.355242423, 
    215413.069274746, 240755.78330707, 266098.497339393, 291441.211371715, 
    316783.92540404, 342126.639436362, 367469.353468685, 392812.06750101, 
    418154.781533332, 443497.495565655, 468840.209597978, 494182.923630302, 
    519525.637662626, 544868.351694949, 570211.065727272, 595553.779759596, 
    620896.493791919, 646239.207824242, 671581.921856566, 696924.635888889, 
    722267.349921212, 747610.063953536, 772952.777985858, 798295.492018182, 
    823638.206050505, 848980.920082828, 874323.634115152, 899666.348147475, 
    925009.062179798, 950351.776212122, 975694.490244445, 1001037.20427677, 
    1026379.91830909, 1051722.63234142, 1077065.34637374, 1102408.06040606, 
    1127750.77443838, 1153093.48847071, 1178436.20250303, 1203778.91653535, 
    1229121.63056768, 1254464.3446, 1279807.05863232, 1305149.77266465, 
    1330492.48669697, 1355835.20072929, 1381177.91476162,
  12592.5486115587, 37777.6458346762, 62962.7430577947, 88147.8402809143, 
    113332.937504033, 138518.034727151, 163703.131950271, 188888.229173389, 
    214073.326396508, 239258.423619627, 264443.520842746, 289628.618065864, 
    314813.715288984, 339998.812512103, 365183.909735221, 390369.006958341, 
    415554.104181459, 440739.201404577, 465924.298627696, 491109.395850816, 
    516294.493073935, 541479.590297053, 566664.687520172, 591849.784743291, 
    617034.88196641, 642219.979189529, 667405.076412648, 692590.173635766, 
    717775.270858885, 742960.368082004, 768145.465305123, 793330.562528242, 
    818515.659751361, 843700.75697448, 868885.854197599, 894070.951420718, 
    919256.048643836, 944441.145866955, 969626.243090074, 994811.340313193, 
    1019996.43753631, 1045181.53475943, 1070366.63198255, 1095551.72920567, 
    1120736.82642879, 1145921.92365191, 1171107.02087503, 1196292.11809814, 
    1221477.21532126, 1246662.31254438, 1271847.4097675, 1297032.50699062, 
    1322217.60421374, 1347402.70143686, 1372587.79865998,
  12513.3139973572, 37539.9419920716, 62566.5699867871, 87593.1979815036, 
    112619.825976219, 137646.453970935, 162673.081965651, 187699.709960367, 
    212726.337955082, 237752.965949799, 262779.593944514, 287806.22193923, 
    312832.849933946, 337859.477928662, 362886.105923377, 387912.733918093, 
    412939.361912809, 437965.989907524, 462992.61790224, 488019.245896956, 
    513045.873891672, 538072.501886388, 563099.129881104, 588125.75787582, 
    613152.385870535, 638179.013865251, 663205.641859967, 688232.269854683, 
    713258.897849399, 738285.525844115, 763312.15383883, 788338.781833546, 
    813365.409828263, 838392.037822978, 863418.665817694, 888445.29381241, 
    913471.921807125, 938498.549801841, 963525.177796558, 988551.805791273, 
    1013578.43378599, 1038605.06178071, 1063631.68977542, 1088658.31777014, 
    1113684.94576485, 1138711.57375957, 1163738.20175428, 1188764.829749, 
    1213791.45774372, 1238818.08573843, 1263844.71373315, 1288871.34172786, 
    1313897.96972258, 1338924.59771729, 1363951.22571201,
  12433.6558553727, 37300.967566118, 62168.2792768644, 87035.5909876119, 
    111902.902698358, 136770.214409105, 161637.526119852, 186504.837830599, 
    211372.149541345, 236239.461252092, 261106.772962839, 285974.084673585, 
    310841.396384333, 335708.708095079, 360576.019805826, 385443.331516573, 
    410310.643227319, 435177.954938065, 460045.266648812, 484912.57835956, 
    509779.890070307, 534647.201781053, 559514.5134918, 584381.825202547, 
    609249.136913294, 634116.44862404, 658983.760334787, 683851.072045534, 
    708718.383756281, 733585.695467028, 758453.007177774, 783320.318888521, 
    808187.630599268, 833054.942310015, 857922.254020761, 882789.565731508, 
    907656.877442255, 932524.189153002, 957391.500863749, 982258.812574495, 
    1007126.12428524, 1031993.43599599, 1056860.74770674, 1081728.05941748, 
    1106595.37112823, 1131462.68283898, 1156329.99454972, 1181197.30626047, 
    1206064.61797122, 1230931.92968196, 1255799.24139271, 1280666.55310346, 
    1305533.8648142, 1330401.17652495, 1355268.4882357 ;

 y_rho =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  37044.2803647582, 37044.2803647582, 37044.2803647582, 37044.2803647582, 
    37044.2803647582, 37044.2803647582, 37044.2803647582, 37044.2803647582, 
    37044.2803647582, 37044.2803647582, 37044.2803647582, 37044.2803647582, 
    37044.2803647582, 37044.2803647582, 37044.2803647582, 37044.2803647582, 
    37044.2803647582, 37044.2803647582, 37044.2803647582, 37044.2803647582, 
    37044.2803647582, 37044.2803647582, 37044.2803647582, 37044.2803647582, 
    37044.2803647582, 37044.2803647582, 37044.2803647582, 37044.2803647582, 
    37044.2803647582, 37044.2803647582, 37044.2803647582, 37044.2803647582, 
    37044.2803647582, 37044.2803647582, 37044.2803647582, 37044.2803647582, 
    37044.2803647582, 37044.2803647582, 37044.2803647582, 37044.2803647582, 
    37044.2803647582, 37044.2803647582, 37044.2803647582, 37044.2803647582, 
    37044.2803647582, 37044.2803647582, 37044.2803647582, 37044.2803647582, 
    37044.2803647582, 37044.2803647582, 37044.2803647582, 37044.2803647582, 
    37044.2803647582, 37044.2803647582, 37044.2803647582, 37044.2803647582,
  74088.5607295167, 74088.5607295167, 74088.5607295167, 74088.5607295167, 
    74088.5607295167, 74088.5607295167, 74088.5607295167, 74088.5607295167, 
    74088.5607295167, 74088.5607295167, 74088.5607295167, 74088.5607295167, 
    74088.5607295167, 74088.5607295167, 74088.5607295167, 74088.5607295167, 
    74088.5607295167, 74088.5607295167, 74088.5607295167, 74088.5607295167, 
    74088.5607295167, 74088.5607295167, 74088.5607295167, 74088.5607295167, 
    74088.5607295167, 74088.5607295167, 74088.5607295167, 74088.5607295167, 
    74088.5607295167, 74088.5607295167, 74088.5607295167, 74088.5607295167, 
    74088.5607295167, 74088.5607295167, 74088.5607295167, 74088.5607295167, 
    74088.5607295167, 74088.5607295167, 74088.5607295167, 74088.5607295167, 
    74088.5607295167, 74088.5607295167, 74088.5607295167, 74088.5607295167, 
    74088.5607295167, 74088.5607295167, 74088.5607295167, 74088.5607295167, 
    74088.5607295167, 74088.5607295167, 74088.5607295167, 74088.5607295167, 
    74088.5607295167, 74088.5607295167, 74088.5607295167, 74088.5607295167,
  111132.841094275, 111132.841094275, 111132.841094275, 111132.841094275, 
    111132.841094275, 111132.841094275, 111132.841094275, 111132.841094275, 
    111132.841094275, 111132.841094275, 111132.841094275, 111132.841094275, 
    111132.841094275, 111132.841094275, 111132.841094275, 111132.841094275, 
    111132.841094275, 111132.841094275, 111132.841094275, 111132.841094275, 
    111132.841094275, 111132.841094275, 111132.841094275, 111132.841094275, 
    111132.841094275, 111132.841094275, 111132.841094275, 111132.841094275, 
    111132.841094275, 111132.841094275, 111132.841094275, 111132.841094275, 
    111132.841094275, 111132.841094275, 111132.841094275, 111132.841094275, 
    111132.841094275, 111132.841094275, 111132.841094275, 111132.841094275, 
    111132.841094275, 111132.841094275, 111132.841094275, 111132.841094275, 
    111132.841094275, 111132.841094275, 111132.841094275, 111132.841094275, 
    111132.841094275, 111132.841094275, 111132.841094275, 111132.841094275, 
    111132.841094275, 111132.841094275, 111132.841094275, 111132.841094275,
  148177.121459033, 148177.121459033, 148177.121459033, 148177.121459033, 
    148177.121459033, 148177.121459033, 148177.121459033, 148177.121459033, 
    148177.121459033, 148177.121459033, 148177.121459033, 148177.121459033, 
    148177.121459033, 148177.121459033, 148177.121459033, 148177.121459033, 
    148177.121459033, 148177.121459033, 148177.121459033, 148177.121459033, 
    148177.121459033, 148177.121459033, 148177.121459033, 148177.121459033, 
    148177.121459033, 148177.121459033, 148177.121459033, 148177.121459033, 
    148177.121459033, 148177.121459033, 148177.121459033, 148177.121459033, 
    148177.121459033, 148177.121459033, 148177.121459033, 148177.121459033, 
    148177.121459033, 148177.121459033, 148177.121459033, 148177.121459033, 
    148177.121459033, 148177.121459033, 148177.121459033, 148177.121459033, 
    148177.121459033, 148177.121459033, 148177.121459033, 148177.121459033, 
    148177.121459033, 148177.121459033, 148177.121459033, 148177.121459033, 
    148177.121459033, 148177.121459033, 148177.121459033, 148177.121459033,
  185221.401823792, 185221.401823792, 185221.401823792, 185221.401823792, 
    185221.401823792, 185221.401823792, 185221.401823792, 185221.401823792, 
    185221.401823792, 185221.401823792, 185221.401823792, 185221.401823792, 
    185221.401823792, 185221.401823792, 185221.401823792, 185221.401823792, 
    185221.401823792, 185221.401823792, 185221.401823792, 185221.401823792, 
    185221.401823792, 185221.401823792, 185221.401823792, 185221.401823792, 
    185221.401823792, 185221.401823792, 185221.401823792, 185221.401823792, 
    185221.401823792, 185221.401823792, 185221.401823792, 185221.401823792, 
    185221.401823792, 185221.401823792, 185221.401823792, 185221.401823792, 
    185221.401823792, 185221.401823792, 185221.401823792, 185221.401823792, 
    185221.401823792, 185221.401823792, 185221.401823792, 185221.401823792, 
    185221.401823792, 185221.401823792, 185221.401823792, 185221.401823792, 
    185221.401823792, 185221.401823792, 185221.401823792, 185221.401823792, 
    185221.401823792, 185221.401823792, 185221.401823792, 185221.401823792,
  222265.682188551, 222265.682188551, 222265.682188551, 222265.682188551, 
    222265.682188551, 222265.682188551, 222265.682188551, 222265.682188551, 
    222265.682188551, 222265.682188551, 222265.682188551, 222265.682188551, 
    222265.682188551, 222265.682188551, 222265.682188551, 222265.682188551, 
    222265.682188551, 222265.682188551, 222265.682188551, 222265.682188551, 
    222265.682188551, 222265.682188551, 222265.682188551, 222265.682188551, 
    222265.682188551, 222265.682188551, 222265.682188551, 222265.682188551, 
    222265.682188551, 222265.682188551, 222265.682188551, 222265.682188551, 
    222265.682188551, 222265.682188551, 222265.682188551, 222265.682188551, 
    222265.682188551, 222265.682188551, 222265.682188551, 222265.682188551, 
    222265.682188551, 222265.682188551, 222265.682188551, 222265.682188551, 
    222265.682188551, 222265.682188551, 222265.682188551, 222265.682188551, 
    222265.682188551, 222265.682188551, 222265.682188551, 222265.682188551, 
    222265.682188551, 222265.682188551, 222265.682188551, 222265.682188551,
  259309.962553309, 259309.962553309, 259309.962553309, 259309.962553309, 
    259309.962553309, 259309.962553309, 259309.962553309, 259309.962553309, 
    259309.962553309, 259309.962553309, 259309.962553309, 259309.962553309, 
    259309.962553309, 259309.962553309, 259309.962553309, 259309.962553309, 
    259309.962553309, 259309.962553309, 259309.962553309, 259309.962553309, 
    259309.962553309, 259309.962553309, 259309.962553309, 259309.962553309, 
    259309.962553309, 259309.962553309, 259309.962553309, 259309.962553309, 
    259309.962553309, 259309.962553309, 259309.962553309, 259309.962553309, 
    259309.962553309, 259309.962553309, 259309.962553309, 259309.962553309, 
    259309.962553309, 259309.962553309, 259309.962553309, 259309.962553309, 
    259309.962553309, 259309.962553309, 259309.962553309, 259309.962553309, 
    259309.962553309, 259309.962553309, 259309.962553309, 259309.962553309, 
    259309.962553309, 259309.962553309, 259309.962553309, 259309.962553309, 
    259309.962553309, 259309.962553309, 259309.962553309, 259309.962553309,
  296354.242918067, 296354.242918067, 296354.242918067, 296354.242918067, 
    296354.242918067, 296354.242918067, 296354.242918067, 296354.242918067, 
    296354.242918067, 296354.242918067, 296354.242918067, 296354.242918067, 
    296354.242918067, 296354.242918067, 296354.242918067, 296354.242918067, 
    296354.242918067, 296354.242918067, 296354.242918067, 296354.242918067, 
    296354.242918067, 296354.242918067, 296354.242918067, 296354.242918067, 
    296354.242918067, 296354.242918067, 296354.242918067, 296354.242918067, 
    296354.242918067, 296354.242918067, 296354.242918067, 296354.242918067, 
    296354.242918067, 296354.242918067, 296354.242918067, 296354.242918067, 
    296354.242918067, 296354.242918067, 296354.242918067, 296354.242918067, 
    296354.242918067, 296354.242918067, 296354.242918067, 296354.242918067, 
    296354.242918067, 296354.242918067, 296354.242918067, 296354.242918067, 
    296354.242918067, 296354.242918067, 296354.242918067, 296354.242918067, 
    296354.242918067, 296354.242918067, 296354.242918067, 296354.242918067,
  333398.523282826, 333398.523282826, 333398.523282826, 333398.523282826, 
    333398.523282826, 333398.523282826, 333398.523282826, 333398.523282826, 
    333398.523282826, 333398.523282826, 333398.523282826, 333398.523282826, 
    333398.523282826, 333398.523282826, 333398.523282826, 333398.523282826, 
    333398.523282826, 333398.523282826, 333398.523282826, 333398.523282826, 
    333398.523282826, 333398.523282826, 333398.523282826, 333398.523282826, 
    333398.523282826, 333398.523282826, 333398.523282826, 333398.523282826, 
    333398.523282826, 333398.523282826, 333398.523282826, 333398.523282826, 
    333398.523282826, 333398.523282826, 333398.523282826, 333398.523282826, 
    333398.523282826, 333398.523282826, 333398.523282826, 333398.523282826, 
    333398.523282826, 333398.523282826, 333398.523282826, 333398.523282826, 
    333398.523282826, 333398.523282826, 333398.523282826, 333398.523282826, 
    333398.523282826, 333398.523282826, 333398.523282826, 333398.523282826, 
    333398.523282826, 333398.523282826, 333398.523282826, 333398.523282826,
  370442.803647584, 370442.803647584, 370442.803647584, 370442.803647584, 
    370442.803647584, 370442.803647584, 370442.803647584, 370442.803647584, 
    370442.803647584, 370442.803647584, 370442.803647584, 370442.803647584, 
    370442.803647584, 370442.803647584, 370442.803647584, 370442.803647584, 
    370442.803647584, 370442.803647584, 370442.803647584, 370442.803647584, 
    370442.803647584, 370442.803647584, 370442.803647584, 370442.803647584, 
    370442.803647584, 370442.803647584, 370442.803647584, 370442.803647584, 
    370442.803647584, 370442.803647584, 370442.803647584, 370442.803647584, 
    370442.803647584, 370442.803647584, 370442.803647584, 370442.803647584, 
    370442.803647584, 370442.803647584, 370442.803647584, 370442.803647584, 
    370442.803647584, 370442.803647584, 370442.803647584, 370442.803647584, 
    370442.803647584, 370442.803647584, 370442.803647584, 370442.803647584, 
    370442.803647584, 370442.803647584, 370442.803647584, 370442.803647584, 
    370442.803647584, 370442.803647584, 370442.803647584, 370442.803647584,
  407487.084012342, 407487.084012342, 407487.084012342, 407487.084012342, 
    407487.084012342, 407487.084012342, 407487.084012342, 407487.084012342, 
    407487.084012342, 407487.084012342, 407487.084012342, 407487.084012342, 
    407487.084012342, 407487.084012342, 407487.084012342, 407487.084012342, 
    407487.084012342, 407487.084012342, 407487.084012342, 407487.084012342, 
    407487.084012342, 407487.084012342, 407487.084012342, 407487.084012342, 
    407487.084012342, 407487.084012342, 407487.084012342, 407487.084012342, 
    407487.084012342, 407487.084012342, 407487.084012342, 407487.084012342, 
    407487.084012342, 407487.084012342, 407487.084012342, 407487.084012342, 
    407487.084012342, 407487.084012342, 407487.084012342, 407487.084012342, 
    407487.084012342, 407487.084012342, 407487.084012342, 407487.084012342, 
    407487.084012342, 407487.084012342, 407487.084012342, 407487.084012342, 
    407487.084012342, 407487.084012342, 407487.084012342, 407487.084012342, 
    407487.084012342, 407487.084012342, 407487.084012342, 407487.084012342,
  444531.364377101, 444531.364377101, 444531.364377101, 444531.364377101, 
    444531.364377101, 444531.364377101, 444531.364377101, 444531.364377101, 
    444531.364377101, 444531.364377101, 444531.364377101, 444531.364377101, 
    444531.364377101, 444531.364377101, 444531.364377101, 444531.364377101, 
    444531.364377101, 444531.364377101, 444531.364377101, 444531.364377101, 
    444531.364377101, 444531.364377101, 444531.364377101, 444531.364377101, 
    444531.364377101, 444531.364377101, 444531.364377101, 444531.364377101, 
    444531.364377101, 444531.364377101, 444531.364377101, 444531.364377101, 
    444531.364377101, 444531.364377101, 444531.364377101, 444531.364377101, 
    444531.364377101, 444531.364377101, 444531.364377101, 444531.364377101, 
    444531.364377101, 444531.364377101, 444531.364377101, 444531.364377101, 
    444531.364377101, 444531.364377101, 444531.364377101, 444531.364377101, 
    444531.364377101, 444531.364377101, 444531.364377101, 444531.364377101, 
    444531.364377101, 444531.364377101, 444531.364377101, 444531.364377101,
  481575.644741859, 481575.644741859, 481575.644741859, 481575.644741859, 
    481575.644741859, 481575.644741859, 481575.644741859, 481575.644741859, 
    481575.644741859, 481575.644741859, 481575.644741859, 481575.644741859, 
    481575.644741859, 481575.644741859, 481575.644741859, 481575.644741859, 
    481575.644741859, 481575.644741859, 481575.644741859, 481575.644741859, 
    481575.644741859, 481575.644741859, 481575.644741859, 481575.644741859, 
    481575.644741859, 481575.644741859, 481575.644741859, 481575.644741859, 
    481575.644741859, 481575.644741859, 481575.644741859, 481575.644741859, 
    481575.644741859, 481575.644741859, 481575.644741859, 481575.644741859, 
    481575.644741859, 481575.644741859, 481575.644741859, 481575.644741859, 
    481575.644741859, 481575.644741859, 481575.644741859, 481575.644741859, 
    481575.644741859, 481575.644741859, 481575.644741859, 481575.644741859, 
    481575.644741859, 481575.644741859, 481575.644741859, 481575.644741859, 
    481575.644741859, 481575.644741859, 481575.644741859, 481575.644741859,
  518619.925106617, 518619.925106617, 518619.925106617, 518619.925106617, 
    518619.925106617, 518619.925106617, 518619.925106617, 518619.925106617, 
    518619.925106617, 518619.925106617, 518619.925106617, 518619.925106617, 
    518619.925106617, 518619.925106617, 518619.925106617, 518619.925106617, 
    518619.925106617, 518619.925106617, 518619.925106617, 518619.925106617, 
    518619.925106617, 518619.925106617, 518619.925106617, 518619.925106617, 
    518619.925106617, 518619.925106617, 518619.925106617, 518619.925106617, 
    518619.925106617, 518619.925106617, 518619.925106617, 518619.925106617, 
    518619.925106617, 518619.925106617, 518619.925106617, 518619.925106617, 
    518619.925106617, 518619.925106617, 518619.925106617, 518619.925106617, 
    518619.925106617, 518619.925106617, 518619.925106617, 518619.925106617, 
    518619.925106617, 518619.925106617, 518619.925106617, 518619.925106617, 
    518619.925106617, 518619.925106617, 518619.925106617, 518619.925106617, 
    518619.925106617, 518619.925106617, 518619.925106617, 518619.925106617,
  555664.205471375, 555664.205471375, 555664.205471375, 555664.205471375, 
    555664.205471375, 555664.205471375, 555664.205471375, 555664.205471375, 
    555664.205471375, 555664.205471375, 555664.205471375, 555664.205471375, 
    555664.205471375, 555664.205471375, 555664.205471375, 555664.205471375, 
    555664.205471375, 555664.205471375, 555664.205471375, 555664.205471375, 
    555664.205471375, 555664.205471375, 555664.205471375, 555664.205471375, 
    555664.205471375, 555664.205471375, 555664.205471375, 555664.205471375, 
    555664.205471375, 555664.205471375, 555664.205471375, 555664.205471375, 
    555664.205471375, 555664.205471375, 555664.205471375, 555664.205471375, 
    555664.205471375, 555664.205471375, 555664.205471375, 555664.205471375, 
    555664.205471375, 555664.205471375, 555664.205471375, 555664.205471375, 
    555664.205471375, 555664.205471375, 555664.205471375, 555664.205471375, 
    555664.205471375, 555664.205471375, 555664.205471375, 555664.205471375, 
    555664.205471375, 555664.205471375, 555664.205471375, 555664.205471375,
  592708.485836134, 592708.485836134, 592708.485836134, 592708.485836134, 
    592708.485836134, 592708.485836134, 592708.485836134, 592708.485836134, 
    592708.485836134, 592708.485836134, 592708.485836134, 592708.485836134, 
    592708.485836134, 592708.485836134, 592708.485836134, 592708.485836134, 
    592708.485836134, 592708.485836134, 592708.485836134, 592708.485836134, 
    592708.485836134, 592708.485836134, 592708.485836134, 592708.485836134, 
    592708.485836134, 592708.485836134, 592708.485836134, 592708.485836134, 
    592708.485836134, 592708.485836134, 592708.485836134, 592708.485836134, 
    592708.485836134, 592708.485836134, 592708.485836134, 592708.485836134, 
    592708.485836134, 592708.485836134, 592708.485836134, 592708.485836134, 
    592708.485836134, 592708.485836134, 592708.485836134, 592708.485836134, 
    592708.485836134, 592708.485836134, 592708.485836134, 592708.485836134, 
    592708.485836134, 592708.485836134, 592708.485836134, 592708.485836134, 
    592708.485836134, 592708.485836134, 592708.485836134, 592708.485836134,
  629752.766200892, 629752.766200892, 629752.766200892, 629752.766200892, 
    629752.766200892, 629752.766200892, 629752.766200892, 629752.766200892, 
    629752.766200892, 629752.766200892, 629752.766200892, 629752.766200892, 
    629752.766200892, 629752.766200892, 629752.766200892, 629752.766200892, 
    629752.766200892, 629752.766200892, 629752.766200892, 629752.766200892, 
    629752.766200892, 629752.766200892, 629752.766200892, 629752.766200892, 
    629752.766200892, 629752.766200892, 629752.766200892, 629752.766200892, 
    629752.766200892, 629752.766200892, 629752.766200892, 629752.766200892, 
    629752.766200892, 629752.766200892, 629752.766200892, 629752.766200892, 
    629752.766200892, 629752.766200892, 629752.766200892, 629752.766200892, 
    629752.766200892, 629752.766200892, 629752.766200892, 629752.766200892, 
    629752.766200892, 629752.766200892, 629752.766200892, 629752.766200892, 
    629752.766200892, 629752.766200892, 629752.766200892, 629752.766200892, 
    629752.766200892, 629752.766200892, 629752.766200892, 629752.766200892,
  666797.04656565, 666797.04656565, 666797.04656565, 666797.04656565, 
    666797.04656565, 666797.04656565, 666797.04656565, 666797.04656565, 
    666797.04656565, 666797.04656565, 666797.04656565, 666797.04656565, 
    666797.04656565, 666797.04656565, 666797.04656565, 666797.04656565, 
    666797.04656565, 666797.04656565, 666797.04656565, 666797.04656565, 
    666797.04656565, 666797.04656565, 666797.04656565, 666797.04656565, 
    666797.04656565, 666797.04656565, 666797.04656565, 666797.04656565, 
    666797.04656565, 666797.04656565, 666797.04656565, 666797.04656565, 
    666797.04656565, 666797.04656565, 666797.04656565, 666797.04656565, 
    666797.04656565, 666797.04656565, 666797.04656565, 666797.04656565, 
    666797.04656565, 666797.04656565, 666797.04656565, 666797.04656565, 
    666797.04656565, 666797.04656565, 666797.04656565, 666797.04656565, 
    666797.04656565, 666797.04656565, 666797.04656565, 666797.04656565, 
    666797.04656565, 666797.04656565, 666797.04656565, 666797.04656565,
  703841.326930409, 703841.326930409, 703841.326930409, 703841.326930409, 
    703841.326930409, 703841.326930409, 703841.326930409, 703841.326930409, 
    703841.326930409, 703841.326930409, 703841.326930409, 703841.326930409, 
    703841.326930409, 703841.326930409, 703841.326930409, 703841.326930409, 
    703841.326930409, 703841.326930409, 703841.326930409, 703841.326930409, 
    703841.326930409, 703841.326930409, 703841.326930409, 703841.326930409, 
    703841.326930409, 703841.326930409, 703841.326930409, 703841.326930409, 
    703841.326930409, 703841.326930409, 703841.326930409, 703841.326930409, 
    703841.326930409, 703841.326930409, 703841.326930409, 703841.326930409, 
    703841.326930409, 703841.326930409, 703841.326930409, 703841.326930409, 
    703841.326930409, 703841.326930409, 703841.326930409, 703841.326930409, 
    703841.326930409, 703841.326930409, 703841.326930409, 703841.326930409, 
    703841.326930409, 703841.326930409, 703841.326930409, 703841.326930409, 
    703841.326930409, 703841.326930409, 703841.326930409, 703841.326930409,
  740885.607295166, 740885.607295166, 740885.607295166, 740885.607295166, 
    740885.607295166, 740885.607295166, 740885.607295166, 740885.607295166, 
    740885.607295166, 740885.607295166, 740885.607295166, 740885.607295166, 
    740885.607295166, 740885.607295166, 740885.607295166, 740885.607295166, 
    740885.607295166, 740885.607295166, 740885.607295166, 740885.607295166, 
    740885.607295166, 740885.607295166, 740885.607295166, 740885.607295166, 
    740885.607295166, 740885.607295166, 740885.607295166, 740885.607295166, 
    740885.607295166, 740885.607295166, 740885.607295166, 740885.607295166, 
    740885.607295166, 740885.607295166, 740885.607295166, 740885.607295166, 
    740885.607295166, 740885.607295166, 740885.607295166, 740885.607295166, 
    740885.607295166, 740885.607295166, 740885.607295166, 740885.607295166, 
    740885.607295166, 740885.607295166, 740885.607295166, 740885.607295166, 
    740885.607295166, 740885.607295166, 740885.607295166, 740885.607295166, 
    740885.607295166, 740885.607295166, 740885.607295166, 740885.607295166,
  777929.887659925, 777929.887659925, 777929.887659925, 777929.887659925, 
    777929.887659925, 777929.887659925, 777929.887659925, 777929.887659925, 
    777929.887659925, 777929.887659925, 777929.887659925, 777929.887659925, 
    777929.887659925, 777929.887659925, 777929.887659925, 777929.887659925, 
    777929.887659925, 777929.887659925, 777929.887659925, 777929.887659925, 
    777929.887659925, 777929.887659925, 777929.887659925, 777929.887659925, 
    777929.887659925, 777929.887659925, 777929.887659925, 777929.887659925, 
    777929.887659925, 777929.887659925, 777929.887659925, 777929.887659925, 
    777929.887659925, 777929.887659925, 777929.887659925, 777929.887659925, 
    777929.887659925, 777929.887659925, 777929.887659925, 777929.887659925, 
    777929.887659925, 777929.887659925, 777929.887659925, 777929.887659925, 
    777929.887659925, 777929.887659925, 777929.887659925, 777929.887659925, 
    777929.887659925, 777929.887659925, 777929.887659925, 777929.887659925, 
    777929.887659925, 777929.887659925, 777929.887659925, 777929.887659925,
  814974.168024684, 814974.168024684, 814974.168024684, 814974.168024684, 
    814974.168024684, 814974.168024684, 814974.168024684, 814974.168024684, 
    814974.168024684, 814974.168024684, 814974.168024684, 814974.168024684, 
    814974.168024684, 814974.168024684, 814974.168024684, 814974.168024684, 
    814974.168024684, 814974.168024684, 814974.168024684, 814974.168024684, 
    814974.168024684, 814974.168024684, 814974.168024684, 814974.168024684, 
    814974.168024684, 814974.168024684, 814974.168024684, 814974.168024684, 
    814974.168024684, 814974.168024684, 814974.168024684, 814974.168024684, 
    814974.168024684, 814974.168024684, 814974.168024684, 814974.168024684, 
    814974.168024684, 814974.168024684, 814974.168024684, 814974.168024684, 
    814974.168024684, 814974.168024684, 814974.168024684, 814974.168024684, 
    814974.168024684, 814974.168024684, 814974.168024684, 814974.168024684, 
    814974.168024684, 814974.168024684, 814974.168024684, 814974.168024684, 
    814974.168024684, 814974.168024684, 814974.168024684, 814974.168024684,
  852018.448389441, 852018.448389441, 852018.448389441, 852018.448389441, 
    852018.448389441, 852018.448389441, 852018.448389441, 852018.448389441, 
    852018.448389441, 852018.448389441, 852018.448389441, 852018.448389441, 
    852018.448389441, 852018.448389441, 852018.448389441, 852018.448389441, 
    852018.448389441, 852018.448389441, 852018.448389441, 852018.448389441, 
    852018.448389441, 852018.448389441, 852018.448389441, 852018.448389441, 
    852018.448389441, 852018.448389441, 852018.448389441, 852018.448389441, 
    852018.448389441, 852018.448389441, 852018.448389441, 852018.448389441, 
    852018.448389441, 852018.448389441, 852018.448389441, 852018.448389441, 
    852018.448389441, 852018.448389441, 852018.448389441, 852018.448389441, 
    852018.448389441, 852018.448389441, 852018.448389441, 852018.448389441, 
    852018.448389441, 852018.448389441, 852018.448389441, 852018.448389441, 
    852018.448389441, 852018.448389441, 852018.448389441, 852018.448389441, 
    852018.448389441, 852018.448389441, 852018.448389441, 852018.448389441,
  889062.7287542, 889062.7287542, 889062.7287542, 889062.7287542, 
    889062.7287542, 889062.7287542, 889062.7287542, 889062.7287542, 
    889062.7287542, 889062.7287542, 889062.7287542, 889062.7287542, 
    889062.7287542, 889062.7287542, 889062.7287542, 889062.7287542, 
    889062.7287542, 889062.7287542, 889062.7287542, 889062.7287542, 
    889062.7287542, 889062.7287542, 889062.7287542, 889062.7287542, 
    889062.7287542, 889062.7287542, 889062.7287542, 889062.7287542, 
    889062.7287542, 889062.7287542, 889062.7287542, 889062.7287542, 
    889062.7287542, 889062.7287542, 889062.7287542, 889062.7287542, 
    889062.7287542, 889062.7287542, 889062.7287542, 889062.7287542, 
    889062.7287542, 889062.7287542, 889062.7287542, 889062.7287542, 
    889062.7287542, 889062.7287542, 889062.7287542, 889062.7287542, 
    889062.7287542, 889062.7287542, 889062.7287542, 889062.7287542, 
    889062.7287542, 889062.7287542, 889062.7287542, 889062.7287542,
  926107.009118958, 926107.009118958, 926107.009118958, 926107.009118958, 
    926107.009118958, 926107.009118958, 926107.009118958, 926107.009118958, 
    926107.009118958, 926107.009118958, 926107.009118958, 926107.009118958, 
    926107.009118958, 926107.009118958, 926107.009118958, 926107.009118958, 
    926107.009118958, 926107.009118958, 926107.009118958, 926107.009118958, 
    926107.009118958, 926107.009118958, 926107.009118958, 926107.009118958, 
    926107.009118958, 926107.009118958, 926107.009118958, 926107.009118958, 
    926107.009118958, 926107.009118958, 926107.009118958, 926107.009118958, 
    926107.009118958, 926107.009118958, 926107.009118958, 926107.009118958, 
    926107.009118958, 926107.009118958, 926107.009118958, 926107.009118958, 
    926107.009118958, 926107.009118958, 926107.009118958, 926107.009118958, 
    926107.009118958, 926107.009118958, 926107.009118958, 926107.009118958, 
    926107.009118958, 926107.009118958, 926107.009118958, 926107.009118958, 
    926107.009118958, 926107.009118958, 926107.009118958, 926107.009118958,
  963151.289483716, 963151.289483716, 963151.289483716, 963151.289483716, 
    963151.289483716, 963151.289483716, 963151.289483716, 963151.289483716, 
    963151.289483716, 963151.289483716, 963151.289483716, 963151.289483716, 
    963151.289483716, 963151.289483716, 963151.289483716, 963151.289483716, 
    963151.289483716, 963151.289483716, 963151.289483716, 963151.289483716, 
    963151.289483716, 963151.289483716, 963151.289483716, 963151.289483716, 
    963151.289483716, 963151.289483716, 963151.289483716, 963151.289483716, 
    963151.289483716, 963151.289483716, 963151.289483716, 963151.289483716, 
    963151.289483716, 963151.289483716, 963151.289483716, 963151.289483716, 
    963151.289483716, 963151.289483716, 963151.289483716, 963151.289483716, 
    963151.289483716, 963151.289483716, 963151.289483716, 963151.289483716, 
    963151.289483716, 963151.289483716, 963151.289483716, 963151.289483716, 
    963151.289483716, 963151.289483716, 963151.289483716, 963151.289483716, 
    963151.289483716, 963151.289483716, 963151.289483716, 963151.289483716,
  1000195.56984848, 1000195.56984848, 1000195.56984848, 1000195.56984848, 
    1000195.56984848, 1000195.56984848, 1000195.56984848, 1000195.56984848, 
    1000195.56984848, 1000195.56984848, 1000195.56984848, 1000195.56984848, 
    1000195.56984848, 1000195.56984848, 1000195.56984848, 1000195.56984848, 
    1000195.56984848, 1000195.56984848, 1000195.56984848, 1000195.56984848, 
    1000195.56984848, 1000195.56984848, 1000195.56984848, 1000195.56984848, 
    1000195.56984848, 1000195.56984848, 1000195.56984848, 1000195.56984848, 
    1000195.56984848, 1000195.56984848, 1000195.56984848, 1000195.56984848, 
    1000195.56984848, 1000195.56984848, 1000195.56984848, 1000195.56984848, 
    1000195.56984848, 1000195.56984848, 1000195.56984848, 1000195.56984848, 
    1000195.56984848, 1000195.56984848, 1000195.56984848, 1000195.56984848, 
    1000195.56984848, 1000195.56984848, 1000195.56984848, 1000195.56984848, 
    1000195.56984848, 1000195.56984848, 1000195.56984848, 1000195.56984848, 
    1000195.56984848, 1000195.56984848, 1000195.56984848, 1000195.56984848,
  1037239.85021323, 1037239.85021323, 1037239.85021323, 1037239.85021323, 
    1037239.85021323, 1037239.85021323, 1037239.85021323, 1037239.85021323, 
    1037239.85021323, 1037239.85021323, 1037239.85021323, 1037239.85021323, 
    1037239.85021323, 1037239.85021323, 1037239.85021323, 1037239.85021323, 
    1037239.85021323, 1037239.85021323, 1037239.85021323, 1037239.85021323, 
    1037239.85021323, 1037239.85021323, 1037239.85021323, 1037239.85021323, 
    1037239.85021323, 1037239.85021323, 1037239.85021323, 1037239.85021323, 
    1037239.85021323, 1037239.85021323, 1037239.85021323, 1037239.85021323, 
    1037239.85021323, 1037239.85021323, 1037239.85021323, 1037239.85021323, 
    1037239.85021323, 1037239.85021323, 1037239.85021323, 1037239.85021323, 
    1037239.85021323, 1037239.85021323, 1037239.85021323, 1037239.85021323, 
    1037239.85021323, 1037239.85021323, 1037239.85021323, 1037239.85021323, 
    1037239.85021323, 1037239.85021323, 1037239.85021323, 1037239.85021323, 
    1037239.85021323, 1037239.85021323, 1037239.85021323, 1037239.85021323,
  1074284.13057799, 1074284.13057799, 1074284.13057799, 1074284.13057799, 
    1074284.13057799, 1074284.13057799, 1074284.13057799, 1074284.13057799, 
    1074284.13057799, 1074284.13057799, 1074284.13057799, 1074284.13057799, 
    1074284.13057799, 1074284.13057799, 1074284.13057799, 1074284.13057799, 
    1074284.13057799, 1074284.13057799, 1074284.13057799, 1074284.13057799, 
    1074284.13057799, 1074284.13057799, 1074284.13057799, 1074284.13057799, 
    1074284.13057799, 1074284.13057799, 1074284.13057799, 1074284.13057799, 
    1074284.13057799, 1074284.13057799, 1074284.13057799, 1074284.13057799, 
    1074284.13057799, 1074284.13057799, 1074284.13057799, 1074284.13057799, 
    1074284.13057799, 1074284.13057799, 1074284.13057799, 1074284.13057799, 
    1074284.13057799, 1074284.13057799, 1074284.13057799, 1074284.13057799, 
    1074284.13057799, 1074284.13057799, 1074284.13057799, 1074284.13057799, 
    1074284.13057799, 1074284.13057799, 1074284.13057799, 1074284.13057799, 
    1074284.13057799, 1074284.13057799, 1074284.13057799, 1074284.13057799,
  1111328.41094275, 1111328.41094275, 1111328.41094275, 1111328.41094275, 
    1111328.41094275, 1111328.41094275, 1111328.41094275, 1111328.41094275, 
    1111328.41094275, 1111328.41094275, 1111328.41094275, 1111328.41094275, 
    1111328.41094275, 1111328.41094275, 1111328.41094275, 1111328.41094275, 
    1111328.41094275, 1111328.41094275, 1111328.41094275, 1111328.41094275, 
    1111328.41094275, 1111328.41094275, 1111328.41094275, 1111328.41094275, 
    1111328.41094275, 1111328.41094275, 1111328.41094275, 1111328.41094275, 
    1111328.41094275, 1111328.41094275, 1111328.41094275, 1111328.41094275, 
    1111328.41094275, 1111328.41094275, 1111328.41094275, 1111328.41094275, 
    1111328.41094275, 1111328.41094275, 1111328.41094275, 1111328.41094275, 
    1111328.41094275, 1111328.41094275, 1111328.41094275, 1111328.41094275, 
    1111328.41094275, 1111328.41094275, 1111328.41094275, 1111328.41094275, 
    1111328.41094275, 1111328.41094275, 1111328.41094275, 1111328.41094275, 
    1111328.41094275, 1111328.41094275, 1111328.41094275, 1111328.41094275,
  1148372.69130751, 1148372.69130751, 1148372.69130751, 1148372.69130751, 
    1148372.69130751, 1148372.69130751, 1148372.69130751, 1148372.69130751, 
    1148372.69130751, 1148372.69130751, 1148372.69130751, 1148372.69130751, 
    1148372.69130751, 1148372.69130751, 1148372.69130751, 1148372.69130751, 
    1148372.69130751, 1148372.69130751, 1148372.69130751, 1148372.69130751, 
    1148372.69130751, 1148372.69130751, 1148372.69130751, 1148372.69130751, 
    1148372.69130751, 1148372.69130751, 1148372.69130751, 1148372.69130751, 
    1148372.69130751, 1148372.69130751, 1148372.69130751, 1148372.69130751, 
    1148372.69130751, 1148372.69130751, 1148372.69130751, 1148372.69130751, 
    1148372.69130751, 1148372.69130751, 1148372.69130751, 1148372.69130751, 
    1148372.69130751, 1148372.69130751, 1148372.69130751, 1148372.69130751, 
    1148372.69130751, 1148372.69130751, 1148372.69130751, 1148372.69130751, 
    1148372.69130751, 1148372.69130751, 1148372.69130751, 1148372.69130751, 
    1148372.69130751, 1148372.69130751, 1148372.69130751, 1148372.69130751,
  1185416.97167227, 1185416.97167227, 1185416.97167227, 1185416.97167227, 
    1185416.97167227, 1185416.97167227, 1185416.97167227, 1185416.97167227, 
    1185416.97167227, 1185416.97167227, 1185416.97167227, 1185416.97167227, 
    1185416.97167227, 1185416.97167227, 1185416.97167227, 1185416.97167227, 
    1185416.97167227, 1185416.97167227, 1185416.97167227, 1185416.97167227, 
    1185416.97167227, 1185416.97167227, 1185416.97167227, 1185416.97167227, 
    1185416.97167227, 1185416.97167227, 1185416.97167227, 1185416.97167227, 
    1185416.97167227, 1185416.97167227, 1185416.97167227, 1185416.97167227, 
    1185416.97167227, 1185416.97167227, 1185416.97167227, 1185416.97167227, 
    1185416.97167227, 1185416.97167227, 1185416.97167227, 1185416.97167227, 
    1185416.97167227, 1185416.97167227, 1185416.97167227, 1185416.97167227, 
    1185416.97167227, 1185416.97167227, 1185416.97167227, 1185416.97167227, 
    1185416.97167227, 1185416.97167227, 1185416.97167227, 1185416.97167227, 
    1185416.97167227, 1185416.97167227, 1185416.97167227, 1185416.97167227,
  1222461.25203703, 1222461.25203703, 1222461.25203703, 1222461.25203703, 
    1222461.25203703, 1222461.25203703, 1222461.25203703, 1222461.25203703, 
    1222461.25203703, 1222461.25203703, 1222461.25203703, 1222461.25203703, 
    1222461.25203703, 1222461.25203703, 1222461.25203703, 1222461.25203703, 
    1222461.25203703, 1222461.25203703, 1222461.25203703, 1222461.25203703, 
    1222461.25203703, 1222461.25203703, 1222461.25203703, 1222461.25203703, 
    1222461.25203703, 1222461.25203703, 1222461.25203703, 1222461.25203703, 
    1222461.25203703, 1222461.25203703, 1222461.25203703, 1222461.25203703, 
    1222461.25203703, 1222461.25203703, 1222461.25203703, 1222461.25203703, 
    1222461.25203703, 1222461.25203703, 1222461.25203703, 1222461.25203703, 
    1222461.25203703, 1222461.25203703, 1222461.25203703, 1222461.25203703, 
    1222461.25203703, 1222461.25203703, 1222461.25203703, 1222461.25203703, 
    1222461.25203703, 1222461.25203703, 1222461.25203703, 1222461.25203703, 
    1222461.25203703, 1222461.25203703, 1222461.25203703, 1222461.25203703,
  1259505.53240178, 1259505.53240178, 1259505.53240178, 1259505.53240178, 
    1259505.53240178, 1259505.53240178, 1259505.53240178, 1259505.53240178, 
    1259505.53240178, 1259505.53240178, 1259505.53240178, 1259505.53240178, 
    1259505.53240178, 1259505.53240178, 1259505.53240178, 1259505.53240178, 
    1259505.53240178, 1259505.53240178, 1259505.53240178, 1259505.53240178, 
    1259505.53240178, 1259505.53240178, 1259505.53240178, 1259505.53240178, 
    1259505.53240178, 1259505.53240178, 1259505.53240178, 1259505.53240178, 
    1259505.53240178, 1259505.53240178, 1259505.53240178, 1259505.53240178, 
    1259505.53240178, 1259505.53240178, 1259505.53240178, 1259505.53240178, 
    1259505.53240178, 1259505.53240178, 1259505.53240178, 1259505.53240178, 
    1259505.53240178, 1259505.53240178, 1259505.53240178, 1259505.53240178, 
    1259505.53240178, 1259505.53240178, 1259505.53240178, 1259505.53240178, 
    1259505.53240178, 1259505.53240178, 1259505.53240178, 1259505.53240178, 
    1259505.53240178, 1259505.53240178, 1259505.53240178, 1259505.53240178,
  1296549.81276654, 1296549.81276654, 1296549.81276654, 1296549.81276654, 
    1296549.81276654, 1296549.81276654, 1296549.81276654, 1296549.81276654, 
    1296549.81276654, 1296549.81276654, 1296549.81276654, 1296549.81276654, 
    1296549.81276654, 1296549.81276654, 1296549.81276654, 1296549.81276654, 
    1296549.81276654, 1296549.81276654, 1296549.81276654, 1296549.81276654, 
    1296549.81276654, 1296549.81276654, 1296549.81276654, 1296549.81276654, 
    1296549.81276654, 1296549.81276654, 1296549.81276654, 1296549.81276654, 
    1296549.81276654, 1296549.81276654, 1296549.81276654, 1296549.81276654, 
    1296549.81276654, 1296549.81276654, 1296549.81276654, 1296549.81276654, 
    1296549.81276654, 1296549.81276654, 1296549.81276654, 1296549.81276654, 
    1296549.81276654, 1296549.81276654, 1296549.81276654, 1296549.81276654, 
    1296549.81276654, 1296549.81276654, 1296549.81276654, 1296549.81276654, 
    1296549.81276654, 1296549.81276654, 1296549.81276654, 1296549.81276654, 
    1296549.81276654, 1296549.81276654, 1296549.81276654, 1296549.81276654,
  1333594.0931313, 1333594.0931313, 1333594.0931313, 1333594.0931313, 
    1333594.0931313, 1333594.0931313, 1333594.0931313, 1333594.0931313, 
    1333594.0931313, 1333594.0931313, 1333594.0931313, 1333594.0931313, 
    1333594.0931313, 1333594.0931313, 1333594.0931313, 1333594.0931313, 
    1333594.0931313, 1333594.0931313, 1333594.0931313, 1333594.0931313, 
    1333594.0931313, 1333594.0931313, 1333594.0931313, 1333594.0931313, 
    1333594.0931313, 1333594.0931313, 1333594.0931313, 1333594.0931313, 
    1333594.0931313, 1333594.0931313, 1333594.0931313, 1333594.0931313, 
    1333594.0931313, 1333594.0931313, 1333594.0931313, 1333594.0931313, 
    1333594.0931313, 1333594.0931313, 1333594.0931313, 1333594.0931313, 
    1333594.0931313, 1333594.0931313, 1333594.0931313, 1333594.0931313, 
    1333594.0931313, 1333594.0931313, 1333594.0931313, 1333594.0931313, 
    1333594.0931313, 1333594.0931313, 1333594.0931313, 1333594.0931313, 
    1333594.0931313, 1333594.0931313, 1333594.0931313, 1333594.0931313,
  1370638.37349606, 1370638.37349606, 1370638.37349606, 1370638.37349606, 
    1370638.37349606, 1370638.37349606, 1370638.37349606, 1370638.37349606, 
    1370638.37349606, 1370638.37349606, 1370638.37349606, 1370638.37349606, 
    1370638.37349606, 1370638.37349606, 1370638.37349606, 1370638.37349606, 
    1370638.37349606, 1370638.37349606, 1370638.37349606, 1370638.37349606, 
    1370638.37349606, 1370638.37349606, 1370638.37349606, 1370638.37349606, 
    1370638.37349606, 1370638.37349606, 1370638.37349606, 1370638.37349606, 
    1370638.37349606, 1370638.37349606, 1370638.37349606, 1370638.37349606, 
    1370638.37349606, 1370638.37349606, 1370638.37349606, 1370638.37349606, 
    1370638.37349606, 1370638.37349606, 1370638.37349606, 1370638.37349606, 
    1370638.37349606, 1370638.37349606, 1370638.37349606, 1370638.37349606, 
    1370638.37349606, 1370638.37349606, 1370638.37349606, 1370638.37349606, 
    1370638.37349606, 1370638.37349606, 1370638.37349606, 1370638.37349606, 
    1370638.37349606, 1370638.37349606, 1370638.37349606, 1370638.37349606,
  1407682.65386082, 1407682.65386082, 1407682.65386082, 1407682.65386082, 
    1407682.65386082, 1407682.65386082, 1407682.65386082, 1407682.65386082, 
    1407682.65386082, 1407682.65386082, 1407682.65386082, 1407682.65386082, 
    1407682.65386082, 1407682.65386082, 1407682.65386082, 1407682.65386082, 
    1407682.65386082, 1407682.65386082, 1407682.65386082, 1407682.65386082, 
    1407682.65386082, 1407682.65386082, 1407682.65386082, 1407682.65386082, 
    1407682.65386082, 1407682.65386082, 1407682.65386082, 1407682.65386082, 
    1407682.65386082, 1407682.65386082, 1407682.65386082, 1407682.65386082, 
    1407682.65386082, 1407682.65386082, 1407682.65386082, 1407682.65386082, 
    1407682.65386082, 1407682.65386082, 1407682.65386082, 1407682.65386082, 
    1407682.65386082, 1407682.65386082, 1407682.65386082, 1407682.65386082, 
    1407682.65386082, 1407682.65386082, 1407682.65386082, 1407682.65386082, 
    1407682.65386082, 1407682.65386082, 1407682.65386082, 1407682.65386082, 
    1407682.65386082, 1407682.65386082, 1407682.65386082, 1407682.65386082,
  1444726.93422558, 1444726.93422558, 1444726.93422558, 1444726.93422558, 
    1444726.93422558, 1444726.93422558, 1444726.93422558, 1444726.93422558, 
    1444726.93422558, 1444726.93422558, 1444726.93422558, 1444726.93422558, 
    1444726.93422558, 1444726.93422558, 1444726.93422558, 1444726.93422558, 
    1444726.93422558, 1444726.93422558, 1444726.93422558, 1444726.93422558, 
    1444726.93422558, 1444726.93422558, 1444726.93422558, 1444726.93422558, 
    1444726.93422558, 1444726.93422558, 1444726.93422558, 1444726.93422558, 
    1444726.93422558, 1444726.93422558, 1444726.93422558, 1444726.93422558, 
    1444726.93422558, 1444726.93422558, 1444726.93422558, 1444726.93422558, 
    1444726.93422558, 1444726.93422558, 1444726.93422558, 1444726.93422558, 
    1444726.93422558, 1444726.93422558, 1444726.93422558, 1444726.93422558, 
    1444726.93422558, 1444726.93422558, 1444726.93422558, 1444726.93422558, 
    1444726.93422558, 1444726.93422558, 1444726.93422558, 1444726.93422558, 
    1444726.93422558, 1444726.93422558, 1444726.93422558, 1444726.93422558,
  1481771.21459033, 1481771.21459033, 1481771.21459033, 1481771.21459033, 
    1481771.21459033, 1481771.21459033, 1481771.21459033, 1481771.21459033, 
    1481771.21459033, 1481771.21459033, 1481771.21459033, 1481771.21459033, 
    1481771.21459033, 1481771.21459033, 1481771.21459033, 1481771.21459033, 
    1481771.21459033, 1481771.21459033, 1481771.21459033, 1481771.21459033, 
    1481771.21459033, 1481771.21459033, 1481771.21459033, 1481771.21459033, 
    1481771.21459033, 1481771.21459033, 1481771.21459033, 1481771.21459033, 
    1481771.21459033, 1481771.21459033, 1481771.21459033, 1481771.21459033, 
    1481771.21459033, 1481771.21459033, 1481771.21459033, 1481771.21459033, 
    1481771.21459033, 1481771.21459033, 1481771.21459033, 1481771.21459033, 
    1481771.21459033, 1481771.21459033, 1481771.21459033, 1481771.21459033, 
    1481771.21459033, 1481771.21459033, 1481771.21459033, 1481771.21459033, 
    1481771.21459033, 1481771.21459033, 1481771.21459033, 1481771.21459033, 
    1481771.21459033, 1481771.21459033, 1481771.21459033, 1481771.21459033,
  1518815.49495509, 1518815.49495509, 1518815.49495509, 1518815.49495509, 
    1518815.49495509, 1518815.49495509, 1518815.49495509, 1518815.49495509, 
    1518815.49495509, 1518815.49495509, 1518815.49495509, 1518815.49495509, 
    1518815.49495509, 1518815.49495509, 1518815.49495509, 1518815.49495509, 
    1518815.49495509, 1518815.49495509, 1518815.49495509, 1518815.49495509, 
    1518815.49495509, 1518815.49495509, 1518815.49495509, 1518815.49495509, 
    1518815.49495509, 1518815.49495509, 1518815.49495509, 1518815.49495509, 
    1518815.49495509, 1518815.49495509, 1518815.49495509, 1518815.49495509, 
    1518815.49495509, 1518815.49495509, 1518815.49495509, 1518815.49495509, 
    1518815.49495509, 1518815.49495509, 1518815.49495509, 1518815.49495509, 
    1518815.49495509, 1518815.49495509, 1518815.49495509, 1518815.49495509, 
    1518815.49495509, 1518815.49495509, 1518815.49495509, 1518815.49495509, 
    1518815.49495509, 1518815.49495509, 1518815.49495509, 1518815.49495509, 
    1518815.49495509, 1518815.49495509, 1518815.49495509, 1518815.49495509,
  1555859.77531985, 1555859.77531985, 1555859.77531985, 1555859.77531985, 
    1555859.77531985, 1555859.77531985, 1555859.77531985, 1555859.77531985, 
    1555859.77531985, 1555859.77531985, 1555859.77531985, 1555859.77531985, 
    1555859.77531985, 1555859.77531985, 1555859.77531985, 1555859.77531985, 
    1555859.77531985, 1555859.77531985, 1555859.77531985, 1555859.77531985, 
    1555859.77531985, 1555859.77531985, 1555859.77531985, 1555859.77531985, 
    1555859.77531985, 1555859.77531985, 1555859.77531985, 1555859.77531985, 
    1555859.77531985, 1555859.77531985, 1555859.77531985, 1555859.77531985, 
    1555859.77531985, 1555859.77531985, 1555859.77531985, 1555859.77531985, 
    1555859.77531985, 1555859.77531985, 1555859.77531985, 1555859.77531985, 
    1555859.77531985, 1555859.77531985, 1555859.77531985, 1555859.77531985, 
    1555859.77531985, 1555859.77531985, 1555859.77531985, 1555859.77531985, 
    1555859.77531985, 1555859.77531985, 1555859.77531985, 1555859.77531985, 
    1555859.77531985, 1555859.77531985, 1555859.77531985, 1555859.77531985,
  1592904.05568461, 1592904.05568461, 1592904.05568461, 1592904.05568461, 
    1592904.05568461, 1592904.05568461, 1592904.05568461, 1592904.05568461, 
    1592904.05568461, 1592904.05568461, 1592904.05568461, 1592904.05568461, 
    1592904.05568461, 1592904.05568461, 1592904.05568461, 1592904.05568461, 
    1592904.05568461, 1592904.05568461, 1592904.05568461, 1592904.05568461, 
    1592904.05568461, 1592904.05568461, 1592904.05568461, 1592904.05568461, 
    1592904.05568461, 1592904.05568461, 1592904.05568461, 1592904.05568461, 
    1592904.05568461, 1592904.05568461, 1592904.05568461, 1592904.05568461, 
    1592904.05568461, 1592904.05568461, 1592904.05568461, 1592904.05568461, 
    1592904.05568461, 1592904.05568461, 1592904.05568461, 1592904.05568461, 
    1592904.05568461, 1592904.05568461, 1592904.05568461, 1592904.05568461, 
    1592904.05568461, 1592904.05568461, 1592904.05568461, 1592904.05568461, 
    1592904.05568461, 1592904.05568461, 1592904.05568461, 1592904.05568461, 
    1592904.05568461, 1592904.05568461, 1592904.05568461, 1592904.05568461,
  1629948.33604937, 1629948.33604937, 1629948.33604937, 1629948.33604937, 
    1629948.33604937, 1629948.33604937, 1629948.33604937, 1629948.33604937, 
    1629948.33604937, 1629948.33604937, 1629948.33604937, 1629948.33604937, 
    1629948.33604937, 1629948.33604937, 1629948.33604937, 1629948.33604937, 
    1629948.33604937, 1629948.33604937, 1629948.33604937, 1629948.33604937, 
    1629948.33604937, 1629948.33604937, 1629948.33604937, 1629948.33604937, 
    1629948.33604937, 1629948.33604937, 1629948.33604937, 1629948.33604937, 
    1629948.33604937, 1629948.33604937, 1629948.33604937, 1629948.33604937, 
    1629948.33604937, 1629948.33604937, 1629948.33604937, 1629948.33604937, 
    1629948.33604937, 1629948.33604937, 1629948.33604937, 1629948.33604937, 
    1629948.33604937, 1629948.33604937, 1629948.33604937, 1629948.33604937, 
    1629948.33604937, 1629948.33604937, 1629948.33604937, 1629948.33604937, 
    1629948.33604937, 1629948.33604937, 1629948.33604937, 1629948.33604937, 
    1629948.33604937, 1629948.33604937, 1629948.33604937, 1629948.33604937,
  1666992.61641413, 1666992.61641413, 1666992.61641413, 1666992.61641413, 
    1666992.61641413, 1666992.61641413, 1666992.61641413, 1666992.61641413, 
    1666992.61641413, 1666992.61641413, 1666992.61641413, 1666992.61641413, 
    1666992.61641413, 1666992.61641413, 1666992.61641413, 1666992.61641413, 
    1666992.61641413, 1666992.61641413, 1666992.61641413, 1666992.61641413, 
    1666992.61641413, 1666992.61641413, 1666992.61641413, 1666992.61641413, 
    1666992.61641413, 1666992.61641413, 1666992.61641413, 1666992.61641413, 
    1666992.61641413, 1666992.61641413, 1666992.61641413, 1666992.61641413, 
    1666992.61641413, 1666992.61641413, 1666992.61641413, 1666992.61641413, 
    1666992.61641413, 1666992.61641413, 1666992.61641413, 1666992.61641413, 
    1666992.61641413, 1666992.61641413, 1666992.61641413, 1666992.61641413, 
    1666992.61641413, 1666992.61641413, 1666992.61641413, 1666992.61641413, 
    1666992.61641413, 1666992.61641413, 1666992.61641413, 1666992.61641413, 
    1666992.61641413, 1666992.61641413, 1666992.61641413, 1666992.61641413,
  1704036.89677889, 1704036.89677889, 1704036.89677889, 1704036.89677889, 
    1704036.89677889, 1704036.89677889, 1704036.89677889, 1704036.89677889, 
    1704036.89677889, 1704036.89677889, 1704036.89677889, 1704036.89677889, 
    1704036.89677889, 1704036.89677889, 1704036.89677889, 1704036.89677889, 
    1704036.89677889, 1704036.89677889, 1704036.89677889, 1704036.89677889, 
    1704036.89677889, 1704036.89677889, 1704036.89677889, 1704036.89677889, 
    1704036.89677889, 1704036.89677889, 1704036.89677889, 1704036.89677889, 
    1704036.89677889, 1704036.89677889, 1704036.89677889, 1704036.89677889, 
    1704036.89677889, 1704036.89677889, 1704036.89677889, 1704036.89677889, 
    1704036.89677889, 1704036.89677889, 1704036.89677889, 1704036.89677889, 
    1704036.89677889, 1704036.89677889, 1704036.89677889, 1704036.89677889, 
    1704036.89677889, 1704036.89677889, 1704036.89677889, 1704036.89677889, 
    1704036.89677889, 1704036.89677889, 1704036.89677889, 1704036.89677889, 
    1704036.89677889, 1704036.89677889, 1704036.89677889, 1704036.89677889,
  1741081.17714364, 1741081.17714364, 1741081.17714364, 1741081.17714364, 
    1741081.17714364, 1741081.17714364, 1741081.17714364, 1741081.17714364, 
    1741081.17714364, 1741081.17714364, 1741081.17714364, 1741081.17714364, 
    1741081.17714364, 1741081.17714364, 1741081.17714364, 1741081.17714364, 
    1741081.17714364, 1741081.17714364, 1741081.17714364, 1741081.17714364, 
    1741081.17714364, 1741081.17714364, 1741081.17714364, 1741081.17714364, 
    1741081.17714364, 1741081.17714364, 1741081.17714364, 1741081.17714364, 
    1741081.17714364, 1741081.17714364, 1741081.17714364, 1741081.17714364, 
    1741081.17714364, 1741081.17714364, 1741081.17714364, 1741081.17714364, 
    1741081.17714364, 1741081.17714364, 1741081.17714364, 1741081.17714364, 
    1741081.17714364, 1741081.17714364, 1741081.17714364, 1741081.17714364, 
    1741081.17714364, 1741081.17714364, 1741081.17714364, 1741081.17714364, 
    1741081.17714364, 1741081.17714364, 1741081.17714364, 1741081.17714364, 
    1741081.17714364, 1741081.17714364, 1741081.17714364, 1741081.17714364,
  1778125.4575084, 1778125.4575084, 1778125.4575084, 1778125.4575084, 
    1778125.4575084, 1778125.4575084, 1778125.4575084, 1778125.4575084, 
    1778125.4575084, 1778125.4575084, 1778125.4575084, 1778125.4575084, 
    1778125.4575084, 1778125.4575084, 1778125.4575084, 1778125.4575084, 
    1778125.4575084, 1778125.4575084, 1778125.4575084, 1778125.4575084, 
    1778125.4575084, 1778125.4575084, 1778125.4575084, 1778125.4575084, 
    1778125.4575084, 1778125.4575084, 1778125.4575084, 1778125.4575084, 
    1778125.4575084, 1778125.4575084, 1778125.4575084, 1778125.4575084, 
    1778125.4575084, 1778125.4575084, 1778125.4575084, 1778125.4575084, 
    1778125.4575084, 1778125.4575084, 1778125.4575084, 1778125.4575084, 
    1778125.4575084, 1778125.4575084, 1778125.4575084, 1778125.4575084, 
    1778125.4575084, 1778125.4575084, 1778125.4575084, 1778125.4575084, 
    1778125.4575084, 1778125.4575084, 1778125.4575084, 1778125.4575084, 
    1778125.4575084, 1778125.4575084, 1778125.4575084, 1778125.4575084,
  1815169.73787316, 1815169.73787316, 1815169.73787316, 1815169.73787316, 
    1815169.73787316, 1815169.73787316, 1815169.73787316, 1815169.73787316, 
    1815169.73787316, 1815169.73787316, 1815169.73787316, 1815169.73787316, 
    1815169.73787316, 1815169.73787316, 1815169.73787316, 1815169.73787316, 
    1815169.73787316, 1815169.73787316, 1815169.73787316, 1815169.73787316, 
    1815169.73787316, 1815169.73787316, 1815169.73787316, 1815169.73787316, 
    1815169.73787316, 1815169.73787316, 1815169.73787316, 1815169.73787316, 
    1815169.73787316, 1815169.73787316, 1815169.73787316, 1815169.73787316, 
    1815169.73787316, 1815169.73787316, 1815169.73787316, 1815169.73787316, 
    1815169.73787316, 1815169.73787316, 1815169.73787316, 1815169.73787316, 
    1815169.73787316, 1815169.73787316, 1815169.73787316, 1815169.73787316, 
    1815169.73787316, 1815169.73787316, 1815169.73787316, 1815169.73787316, 
    1815169.73787316, 1815169.73787316, 1815169.73787316, 1815169.73787316, 
    1815169.73787316, 1815169.73787316, 1815169.73787316, 1815169.73787316,
  1852214.01823792, 1852214.01823792, 1852214.01823792, 1852214.01823792, 
    1852214.01823792, 1852214.01823792, 1852214.01823792, 1852214.01823792, 
    1852214.01823792, 1852214.01823792, 1852214.01823792, 1852214.01823792, 
    1852214.01823792, 1852214.01823792, 1852214.01823792, 1852214.01823792, 
    1852214.01823792, 1852214.01823792, 1852214.01823792, 1852214.01823792, 
    1852214.01823792, 1852214.01823792, 1852214.01823792, 1852214.01823792, 
    1852214.01823792, 1852214.01823792, 1852214.01823792, 1852214.01823792, 
    1852214.01823792, 1852214.01823792, 1852214.01823792, 1852214.01823792, 
    1852214.01823792, 1852214.01823792, 1852214.01823792, 1852214.01823792, 
    1852214.01823792, 1852214.01823792, 1852214.01823792, 1852214.01823792, 
    1852214.01823792, 1852214.01823792, 1852214.01823792, 1852214.01823792, 
    1852214.01823792, 1852214.01823792, 1852214.01823792, 1852214.01823792, 
    1852214.01823792, 1852214.01823792, 1852214.01823792, 1852214.01823792, 
    1852214.01823792, 1852214.01823792, 1852214.01823792, 1852214.01823792,
  1889258.29860268, 1889258.29860268, 1889258.29860268, 1889258.29860268, 
    1889258.29860268, 1889258.29860268, 1889258.29860268, 1889258.29860268, 
    1889258.29860268, 1889258.29860268, 1889258.29860268, 1889258.29860268, 
    1889258.29860268, 1889258.29860268, 1889258.29860268, 1889258.29860268, 
    1889258.29860268, 1889258.29860268, 1889258.29860268, 1889258.29860268, 
    1889258.29860268, 1889258.29860268, 1889258.29860268, 1889258.29860268, 
    1889258.29860268, 1889258.29860268, 1889258.29860268, 1889258.29860268, 
    1889258.29860268, 1889258.29860268, 1889258.29860268, 1889258.29860268, 
    1889258.29860268, 1889258.29860268, 1889258.29860268, 1889258.29860268, 
    1889258.29860268, 1889258.29860268, 1889258.29860268, 1889258.29860268, 
    1889258.29860268, 1889258.29860268, 1889258.29860268, 1889258.29860268, 
    1889258.29860268, 1889258.29860268, 1889258.29860268, 1889258.29860268, 
    1889258.29860268, 1889258.29860268, 1889258.29860268, 1889258.29860268, 
    1889258.29860268, 1889258.29860268, 1889258.29860268, 1889258.29860268,
  1926302.57896744, 1926302.57896744, 1926302.57896744, 1926302.57896744, 
    1926302.57896744, 1926302.57896744, 1926302.57896744, 1926302.57896744, 
    1926302.57896744, 1926302.57896744, 1926302.57896744, 1926302.57896744, 
    1926302.57896744, 1926302.57896744, 1926302.57896744, 1926302.57896744, 
    1926302.57896744, 1926302.57896744, 1926302.57896744, 1926302.57896744, 
    1926302.57896744, 1926302.57896744, 1926302.57896744, 1926302.57896744, 
    1926302.57896744, 1926302.57896744, 1926302.57896744, 1926302.57896744, 
    1926302.57896744, 1926302.57896744, 1926302.57896744, 1926302.57896744, 
    1926302.57896744, 1926302.57896744, 1926302.57896744, 1926302.57896744, 
    1926302.57896744, 1926302.57896744, 1926302.57896744, 1926302.57896744, 
    1926302.57896744, 1926302.57896744, 1926302.57896744, 1926302.57896744, 
    1926302.57896744, 1926302.57896744, 1926302.57896744, 1926302.57896744, 
    1926302.57896744, 1926302.57896744, 1926302.57896744, 1926302.57896744, 
    1926302.57896744, 1926302.57896744, 1926302.57896744, 1926302.57896744,
  1963346.85933219, 1963346.85933219, 1963346.85933219, 1963346.85933219, 
    1963346.85933219, 1963346.85933219, 1963346.85933219, 1963346.85933219, 
    1963346.85933219, 1963346.85933219, 1963346.85933219, 1963346.85933219, 
    1963346.85933219, 1963346.85933219, 1963346.85933219, 1963346.85933219, 
    1963346.85933219, 1963346.85933219, 1963346.85933219, 1963346.85933219, 
    1963346.85933219, 1963346.85933219, 1963346.85933219, 1963346.85933219, 
    1963346.85933219, 1963346.85933219, 1963346.85933219, 1963346.85933219, 
    1963346.85933219, 1963346.85933219, 1963346.85933219, 1963346.85933219, 
    1963346.85933219, 1963346.85933219, 1963346.85933219, 1963346.85933219, 
    1963346.85933219, 1963346.85933219, 1963346.85933219, 1963346.85933219, 
    1963346.85933219, 1963346.85933219, 1963346.85933219, 1963346.85933219, 
    1963346.85933219, 1963346.85933219, 1963346.85933219, 1963346.85933219, 
    1963346.85933219, 1963346.85933219, 1963346.85933219, 1963346.85933219, 
    1963346.85933219, 1963346.85933219, 1963346.85933219, 1963346.85933219,
  2000391.13969695, 2000391.13969695, 2000391.13969695, 2000391.13969695, 
    2000391.13969695, 2000391.13969695, 2000391.13969695, 2000391.13969695, 
    2000391.13969695, 2000391.13969695, 2000391.13969695, 2000391.13969695, 
    2000391.13969695, 2000391.13969695, 2000391.13969695, 2000391.13969695, 
    2000391.13969695, 2000391.13969695, 2000391.13969695, 2000391.13969695, 
    2000391.13969695, 2000391.13969695, 2000391.13969695, 2000391.13969695, 
    2000391.13969695, 2000391.13969695, 2000391.13969695, 2000391.13969695, 
    2000391.13969695, 2000391.13969695, 2000391.13969695, 2000391.13969695, 
    2000391.13969695, 2000391.13969695, 2000391.13969695, 2000391.13969695, 
    2000391.13969695, 2000391.13969695, 2000391.13969695, 2000391.13969695, 
    2000391.13969695, 2000391.13969695, 2000391.13969695, 2000391.13969695, 
    2000391.13969695, 2000391.13969695, 2000391.13969695, 2000391.13969695, 
    2000391.13969695, 2000391.13969695, 2000391.13969695, 2000391.13969695, 
    2000391.13969695, 2000391.13969695, 2000391.13969695, 2000391.13969695 ;

 y_u =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  37044.2803647582, 37044.2803647582, 37044.2803647582, 37044.2803647582, 
    37044.2803647582, 37044.2803647582, 37044.2803647582, 37044.2803647582, 
    37044.2803647582, 37044.2803647582, 37044.2803647582, 37044.2803647582, 
    37044.2803647582, 37044.2803647582, 37044.2803647582, 37044.2803647582, 
    37044.2803647582, 37044.2803647582, 37044.2803647582, 37044.2803647582, 
    37044.2803647582, 37044.2803647582, 37044.2803647582, 37044.2803647582, 
    37044.2803647582, 37044.2803647582, 37044.2803647582, 37044.2803647582, 
    37044.2803647582, 37044.2803647582, 37044.2803647582, 37044.2803647582, 
    37044.2803647582, 37044.2803647582, 37044.2803647582, 37044.2803647582, 
    37044.2803647582, 37044.2803647582, 37044.2803647582, 37044.2803647582, 
    37044.2803647582, 37044.2803647582, 37044.2803647582, 37044.2803647582, 
    37044.2803647582, 37044.2803647582, 37044.2803647582, 37044.2803647582, 
    37044.2803647582, 37044.2803647582, 37044.2803647582, 37044.2803647582, 
    37044.2803647582, 37044.2803647582, 37044.2803647582,
  74088.5607295167, 74088.5607295167, 74088.5607295167, 74088.5607295167, 
    74088.5607295167, 74088.5607295167, 74088.5607295167, 74088.5607295167, 
    74088.5607295167, 74088.5607295167, 74088.5607295167, 74088.5607295167, 
    74088.5607295167, 74088.5607295167, 74088.5607295167, 74088.5607295167, 
    74088.5607295167, 74088.5607295167, 74088.5607295167, 74088.5607295167, 
    74088.5607295167, 74088.5607295167, 74088.5607295167, 74088.5607295167, 
    74088.5607295167, 74088.5607295167, 74088.5607295167, 74088.5607295167, 
    74088.5607295167, 74088.5607295167, 74088.5607295167, 74088.5607295167, 
    74088.5607295167, 74088.5607295167, 74088.5607295167, 74088.5607295167, 
    74088.5607295167, 74088.5607295167, 74088.5607295167, 74088.5607295167, 
    74088.5607295167, 74088.5607295167, 74088.5607295167, 74088.5607295167, 
    74088.5607295167, 74088.5607295167, 74088.5607295167, 74088.5607295167, 
    74088.5607295167, 74088.5607295167, 74088.5607295167, 74088.5607295167, 
    74088.5607295167, 74088.5607295167, 74088.5607295167,
  111132.841094275, 111132.841094275, 111132.841094275, 111132.841094275, 
    111132.841094275, 111132.841094275, 111132.841094275, 111132.841094275, 
    111132.841094275, 111132.841094275, 111132.841094275, 111132.841094275, 
    111132.841094275, 111132.841094275, 111132.841094275, 111132.841094275, 
    111132.841094275, 111132.841094275, 111132.841094275, 111132.841094275, 
    111132.841094275, 111132.841094275, 111132.841094275, 111132.841094275, 
    111132.841094275, 111132.841094275, 111132.841094275, 111132.841094275, 
    111132.841094275, 111132.841094275, 111132.841094275, 111132.841094275, 
    111132.841094275, 111132.841094275, 111132.841094275, 111132.841094275, 
    111132.841094275, 111132.841094275, 111132.841094275, 111132.841094275, 
    111132.841094275, 111132.841094275, 111132.841094275, 111132.841094275, 
    111132.841094275, 111132.841094275, 111132.841094275, 111132.841094275, 
    111132.841094275, 111132.841094275, 111132.841094275, 111132.841094275, 
    111132.841094275, 111132.841094275, 111132.841094275,
  148177.121459033, 148177.121459033, 148177.121459033, 148177.121459033, 
    148177.121459033, 148177.121459033, 148177.121459033, 148177.121459033, 
    148177.121459033, 148177.121459033, 148177.121459033, 148177.121459033, 
    148177.121459033, 148177.121459033, 148177.121459033, 148177.121459033, 
    148177.121459033, 148177.121459033, 148177.121459033, 148177.121459033, 
    148177.121459033, 148177.121459033, 148177.121459033, 148177.121459033, 
    148177.121459033, 148177.121459033, 148177.121459033, 148177.121459033, 
    148177.121459033, 148177.121459033, 148177.121459033, 148177.121459033, 
    148177.121459033, 148177.121459033, 148177.121459033, 148177.121459033, 
    148177.121459033, 148177.121459033, 148177.121459033, 148177.121459033, 
    148177.121459033, 148177.121459033, 148177.121459033, 148177.121459033, 
    148177.121459033, 148177.121459033, 148177.121459033, 148177.121459033, 
    148177.121459033, 148177.121459033, 148177.121459033, 148177.121459033, 
    148177.121459033, 148177.121459033, 148177.121459033,
  185221.401823792, 185221.401823792, 185221.401823792, 185221.401823792, 
    185221.401823792, 185221.401823792, 185221.401823792, 185221.401823792, 
    185221.401823792, 185221.401823792, 185221.401823792, 185221.401823792, 
    185221.401823792, 185221.401823792, 185221.401823792, 185221.401823792, 
    185221.401823792, 185221.401823792, 185221.401823792, 185221.401823792, 
    185221.401823792, 185221.401823792, 185221.401823792, 185221.401823792, 
    185221.401823792, 185221.401823792, 185221.401823792, 185221.401823792, 
    185221.401823792, 185221.401823792, 185221.401823792, 185221.401823792, 
    185221.401823792, 185221.401823792, 185221.401823792, 185221.401823792, 
    185221.401823792, 185221.401823792, 185221.401823792, 185221.401823792, 
    185221.401823792, 185221.401823792, 185221.401823792, 185221.401823792, 
    185221.401823792, 185221.401823792, 185221.401823792, 185221.401823792, 
    185221.401823792, 185221.401823792, 185221.401823792, 185221.401823792, 
    185221.401823792, 185221.401823792, 185221.401823792,
  222265.682188551, 222265.682188551, 222265.682188551, 222265.682188551, 
    222265.682188551, 222265.682188551, 222265.682188551, 222265.682188551, 
    222265.682188551, 222265.682188551, 222265.682188551, 222265.682188551, 
    222265.682188551, 222265.682188551, 222265.682188551, 222265.682188551, 
    222265.682188551, 222265.682188551, 222265.682188551, 222265.682188551, 
    222265.682188551, 222265.682188551, 222265.682188551, 222265.682188551, 
    222265.682188551, 222265.682188551, 222265.682188551, 222265.682188551, 
    222265.682188551, 222265.682188551, 222265.682188551, 222265.682188551, 
    222265.682188551, 222265.682188551, 222265.682188551, 222265.682188551, 
    222265.682188551, 222265.682188551, 222265.682188551, 222265.682188551, 
    222265.682188551, 222265.682188551, 222265.682188551, 222265.682188551, 
    222265.682188551, 222265.682188551, 222265.682188551, 222265.682188551, 
    222265.682188551, 222265.682188551, 222265.682188551, 222265.682188551, 
    222265.682188551, 222265.682188551, 222265.682188551,
  259309.962553309, 259309.962553309, 259309.962553309, 259309.962553309, 
    259309.962553309, 259309.962553309, 259309.962553309, 259309.962553309, 
    259309.962553309, 259309.962553309, 259309.962553309, 259309.962553309, 
    259309.962553309, 259309.962553309, 259309.962553309, 259309.962553309, 
    259309.962553309, 259309.962553309, 259309.962553309, 259309.962553309, 
    259309.962553309, 259309.962553309, 259309.962553309, 259309.962553309, 
    259309.962553309, 259309.962553309, 259309.962553309, 259309.962553309, 
    259309.962553309, 259309.962553309, 259309.962553309, 259309.962553309, 
    259309.962553309, 259309.962553309, 259309.962553309, 259309.962553309, 
    259309.962553309, 259309.962553309, 259309.962553309, 259309.962553309, 
    259309.962553309, 259309.962553309, 259309.962553309, 259309.962553309, 
    259309.962553309, 259309.962553309, 259309.962553309, 259309.962553309, 
    259309.962553309, 259309.962553309, 259309.962553309, 259309.962553309, 
    259309.962553309, 259309.962553309, 259309.962553309,
  296354.242918067, 296354.242918067, 296354.242918067, 296354.242918067, 
    296354.242918067, 296354.242918067, 296354.242918067, 296354.242918067, 
    296354.242918067, 296354.242918067, 296354.242918067, 296354.242918067, 
    296354.242918067, 296354.242918067, 296354.242918067, 296354.242918067, 
    296354.242918067, 296354.242918067, 296354.242918067, 296354.242918067, 
    296354.242918067, 296354.242918067, 296354.242918067, 296354.242918067, 
    296354.242918067, 296354.242918067, 296354.242918067, 296354.242918067, 
    296354.242918067, 296354.242918067, 296354.242918067, 296354.242918067, 
    296354.242918067, 296354.242918067, 296354.242918067, 296354.242918067, 
    296354.242918067, 296354.242918067, 296354.242918067, 296354.242918067, 
    296354.242918067, 296354.242918067, 296354.242918067, 296354.242918067, 
    296354.242918067, 296354.242918067, 296354.242918067, 296354.242918067, 
    296354.242918067, 296354.242918067, 296354.242918067, 296354.242918067, 
    296354.242918067, 296354.242918067, 296354.242918067,
  333398.523282826, 333398.523282826, 333398.523282826, 333398.523282826, 
    333398.523282826, 333398.523282826, 333398.523282826, 333398.523282826, 
    333398.523282826, 333398.523282826, 333398.523282826, 333398.523282826, 
    333398.523282826, 333398.523282826, 333398.523282826, 333398.523282826, 
    333398.523282826, 333398.523282826, 333398.523282826, 333398.523282826, 
    333398.523282826, 333398.523282826, 333398.523282826, 333398.523282826, 
    333398.523282826, 333398.523282826, 333398.523282826, 333398.523282826, 
    333398.523282826, 333398.523282826, 333398.523282826, 333398.523282826, 
    333398.523282826, 333398.523282826, 333398.523282826, 333398.523282826, 
    333398.523282826, 333398.523282826, 333398.523282826, 333398.523282826, 
    333398.523282826, 333398.523282826, 333398.523282826, 333398.523282826, 
    333398.523282826, 333398.523282826, 333398.523282826, 333398.523282826, 
    333398.523282826, 333398.523282826, 333398.523282826, 333398.523282826, 
    333398.523282826, 333398.523282826, 333398.523282826,
  370442.803647584, 370442.803647584, 370442.803647584, 370442.803647584, 
    370442.803647584, 370442.803647584, 370442.803647584, 370442.803647584, 
    370442.803647584, 370442.803647584, 370442.803647584, 370442.803647584, 
    370442.803647584, 370442.803647584, 370442.803647584, 370442.803647584, 
    370442.803647584, 370442.803647584, 370442.803647584, 370442.803647584, 
    370442.803647584, 370442.803647584, 370442.803647584, 370442.803647584, 
    370442.803647584, 370442.803647584, 370442.803647584, 370442.803647584, 
    370442.803647584, 370442.803647584, 370442.803647584, 370442.803647584, 
    370442.803647584, 370442.803647584, 370442.803647584, 370442.803647584, 
    370442.803647584, 370442.803647584, 370442.803647584, 370442.803647584, 
    370442.803647584, 370442.803647584, 370442.803647584, 370442.803647584, 
    370442.803647584, 370442.803647584, 370442.803647584, 370442.803647584, 
    370442.803647584, 370442.803647584, 370442.803647584, 370442.803647584, 
    370442.803647584, 370442.803647584, 370442.803647584,
  407487.084012342, 407487.084012342, 407487.084012342, 407487.084012342, 
    407487.084012342, 407487.084012342, 407487.084012342, 407487.084012342, 
    407487.084012342, 407487.084012342, 407487.084012342, 407487.084012342, 
    407487.084012342, 407487.084012342, 407487.084012342, 407487.084012342, 
    407487.084012342, 407487.084012342, 407487.084012342, 407487.084012342, 
    407487.084012342, 407487.084012342, 407487.084012342, 407487.084012342, 
    407487.084012342, 407487.084012342, 407487.084012342, 407487.084012342, 
    407487.084012342, 407487.084012342, 407487.084012342, 407487.084012342, 
    407487.084012342, 407487.084012342, 407487.084012342, 407487.084012342, 
    407487.084012342, 407487.084012342, 407487.084012342, 407487.084012342, 
    407487.084012342, 407487.084012342, 407487.084012342, 407487.084012342, 
    407487.084012342, 407487.084012342, 407487.084012342, 407487.084012342, 
    407487.084012342, 407487.084012342, 407487.084012342, 407487.084012342, 
    407487.084012342, 407487.084012342, 407487.084012342,
  444531.364377101, 444531.364377101, 444531.364377101, 444531.364377101, 
    444531.364377101, 444531.364377101, 444531.364377101, 444531.364377101, 
    444531.364377101, 444531.364377101, 444531.364377101, 444531.364377101, 
    444531.364377101, 444531.364377101, 444531.364377101, 444531.364377101, 
    444531.364377101, 444531.364377101, 444531.364377101, 444531.364377101, 
    444531.364377101, 444531.364377101, 444531.364377101, 444531.364377101, 
    444531.364377101, 444531.364377101, 444531.364377101, 444531.364377101, 
    444531.364377101, 444531.364377101, 444531.364377101, 444531.364377101, 
    444531.364377101, 444531.364377101, 444531.364377101, 444531.364377101, 
    444531.364377101, 444531.364377101, 444531.364377101, 444531.364377101, 
    444531.364377101, 444531.364377101, 444531.364377101, 444531.364377101, 
    444531.364377101, 444531.364377101, 444531.364377101, 444531.364377101, 
    444531.364377101, 444531.364377101, 444531.364377101, 444531.364377101, 
    444531.364377101, 444531.364377101, 444531.364377101,
  481575.644741859, 481575.644741859, 481575.644741859, 481575.644741859, 
    481575.644741859, 481575.644741859, 481575.644741859, 481575.644741859, 
    481575.644741859, 481575.644741859, 481575.644741859, 481575.644741859, 
    481575.644741859, 481575.644741859, 481575.644741859, 481575.644741859, 
    481575.644741859, 481575.644741859, 481575.644741859, 481575.644741859, 
    481575.644741859, 481575.644741859, 481575.644741859, 481575.644741859, 
    481575.644741859, 481575.644741859, 481575.644741859, 481575.644741859, 
    481575.644741859, 481575.644741859, 481575.644741859, 481575.644741859, 
    481575.644741859, 481575.644741859, 481575.644741859, 481575.644741859, 
    481575.644741859, 481575.644741859, 481575.644741859, 481575.644741859, 
    481575.644741859, 481575.644741859, 481575.644741859, 481575.644741859, 
    481575.644741859, 481575.644741859, 481575.644741859, 481575.644741859, 
    481575.644741859, 481575.644741859, 481575.644741859, 481575.644741859, 
    481575.644741859, 481575.644741859, 481575.644741859,
  518619.925106617, 518619.925106617, 518619.925106617, 518619.925106617, 
    518619.925106617, 518619.925106617, 518619.925106617, 518619.925106617, 
    518619.925106617, 518619.925106617, 518619.925106617, 518619.925106617, 
    518619.925106617, 518619.925106617, 518619.925106617, 518619.925106617, 
    518619.925106617, 518619.925106617, 518619.925106617, 518619.925106617, 
    518619.925106617, 518619.925106617, 518619.925106617, 518619.925106617, 
    518619.925106617, 518619.925106617, 518619.925106617, 518619.925106617, 
    518619.925106617, 518619.925106617, 518619.925106617, 518619.925106617, 
    518619.925106617, 518619.925106617, 518619.925106617, 518619.925106617, 
    518619.925106617, 518619.925106617, 518619.925106617, 518619.925106617, 
    518619.925106617, 518619.925106617, 518619.925106617, 518619.925106617, 
    518619.925106617, 518619.925106617, 518619.925106617, 518619.925106617, 
    518619.925106617, 518619.925106617, 518619.925106617, 518619.925106617, 
    518619.925106617, 518619.925106617, 518619.925106617,
  555664.205471375, 555664.205471375, 555664.205471375, 555664.205471375, 
    555664.205471375, 555664.205471375, 555664.205471375, 555664.205471375, 
    555664.205471375, 555664.205471375, 555664.205471375, 555664.205471375, 
    555664.205471375, 555664.205471375, 555664.205471375, 555664.205471375, 
    555664.205471375, 555664.205471375, 555664.205471375, 555664.205471375, 
    555664.205471375, 555664.205471375, 555664.205471375, 555664.205471375, 
    555664.205471375, 555664.205471375, 555664.205471375, 555664.205471375, 
    555664.205471375, 555664.205471375, 555664.205471375, 555664.205471375, 
    555664.205471375, 555664.205471375, 555664.205471375, 555664.205471375, 
    555664.205471375, 555664.205471375, 555664.205471375, 555664.205471375, 
    555664.205471375, 555664.205471375, 555664.205471375, 555664.205471375, 
    555664.205471375, 555664.205471375, 555664.205471375, 555664.205471375, 
    555664.205471375, 555664.205471375, 555664.205471375, 555664.205471375, 
    555664.205471375, 555664.205471375, 555664.205471375,
  592708.485836134, 592708.485836134, 592708.485836134, 592708.485836134, 
    592708.485836134, 592708.485836134, 592708.485836134, 592708.485836134, 
    592708.485836134, 592708.485836134, 592708.485836134, 592708.485836134, 
    592708.485836134, 592708.485836134, 592708.485836134, 592708.485836134, 
    592708.485836134, 592708.485836134, 592708.485836134, 592708.485836134, 
    592708.485836134, 592708.485836134, 592708.485836134, 592708.485836134, 
    592708.485836134, 592708.485836134, 592708.485836134, 592708.485836134, 
    592708.485836134, 592708.485836134, 592708.485836134, 592708.485836134, 
    592708.485836134, 592708.485836134, 592708.485836134, 592708.485836134, 
    592708.485836134, 592708.485836134, 592708.485836134, 592708.485836134, 
    592708.485836134, 592708.485836134, 592708.485836134, 592708.485836134, 
    592708.485836134, 592708.485836134, 592708.485836134, 592708.485836134, 
    592708.485836134, 592708.485836134, 592708.485836134, 592708.485836134, 
    592708.485836134, 592708.485836134, 592708.485836134,
  629752.766200892, 629752.766200892, 629752.766200892, 629752.766200892, 
    629752.766200892, 629752.766200892, 629752.766200892, 629752.766200892, 
    629752.766200892, 629752.766200892, 629752.766200892, 629752.766200892, 
    629752.766200892, 629752.766200892, 629752.766200892, 629752.766200892, 
    629752.766200892, 629752.766200892, 629752.766200892, 629752.766200892, 
    629752.766200892, 629752.766200892, 629752.766200892, 629752.766200892, 
    629752.766200892, 629752.766200892, 629752.766200892, 629752.766200892, 
    629752.766200892, 629752.766200892, 629752.766200892, 629752.766200892, 
    629752.766200892, 629752.766200892, 629752.766200892, 629752.766200892, 
    629752.766200892, 629752.766200892, 629752.766200892, 629752.766200892, 
    629752.766200892, 629752.766200892, 629752.766200892, 629752.766200892, 
    629752.766200892, 629752.766200892, 629752.766200892, 629752.766200892, 
    629752.766200892, 629752.766200892, 629752.766200892, 629752.766200892, 
    629752.766200892, 629752.766200892, 629752.766200892,
  666797.04656565, 666797.04656565, 666797.04656565, 666797.04656565, 
    666797.04656565, 666797.04656565, 666797.04656565, 666797.04656565, 
    666797.04656565, 666797.04656565, 666797.04656565, 666797.04656565, 
    666797.04656565, 666797.04656565, 666797.04656565, 666797.04656565, 
    666797.04656565, 666797.04656565, 666797.04656565, 666797.04656565, 
    666797.04656565, 666797.04656565, 666797.04656565, 666797.04656565, 
    666797.04656565, 666797.04656565, 666797.04656565, 666797.04656565, 
    666797.04656565, 666797.04656565, 666797.04656565, 666797.04656565, 
    666797.04656565, 666797.04656565, 666797.04656565, 666797.04656565, 
    666797.04656565, 666797.04656565, 666797.04656565, 666797.04656565, 
    666797.04656565, 666797.04656565, 666797.04656565, 666797.04656565, 
    666797.04656565, 666797.04656565, 666797.04656565, 666797.04656565, 
    666797.04656565, 666797.04656565, 666797.04656565, 666797.04656565, 
    666797.04656565, 666797.04656565, 666797.04656565,
  703841.326930409, 703841.326930409, 703841.326930409, 703841.326930409, 
    703841.326930409, 703841.326930409, 703841.326930409, 703841.326930409, 
    703841.326930409, 703841.326930409, 703841.326930409, 703841.326930409, 
    703841.326930409, 703841.326930409, 703841.326930409, 703841.326930409, 
    703841.326930409, 703841.326930409, 703841.326930409, 703841.326930409, 
    703841.326930409, 703841.326930409, 703841.326930409, 703841.326930409, 
    703841.326930409, 703841.326930409, 703841.326930409, 703841.326930409, 
    703841.326930409, 703841.326930409, 703841.326930409, 703841.326930409, 
    703841.326930409, 703841.326930409, 703841.326930409, 703841.326930409, 
    703841.326930409, 703841.326930409, 703841.326930409, 703841.326930409, 
    703841.326930409, 703841.326930409, 703841.326930409, 703841.326930409, 
    703841.326930409, 703841.326930409, 703841.326930409, 703841.326930409, 
    703841.326930409, 703841.326930409, 703841.326930409, 703841.326930409, 
    703841.326930409, 703841.326930409, 703841.326930409,
  740885.607295166, 740885.607295166, 740885.607295166, 740885.607295166, 
    740885.607295166, 740885.607295166, 740885.607295166, 740885.607295166, 
    740885.607295166, 740885.607295166, 740885.607295166, 740885.607295166, 
    740885.607295166, 740885.607295166, 740885.607295166, 740885.607295166, 
    740885.607295166, 740885.607295166, 740885.607295166, 740885.607295166, 
    740885.607295166, 740885.607295166, 740885.607295166, 740885.607295166, 
    740885.607295166, 740885.607295166, 740885.607295166, 740885.607295166, 
    740885.607295166, 740885.607295166, 740885.607295166, 740885.607295166, 
    740885.607295166, 740885.607295166, 740885.607295166, 740885.607295166, 
    740885.607295166, 740885.607295166, 740885.607295166, 740885.607295166, 
    740885.607295166, 740885.607295166, 740885.607295166, 740885.607295166, 
    740885.607295166, 740885.607295166, 740885.607295166, 740885.607295166, 
    740885.607295166, 740885.607295166, 740885.607295166, 740885.607295166, 
    740885.607295166, 740885.607295166, 740885.607295166,
  777929.887659925, 777929.887659925, 777929.887659925, 777929.887659925, 
    777929.887659925, 777929.887659925, 777929.887659925, 777929.887659925, 
    777929.887659925, 777929.887659925, 777929.887659925, 777929.887659925, 
    777929.887659925, 777929.887659925, 777929.887659925, 777929.887659925, 
    777929.887659925, 777929.887659925, 777929.887659925, 777929.887659925, 
    777929.887659925, 777929.887659925, 777929.887659925, 777929.887659925, 
    777929.887659925, 777929.887659925, 777929.887659925, 777929.887659925, 
    777929.887659925, 777929.887659925, 777929.887659925, 777929.887659925, 
    777929.887659925, 777929.887659925, 777929.887659925, 777929.887659925, 
    777929.887659925, 777929.887659925, 777929.887659925, 777929.887659925, 
    777929.887659925, 777929.887659925, 777929.887659925, 777929.887659925, 
    777929.887659925, 777929.887659925, 777929.887659925, 777929.887659925, 
    777929.887659925, 777929.887659925, 777929.887659925, 777929.887659925, 
    777929.887659925, 777929.887659925, 777929.887659925,
  814974.168024684, 814974.168024684, 814974.168024684, 814974.168024684, 
    814974.168024684, 814974.168024684, 814974.168024684, 814974.168024684, 
    814974.168024684, 814974.168024684, 814974.168024684, 814974.168024684, 
    814974.168024684, 814974.168024684, 814974.168024684, 814974.168024684, 
    814974.168024684, 814974.168024684, 814974.168024684, 814974.168024684, 
    814974.168024684, 814974.168024684, 814974.168024684, 814974.168024684, 
    814974.168024684, 814974.168024684, 814974.168024684, 814974.168024684, 
    814974.168024684, 814974.168024684, 814974.168024684, 814974.168024684, 
    814974.168024684, 814974.168024684, 814974.168024684, 814974.168024684, 
    814974.168024684, 814974.168024684, 814974.168024684, 814974.168024684, 
    814974.168024684, 814974.168024684, 814974.168024684, 814974.168024684, 
    814974.168024684, 814974.168024684, 814974.168024684, 814974.168024684, 
    814974.168024684, 814974.168024684, 814974.168024684, 814974.168024684, 
    814974.168024684, 814974.168024684, 814974.168024684,
  852018.448389441, 852018.448389441, 852018.448389441, 852018.448389441, 
    852018.448389441, 852018.448389441, 852018.448389441, 852018.448389441, 
    852018.448389441, 852018.448389441, 852018.448389441, 852018.448389441, 
    852018.448389441, 852018.448389441, 852018.448389441, 852018.448389441, 
    852018.448389441, 852018.448389441, 852018.448389441, 852018.448389441, 
    852018.448389441, 852018.448389441, 852018.448389441, 852018.448389441, 
    852018.448389441, 852018.448389441, 852018.448389441, 852018.448389441, 
    852018.448389441, 852018.448389441, 852018.448389441, 852018.448389441, 
    852018.448389441, 852018.448389441, 852018.448389441, 852018.448389441, 
    852018.448389441, 852018.448389441, 852018.448389441, 852018.448389441, 
    852018.448389441, 852018.448389441, 852018.448389441, 852018.448389441, 
    852018.448389441, 852018.448389441, 852018.448389441, 852018.448389441, 
    852018.448389441, 852018.448389441, 852018.448389441, 852018.448389441, 
    852018.448389441, 852018.448389441, 852018.448389441,
  889062.7287542, 889062.7287542, 889062.7287542, 889062.7287542, 
    889062.7287542, 889062.7287542, 889062.7287542, 889062.7287542, 
    889062.7287542, 889062.7287542, 889062.7287542, 889062.7287542, 
    889062.7287542, 889062.7287542, 889062.7287542, 889062.7287542, 
    889062.7287542, 889062.7287542, 889062.7287542, 889062.7287542, 
    889062.7287542, 889062.7287542, 889062.7287542, 889062.7287542, 
    889062.7287542, 889062.7287542, 889062.7287542, 889062.7287542, 
    889062.7287542, 889062.7287542, 889062.7287542, 889062.7287542, 
    889062.7287542, 889062.7287542, 889062.7287542, 889062.7287542, 
    889062.7287542, 889062.7287542, 889062.7287542, 889062.7287542, 
    889062.7287542, 889062.7287542, 889062.7287542, 889062.7287542, 
    889062.7287542, 889062.7287542, 889062.7287542, 889062.7287542, 
    889062.7287542, 889062.7287542, 889062.7287542, 889062.7287542, 
    889062.7287542, 889062.7287542, 889062.7287542,
  926107.009118958, 926107.009118958, 926107.009118958, 926107.009118958, 
    926107.009118958, 926107.009118958, 926107.009118958, 926107.009118958, 
    926107.009118958, 926107.009118958, 926107.009118958, 926107.009118958, 
    926107.009118958, 926107.009118958, 926107.009118958, 926107.009118958, 
    926107.009118958, 926107.009118958, 926107.009118958, 926107.009118958, 
    926107.009118958, 926107.009118958, 926107.009118958, 926107.009118958, 
    926107.009118958, 926107.009118958, 926107.009118958, 926107.009118958, 
    926107.009118958, 926107.009118958, 926107.009118958, 926107.009118958, 
    926107.009118958, 926107.009118958, 926107.009118958, 926107.009118958, 
    926107.009118958, 926107.009118958, 926107.009118958, 926107.009118958, 
    926107.009118958, 926107.009118958, 926107.009118958, 926107.009118958, 
    926107.009118958, 926107.009118958, 926107.009118958, 926107.009118958, 
    926107.009118958, 926107.009118958, 926107.009118958, 926107.009118958, 
    926107.009118958, 926107.009118958, 926107.009118958,
  963151.289483716, 963151.289483716, 963151.289483716, 963151.289483716, 
    963151.289483716, 963151.289483716, 963151.289483716, 963151.289483716, 
    963151.289483716, 963151.289483716, 963151.289483716, 963151.289483716, 
    963151.289483716, 963151.289483716, 963151.289483716, 963151.289483716, 
    963151.289483716, 963151.289483716, 963151.289483716, 963151.289483716, 
    963151.289483716, 963151.289483716, 963151.289483716, 963151.289483716, 
    963151.289483716, 963151.289483716, 963151.289483716, 963151.289483716, 
    963151.289483716, 963151.289483716, 963151.289483716, 963151.289483716, 
    963151.289483716, 963151.289483716, 963151.289483716, 963151.289483716, 
    963151.289483716, 963151.289483716, 963151.289483716, 963151.289483716, 
    963151.289483716, 963151.289483716, 963151.289483716, 963151.289483716, 
    963151.289483716, 963151.289483716, 963151.289483716, 963151.289483716, 
    963151.289483716, 963151.289483716, 963151.289483716, 963151.289483716, 
    963151.289483716, 963151.289483716, 963151.289483716,
  1000195.56984848, 1000195.56984848, 1000195.56984848, 1000195.56984848, 
    1000195.56984848, 1000195.56984848, 1000195.56984848, 1000195.56984848, 
    1000195.56984848, 1000195.56984848, 1000195.56984848, 1000195.56984848, 
    1000195.56984848, 1000195.56984848, 1000195.56984848, 1000195.56984848, 
    1000195.56984848, 1000195.56984848, 1000195.56984848, 1000195.56984848, 
    1000195.56984848, 1000195.56984848, 1000195.56984848, 1000195.56984848, 
    1000195.56984848, 1000195.56984848, 1000195.56984848, 1000195.56984848, 
    1000195.56984848, 1000195.56984848, 1000195.56984848, 1000195.56984848, 
    1000195.56984848, 1000195.56984848, 1000195.56984848, 1000195.56984848, 
    1000195.56984848, 1000195.56984848, 1000195.56984848, 1000195.56984848, 
    1000195.56984848, 1000195.56984848, 1000195.56984848, 1000195.56984848, 
    1000195.56984848, 1000195.56984848, 1000195.56984848, 1000195.56984848, 
    1000195.56984848, 1000195.56984848, 1000195.56984848, 1000195.56984848, 
    1000195.56984848, 1000195.56984848, 1000195.56984848,
  1037239.85021323, 1037239.85021323, 1037239.85021323, 1037239.85021323, 
    1037239.85021323, 1037239.85021323, 1037239.85021323, 1037239.85021323, 
    1037239.85021323, 1037239.85021323, 1037239.85021323, 1037239.85021323, 
    1037239.85021323, 1037239.85021323, 1037239.85021323, 1037239.85021323, 
    1037239.85021323, 1037239.85021323, 1037239.85021323, 1037239.85021323, 
    1037239.85021323, 1037239.85021323, 1037239.85021323, 1037239.85021323, 
    1037239.85021323, 1037239.85021323, 1037239.85021323, 1037239.85021323, 
    1037239.85021323, 1037239.85021323, 1037239.85021323, 1037239.85021323, 
    1037239.85021323, 1037239.85021323, 1037239.85021323, 1037239.85021323, 
    1037239.85021323, 1037239.85021323, 1037239.85021323, 1037239.85021323, 
    1037239.85021323, 1037239.85021323, 1037239.85021323, 1037239.85021323, 
    1037239.85021323, 1037239.85021323, 1037239.85021323, 1037239.85021323, 
    1037239.85021323, 1037239.85021323, 1037239.85021323, 1037239.85021323, 
    1037239.85021323, 1037239.85021323, 1037239.85021323,
  1074284.13057799, 1074284.13057799, 1074284.13057799, 1074284.13057799, 
    1074284.13057799, 1074284.13057799, 1074284.13057799, 1074284.13057799, 
    1074284.13057799, 1074284.13057799, 1074284.13057799, 1074284.13057799, 
    1074284.13057799, 1074284.13057799, 1074284.13057799, 1074284.13057799, 
    1074284.13057799, 1074284.13057799, 1074284.13057799, 1074284.13057799, 
    1074284.13057799, 1074284.13057799, 1074284.13057799, 1074284.13057799, 
    1074284.13057799, 1074284.13057799, 1074284.13057799, 1074284.13057799, 
    1074284.13057799, 1074284.13057799, 1074284.13057799, 1074284.13057799, 
    1074284.13057799, 1074284.13057799, 1074284.13057799, 1074284.13057799, 
    1074284.13057799, 1074284.13057799, 1074284.13057799, 1074284.13057799, 
    1074284.13057799, 1074284.13057799, 1074284.13057799, 1074284.13057799, 
    1074284.13057799, 1074284.13057799, 1074284.13057799, 1074284.13057799, 
    1074284.13057799, 1074284.13057799, 1074284.13057799, 1074284.13057799, 
    1074284.13057799, 1074284.13057799, 1074284.13057799,
  1111328.41094275, 1111328.41094275, 1111328.41094275, 1111328.41094275, 
    1111328.41094275, 1111328.41094275, 1111328.41094275, 1111328.41094275, 
    1111328.41094275, 1111328.41094275, 1111328.41094275, 1111328.41094275, 
    1111328.41094275, 1111328.41094275, 1111328.41094275, 1111328.41094275, 
    1111328.41094275, 1111328.41094275, 1111328.41094275, 1111328.41094275, 
    1111328.41094275, 1111328.41094275, 1111328.41094275, 1111328.41094275, 
    1111328.41094275, 1111328.41094275, 1111328.41094275, 1111328.41094275, 
    1111328.41094275, 1111328.41094275, 1111328.41094275, 1111328.41094275, 
    1111328.41094275, 1111328.41094275, 1111328.41094275, 1111328.41094275, 
    1111328.41094275, 1111328.41094275, 1111328.41094275, 1111328.41094275, 
    1111328.41094275, 1111328.41094275, 1111328.41094275, 1111328.41094275, 
    1111328.41094275, 1111328.41094275, 1111328.41094275, 1111328.41094275, 
    1111328.41094275, 1111328.41094275, 1111328.41094275, 1111328.41094275, 
    1111328.41094275, 1111328.41094275, 1111328.41094275,
  1148372.69130751, 1148372.69130751, 1148372.69130751, 1148372.69130751, 
    1148372.69130751, 1148372.69130751, 1148372.69130751, 1148372.69130751, 
    1148372.69130751, 1148372.69130751, 1148372.69130751, 1148372.69130751, 
    1148372.69130751, 1148372.69130751, 1148372.69130751, 1148372.69130751, 
    1148372.69130751, 1148372.69130751, 1148372.69130751, 1148372.69130751, 
    1148372.69130751, 1148372.69130751, 1148372.69130751, 1148372.69130751, 
    1148372.69130751, 1148372.69130751, 1148372.69130751, 1148372.69130751, 
    1148372.69130751, 1148372.69130751, 1148372.69130751, 1148372.69130751, 
    1148372.69130751, 1148372.69130751, 1148372.69130751, 1148372.69130751, 
    1148372.69130751, 1148372.69130751, 1148372.69130751, 1148372.69130751, 
    1148372.69130751, 1148372.69130751, 1148372.69130751, 1148372.69130751, 
    1148372.69130751, 1148372.69130751, 1148372.69130751, 1148372.69130751, 
    1148372.69130751, 1148372.69130751, 1148372.69130751, 1148372.69130751, 
    1148372.69130751, 1148372.69130751, 1148372.69130751,
  1185416.97167227, 1185416.97167227, 1185416.97167227, 1185416.97167227, 
    1185416.97167227, 1185416.97167227, 1185416.97167227, 1185416.97167227, 
    1185416.97167227, 1185416.97167227, 1185416.97167227, 1185416.97167227, 
    1185416.97167227, 1185416.97167227, 1185416.97167227, 1185416.97167227, 
    1185416.97167227, 1185416.97167227, 1185416.97167227, 1185416.97167227, 
    1185416.97167227, 1185416.97167227, 1185416.97167227, 1185416.97167227, 
    1185416.97167227, 1185416.97167227, 1185416.97167227, 1185416.97167227, 
    1185416.97167227, 1185416.97167227, 1185416.97167227, 1185416.97167227, 
    1185416.97167227, 1185416.97167227, 1185416.97167227, 1185416.97167227, 
    1185416.97167227, 1185416.97167227, 1185416.97167227, 1185416.97167227, 
    1185416.97167227, 1185416.97167227, 1185416.97167227, 1185416.97167227, 
    1185416.97167227, 1185416.97167227, 1185416.97167227, 1185416.97167227, 
    1185416.97167227, 1185416.97167227, 1185416.97167227, 1185416.97167227, 
    1185416.97167227, 1185416.97167227, 1185416.97167227,
  1222461.25203703, 1222461.25203703, 1222461.25203703, 1222461.25203703, 
    1222461.25203703, 1222461.25203703, 1222461.25203703, 1222461.25203703, 
    1222461.25203703, 1222461.25203703, 1222461.25203703, 1222461.25203703, 
    1222461.25203703, 1222461.25203703, 1222461.25203703, 1222461.25203703, 
    1222461.25203703, 1222461.25203703, 1222461.25203703, 1222461.25203703, 
    1222461.25203703, 1222461.25203703, 1222461.25203703, 1222461.25203703, 
    1222461.25203703, 1222461.25203703, 1222461.25203703, 1222461.25203703, 
    1222461.25203703, 1222461.25203703, 1222461.25203703, 1222461.25203703, 
    1222461.25203703, 1222461.25203703, 1222461.25203703, 1222461.25203703, 
    1222461.25203703, 1222461.25203703, 1222461.25203703, 1222461.25203703, 
    1222461.25203703, 1222461.25203703, 1222461.25203703, 1222461.25203703, 
    1222461.25203703, 1222461.25203703, 1222461.25203703, 1222461.25203703, 
    1222461.25203703, 1222461.25203703, 1222461.25203703, 1222461.25203703, 
    1222461.25203703, 1222461.25203703, 1222461.25203703,
  1259505.53240178, 1259505.53240178, 1259505.53240178, 1259505.53240178, 
    1259505.53240178, 1259505.53240178, 1259505.53240178, 1259505.53240178, 
    1259505.53240178, 1259505.53240178, 1259505.53240178, 1259505.53240178, 
    1259505.53240178, 1259505.53240178, 1259505.53240178, 1259505.53240178, 
    1259505.53240178, 1259505.53240178, 1259505.53240178, 1259505.53240178, 
    1259505.53240178, 1259505.53240178, 1259505.53240178, 1259505.53240178, 
    1259505.53240178, 1259505.53240178, 1259505.53240178, 1259505.53240178, 
    1259505.53240178, 1259505.53240178, 1259505.53240178, 1259505.53240178, 
    1259505.53240178, 1259505.53240178, 1259505.53240178, 1259505.53240178, 
    1259505.53240178, 1259505.53240178, 1259505.53240178, 1259505.53240178, 
    1259505.53240178, 1259505.53240178, 1259505.53240178, 1259505.53240178, 
    1259505.53240178, 1259505.53240178, 1259505.53240178, 1259505.53240178, 
    1259505.53240178, 1259505.53240178, 1259505.53240178, 1259505.53240178, 
    1259505.53240178, 1259505.53240178, 1259505.53240178,
  1296549.81276654, 1296549.81276654, 1296549.81276654, 1296549.81276654, 
    1296549.81276654, 1296549.81276654, 1296549.81276654, 1296549.81276654, 
    1296549.81276654, 1296549.81276654, 1296549.81276654, 1296549.81276654, 
    1296549.81276654, 1296549.81276654, 1296549.81276654, 1296549.81276654, 
    1296549.81276654, 1296549.81276654, 1296549.81276654, 1296549.81276654, 
    1296549.81276654, 1296549.81276654, 1296549.81276654, 1296549.81276654, 
    1296549.81276654, 1296549.81276654, 1296549.81276654, 1296549.81276654, 
    1296549.81276654, 1296549.81276654, 1296549.81276654, 1296549.81276654, 
    1296549.81276654, 1296549.81276654, 1296549.81276654, 1296549.81276654, 
    1296549.81276654, 1296549.81276654, 1296549.81276654, 1296549.81276654, 
    1296549.81276654, 1296549.81276654, 1296549.81276654, 1296549.81276654, 
    1296549.81276654, 1296549.81276654, 1296549.81276654, 1296549.81276654, 
    1296549.81276654, 1296549.81276654, 1296549.81276654, 1296549.81276654, 
    1296549.81276654, 1296549.81276654, 1296549.81276654,
  1333594.0931313, 1333594.0931313, 1333594.0931313, 1333594.0931313, 
    1333594.0931313, 1333594.0931313, 1333594.0931313, 1333594.0931313, 
    1333594.0931313, 1333594.0931313, 1333594.0931313, 1333594.0931313, 
    1333594.0931313, 1333594.0931313, 1333594.0931313, 1333594.0931313, 
    1333594.0931313, 1333594.0931313, 1333594.0931313, 1333594.0931313, 
    1333594.0931313, 1333594.0931313, 1333594.0931313, 1333594.0931313, 
    1333594.0931313, 1333594.0931313, 1333594.0931313, 1333594.0931313, 
    1333594.0931313, 1333594.0931313, 1333594.0931313, 1333594.0931313, 
    1333594.0931313, 1333594.0931313, 1333594.0931313, 1333594.0931313, 
    1333594.0931313, 1333594.0931313, 1333594.0931313, 1333594.0931313, 
    1333594.0931313, 1333594.0931313, 1333594.0931313, 1333594.0931313, 
    1333594.0931313, 1333594.0931313, 1333594.0931313, 1333594.0931313, 
    1333594.0931313, 1333594.0931313, 1333594.0931313, 1333594.0931313, 
    1333594.0931313, 1333594.0931313, 1333594.0931313,
  1370638.37349606, 1370638.37349606, 1370638.37349606, 1370638.37349606, 
    1370638.37349606, 1370638.37349606, 1370638.37349606, 1370638.37349606, 
    1370638.37349606, 1370638.37349606, 1370638.37349606, 1370638.37349606, 
    1370638.37349606, 1370638.37349606, 1370638.37349606, 1370638.37349606, 
    1370638.37349606, 1370638.37349606, 1370638.37349606, 1370638.37349606, 
    1370638.37349606, 1370638.37349606, 1370638.37349606, 1370638.37349606, 
    1370638.37349606, 1370638.37349606, 1370638.37349606, 1370638.37349606, 
    1370638.37349606, 1370638.37349606, 1370638.37349606, 1370638.37349606, 
    1370638.37349606, 1370638.37349606, 1370638.37349606, 1370638.37349606, 
    1370638.37349606, 1370638.37349606, 1370638.37349606, 1370638.37349606, 
    1370638.37349606, 1370638.37349606, 1370638.37349606, 1370638.37349606, 
    1370638.37349606, 1370638.37349606, 1370638.37349606, 1370638.37349606, 
    1370638.37349606, 1370638.37349606, 1370638.37349606, 1370638.37349606, 
    1370638.37349606, 1370638.37349606, 1370638.37349606,
  1407682.65386082, 1407682.65386082, 1407682.65386082, 1407682.65386082, 
    1407682.65386082, 1407682.65386082, 1407682.65386082, 1407682.65386082, 
    1407682.65386082, 1407682.65386082, 1407682.65386082, 1407682.65386082, 
    1407682.65386082, 1407682.65386082, 1407682.65386082, 1407682.65386082, 
    1407682.65386082, 1407682.65386082, 1407682.65386082, 1407682.65386082, 
    1407682.65386082, 1407682.65386082, 1407682.65386082, 1407682.65386082, 
    1407682.65386082, 1407682.65386082, 1407682.65386082, 1407682.65386082, 
    1407682.65386082, 1407682.65386082, 1407682.65386082, 1407682.65386082, 
    1407682.65386082, 1407682.65386082, 1407682.65386082, 1407682.65386082, 
    1407682.65386082, 1407682.65386082, 1407682.65386082, 1407682.65386082, 
    1407682.65386082, 1407682.65386082, 1407682.65386082, 1407682.65386082, 
    1407682.65386082, 1407682.65386082, 1407682.65386082, 1407682.65386082, 
    1407682.65386082, 1407682.65386082, 1407682.65386082, 1407682.65386082, 
    1407682.65386082, 1407682.65386082, 1407682.65386082,
  1444726.93422558, 1444726.93422558, 1444726.93422558, 1444726.93422558, 
    1444726.93422558, 1444726.93422558, 1444726.93422558, 1444726.93422558, 
    1444726.93422558, 1444726.93422558, 1444726.93422558, 1444726.93422558, 
    1444726.93422558, 1444726.93422558, 1444726.93422558, 1444726.93422558, 
    1444726.93422558, 1444726.93422558, 1444726.93422558, 1444726.93422558, 
    1444726.93422558, 1444726.93422558, 1444726.93422558, 1444726.93422558, 
    1444726.93422558, 1444726.93422558, 1444726.93422558, 1444726.93422558, 
    1444726.93422558, 1444726.93422558, 1444726.93422558, 1444726.93422558, 
    1444726.93422558, 1444726.93422558, 1444726.93422558, 1444726.93422558, 
    1444726.93422558, 1444726.93422558, 1444726.93422558, 1444726.93422558, 
    1444726.93422558, 1444726.93422558, 1444726.93422558, 1444726.93422558, 
    1444726.93422558, 1444726.93422558, 1444726.93422558, 1444726.93422558, 
    1444726.93422558, 1444726.93422558, 1444726.93422558, 1444726.93422558, 
    1444726.93422558, 1444726.93422558, 1444726.93422558,
  1481771.21459033, 1481771.21459033, 1481771.21459033, 1481771.21459033, 
    1481771.21459033, 1481771.21459033, 1481771.21459033, 1481771.21459033, 
    1481771.21459033, 1481771.21459033, 1481771.21459033, 1481771.21459033, 
    1481771.21459033, 1481771.21459033, 1481771.21459033, 1481771.21459033, 
    1481771.21459033, 1481771.21459033, 1481771.21459033, 1481771.21459033, 
    1481771.21459033, 1481771.21459033, 1481771.21459033, 1481771.21459033, 
    1481771.21459033, 1481771.21459033, 1481771.21459033, 1481771.21459033, 
    1481771.21459033, 1481771.21459033, 1481771.21459033, 1481771.21459033, 
    1481771.21459033, 1481771.21459033, 1481771.21459033, 1481771.21459033, 
    1481771.21459033, 1481771.21459033, 1481771.21459033, 1481771.21459033, 
    1481771.21459033, 1481771.21459033, 1481771.21459033, 1481771.21459033, 
    1481771.21459033, 1481771.21459033, 1481771.21459033, 1481771.21459033, 
    1481771.21459033, 1481771.21459033, 1481771.21459033, 1481771.21459033, 
    1481771.21459033, 1481771.21459033, 1481771.21459033,
  1518815.49495509, 1518815.49495509, 1518815.49495509, 1518815.49495509, 
    1518815.49495509, 1518815.49495509, 1518815.49495509, 1518815.49495509, 
    1518815.49495509, 1518815.49495509, 1518815.49495509, 1518815.49495509, 
    1518815.49495509, 1518815.49495509, 1518815.49495509, 1518815.49495509, 
    1518815.49495509, 1518815.49495509, 1518815.49495509, 1518815.49495509, 
    1518815.49495509, 1518815.49495509, 1518815.49495509, 1518815.49495509, 
    1518815.49495509, 1518815.49495509, 1518815.49495509, 1518815.49495509, 
    1518815.49495509, 1518815.49495509, 1518815.49495509, 1518815.49495509, 
    1518815.49495509, 1518815.49495509, 1518815.49495509, 1518815.49495509, 
    1518815.49495509, 1518815.49495509, 1518815.49495509, 1518815.49495509, 
    1518815.49495509, 1518815.49495509, 1518815.49495509, 1518815.49495509, 
    1518815.49495509, 1518815.49495509, 1518815.49495509, 1518815.49495509, 
    1518815.49495509, 1518815.49495509, 1518815.49495509, 1518815.49495509, 
    1518815.49495509, 1518815.49495509, 1518815.49495509,
  1555859.77531985, 1555859.77531985, 1555859.77531985, 1555859.77531985, 
    1555859.77531985, 1555859.77531985, 1555859.77531985, 1555859.77531985, 
    1555859.77531985, 1555859.77531985, 1555859.77531985, 1555859.77531985, 
    1555859.77531985, 1555859.77531985, 1555859.77531985, 1555859.77531985, 
    1555859.77531985, 1555859.77531985, 1555859.77531985, 1555859.77531985, 
    1555859.77531985, 1555859.77531985, 1555859.77531985, 1555859.77531985, 
    1555859.77531985, 1555859.77531985, 1555859.77531985, 1555859.77531985, 
    1555859.77531985, 1555859.77531985, 1555859.77531985, 1555859.77531985, 
    1555859.77531985, 1555859.77531985, 1555859.77531985, 1555859.77531985, 
    1555859.77531985, 1555859.77531985, 1555859.77531985, 1555859.77531985, 
    1555859.77531985, 1555859.77531985, 1555859.77531985, 1555859.77531985, 
    1555859.77531985, 1555859.77531985, 1555859.77531985, 1555859.77531985, 
    1555859.77531985, 1555859.77531985, 1555859.77531985, 1555859.77531985, 
    1555859.77531985, 1555859.77531985, 1555859.77531985,
  1592904.05568461, 1592904.05568461, 1592904.05568461, 1592904.05568461, 
    1592904.05568461, 1592904.05568461, 1592904.05568461, 1592904.05568461, 
    1592904.05568461, 1592904.05568461, 1592904.05568461, 1592904.05568461, 
    1592904.05568461, 1592904.05568461, 1592904.05568461, 1592904.05568461, 
    1592904.05568461, 1592904.05568461, 1592904.05568461, 1592904.05568461, 
    1592904.05568461, 1592904.05568461, 1592904.05568461, 1592904.05568461, 
    1592904.05568461, 1592904.05568461, 1592904.05568461, 1592904.05568461, 
    1592904.05568461, 1592904.05568461, 1592904.05568461, 1592904.05568461, 
    1592904.05568461, 1592904.05568461, 1592904.05568461, 1592904.05568461, 
    1592904.05568461, 1592904.05568461, 1592904.05568461, 1592904.05568461, 
    1592904.05568461, 1592904.05568461, 1592904.05568461, 1592904.05568461, 
    1592904.05568461, 1592904.05568461, 1592904.05568461, 1592904.05568461, 
    1592904.05568461, 1592904.05568461, 1592904.05568461, 1592904.05568461, 
    1592904.05568461, 1592904.05568461, 1592904.05568461,
  1629948.33604937, 1629948.33604937, 1629948.33604937, 1629948.33604937, 
    1629948.33604937, 1629948.33604937, 1629948.33604937, 1629948.33604937, 
    1629948.33604937, 1629948.33604937, 1629948.33604937, 1629948.33604937, 
    1629948.33604937, 1629948.33604937, 1629948.33604937, 1629948.33604937, 
    1629948.33604937, 1629948.33604937, 1629948.33604937, 1629948.33604937, 
    1629948.33604937, 1629948.33604937, 1629948.33604937, 1629948.33604937, 
    1629948.33604937, 1629948.33604937, 1629948.33604937, 1629948.33604937, 
    1629948.33604937, 1629948.33604937, 1629948.33604937, 1629948.33604937, 
    1629948.33604937, 1629948.33604937, 1629948.33604937, 1629948.33604937, 
    1629948.33604937, 1629948.33604937, 1629948.33604937, 1629948.33604937, 
    1629948.33604937, 1629948.33604937, 1629948.33604937, 1629948.33604937, 
    1629948.33604937, 1629948.33604937, 1629948.33604937, 1629948.33604937, 
    1629948.33604937, 1629948.33604937, 1629948.33604937, 1629948.33604937, 
    1629948.33604937, 1629948.33604937, 1629948.33604937,
  1666992.61641413, 1666992.61641413, 1666992.61641413, 1666992.61641413, 
    1666992.61641413, 1666992.61641413, 1666992.61641413, 1666992.61641413, 
    1666992.61641413, 1666992.61641413, 1666992.61641413, 1666992.61641413, 
    1666992.61641413, 1666992.61641413, 1666992.61641413, 1666992.61641413, 
    1666992.61641413, 1666992.61641413, 1666992.61641413, 1666992.61641413, 
    1666992.61641413, 1666992.61641413, 1666992.61641413, 1666992.61641413, 
    1666992.61641413, 1666992.61641413, 1666992.61641413, 1666992.61641413, 
    1666992.61641413, 1666992.61641413, 1666992.61641413, 1666992.61641413, 
    1666992.61641413, 1666992.61641413, 1666992.61641413, 1666992.61641413, 
    1666992.61641413, 1666992.61641413, 1666992.61641413, 1666992.61641413, 
    1666992.61641413, 1666992.61641413, 1666992.61641413, 1666992.61641413, 
    1666992.61641413, 1666992.61641413, 1666992.61641413, 1666992.61641413, 
    1666992.61641413, 1666992.61641413, 1666992.61641413, 1666992.61641413, 
    1666992.61641413, 1666992.61641413, 1666992.61641413,
  1704036.89677889, 1704036.89677889, 1704036.89677889, 1704036.89677889, 
    1704036.89677889, 1704036.89677889, 1704036.89677889, 1704036.89677889, 
    1704036.89677889, 1704036.89677889, 1704036.89677889, 1704036.89677889, 
    1704036.89677889, 1704036.89677889, 1704036.89677889, 1704036.89677889, 
    1704036.89677889, 1704036.89677889, 1704036.89677889, 1704036.89677889, 
    1704036.89677889, 1704036.89677889, 1704036.89677889, 1704036.89677889, 
    1704036.89677889, 1704036.89677889, 1704036.89677889, 1704036.89677889, 
    1704036.89677889, 1704036.89677889, 1704036.89677889, 1704036.89677889, 
    1704036.89677889, 1704036.89677889, 1704036.89677889, 1704036.89677889, 
    1704036.89677889, 1704036.89677889, 1704036.89677889, 1704036.89677889, 
    1704036.89677889, 1704036.89677889, 1704036.89677889, 1704036.89677889, 
    1704036.89677889, 1704036.89677889, 1704036.89677889, 1704036.89677889, 
    1704036.89677889, 1704036.89677889, 1704036.89677889, 1704036.89677889, 
    1704036.89677889, 1704036.89677889, 1704036.89677889,
  1741081.17714364, 1741081.17714364, 1741081.17714364, 1741081.17714364, 
    1741081.17714364, 1741081.17714364, 1741081.17714364, 1741081.17714364, 
    1741081.17714364, 1741081.17714364, 1741081.17714364, 1741081.17714364, 
    1741081.17714364, 1741081.17714364, 1741081.17714364, 1741081.17714364, 
    1741081.17714364, 1741081.17714364, 1741081.17714364, 1741081.17714364, 
    1741081.17714364, 1741081.17714364, 1741081.17714364, 1741081.17714364, 
    1741081.17714364, 1741081.17714364, 1741081.17714364, 1741081.17714364, 
    1741081.17714364, 1741081.17714364, 1741081.17714364, 1741081.17714364, 
    1741081.17714364, 1741081.17714364, 1741081.17714364, 1741081.17714364, 
    1741081.17714364, 1741081.17714364, 1741081.17714364, 1741081.17714364, 
    1741081.17714364, 1741081.17714364, 1741081.17714364, 1741081.17714364, 
    1741081.17714364, 1741081.17714364, 1741081.17714364, 1741081.17714364, 
    1741081.17714364, 1741081.17714364, 1741081.17714364, 1741081.17714364, 
    1741081.17714364, 1741081.17714364, 1741081.17714364,
  1778125.4575084, 1778125.4575084, 1778125.4575084, 1778125.4575084, 
    1778125.4575084, 1778125.4575084, 1778125.4575084, 1778125.4575084, 
    1778125.4575084, 1778125.4575084, 1778125.4575084, 1778125.4575084, 
    1778125.4575084, 1778125.4575084, 1778125.4575084, 1778125.4575084, 
    1778125.4575084, 1778125.4575084, 1778125.4575084, 1778125.4575084, 
    1778125.4575084, 1778125.4575084, 1778125.4575084, 1778125.4575084, 
    1778125.4575084, 1778125.4575084, 1778125.4575084, 1778125.4575084, 
    1778125.4575084, 1778125.4575084, 1778125.4575084, 1778125.4575084, 
    1778125.4575084, 1778125.4575084, 1778125.4575084, 1778125.4575084, 
    1778125.4575084, 1778125.4575084, 1778125.4575084, 1778125.4575084, 
    1778125.4575084, 1778125.4575084, 1778125.4575084, 1778125.4575084, 
    1778125.4575084, 1778125.4575084, 1778125.4575084, 1778125.4575084, 
    1778125.4575084, 1778125.4575084, 1778125.4575084, 1778125.4575084, 
    1778125.4575084, 1778125.4575084, 1778125.4575084,
  1815169.73787316, 1815169.73787316, 1815169.73787316, 1815169.73787316, 
    1815169.73787316, 1815169.73787316, 1815169.73787316, 1815169.73787316, 
    1815169.73787316, 1815169.73787316, 1815169.73787316, 1815169.73787316, 
    1815169.73787316, 1815169.73787316, 1815169.73787316, 1815169.73787316, 
    1815169.73787316, 1815169.73787316, 1815169.73787316, 1815169.73787316, 
    1815169.73787316, 1815169.73787316, 1815169.73787316, 1815169.73787316, 
    1815169.73787316, 1815169.73787316, 1815169.73787316, 1815169.73787316, 
    1815169.73787316, 1815169.73787316, 1815169.73787316, 1815169.73787316, 
    1815169.73787316, 1815169.73787316, 1815169.73787316, 1815169.73787316, 
    1815169.73787316, 1815169.73787316, 1815169.73787316, 1815169.73787316, 
    1815169.73787316, 1815169.73787316, 1815169.73787316, 1815169.73787316, 
    1815169.73787316, 1815169.73787316, 1815169.73787316, 1815169.73787316, 
    1815169.73787316, 1815169.73787316, 1815169.73787316, 1815169.73787316, 
    1815169.73787316, 1815169.73787316, 1815169.73787316,
  1852214.01823792, 1852214.01823792, 1852214.01823792, 1852214.01823792, 
    1852214.01823792, 1852214.01823792, 1852214.01823792, 1852214.01823792, 
    1852214.01823792, 1852214.01823792, 1852214.01823792, 1852214.01823792, 
    1852214.01823792, 1852214.01823792, 1852214.01823792, 1852214.01823792, 
    1852214.01823792, 1852214.01823792, 1852214.01823792, 1852214.01823792, 
    1852214.01823792, 1852214.01823792, 1852214.01823792, 1852214.01823792, 
    1852214.01823792, 1852214.01823792, 1852214.01823792, 1852214.01823792, 
    1852214.01823792, 1852214.01823792, 1852214.01823792, 1852214.01823792, 
    1852214.01823792, 1852214.01823792, 1852214.01823792, 1852214.01823792, 
    1852214.01823792, 1852214.01823792, 1852214.01823792, 1852214.01823792, 
    1852214.01823792, 1852214.01823792, 1852214.01823792, 1852214.01823792, 
    1852214.01823792, 1852214.01823792, 1852214.01823792, 1852214.01823792, 
    1852214.01823792, 1852214.01823792, 1852214.01823792, 1852214.01823792, 
    1852214.01823792, 1852214.01823792, 1852214.01823792,
  1889258.29860268, 1889258.29860268, 1889258.29860268, 1889258.29860268, 
    1889258.29860268, 1889258.29860268, 1889258.29860268, 1889258.29860268, 
    1889258.29860268, 1889258.29860268, 1889258.29860268, 1889258.29860268, 
    1889258.29860268, 1889258.29860268, 1889258.29860268, 1889258.29860268, 
    1889258.29860268, 1889258.29860268, 1889258.29860268, 1889258.29860268, 
    1889258.29860268, 1889258.29860268, 1889258.29860268, 1889258.29860268, 
    1889258.29860268, 1889258.29860268, 1889258.29860268, 1889258.29860268, 
    1889258.29860268, 1889258.29860268, 1889258.29860268, 1889258.29860268, 
    1889258.29860268, 1889258.29860268, 1889258.29860268, 1889258.29860268, 
    1889258.29860268, 1889258.29860268, 1889258.29860268, 1889258.29860268, 
    1889258.29860268, 1889258.29860268, 1889258.29860268, 1889258.29860268, 
    1889258.29860268, 1889258.29860268, 1889258.29860268, 1889258.29860268, 
    1889258.29860268, 1889258.29860268, 1889258.29860268, 1889258.29860268, 
    1889258.29860268, 1889258.29860268, 1889258.29860268,
  1926302.57896744, 1926302.57896744, 1926302.57896744, 1926302.57896744, 
    1926302.57896744, 1926302.57896744, 1926302.57896744, 1926302.57896744, 
    1926302.57896744, 1926302.57896744, 1926302.57896744, 1926302.57896744, 
    1926302.57896744, 1926302.57896744, 1926302.57896744, 1926302.57896744, 
    1926302.57896744, 1926302.57896744, 1926302.57896744, 1926302.57896744, 
    1926302.57896744, 1926302.57896744, 1926302.57896744, 1926302.57896744, 
    1926302.57896744, 1926302.57896744, 1926302.57896744, 1926302.57896744, 
    1926302.57896744, 1926302.57896744, 1926302.57896744, 1926302.57896744, 
    1926302.57896744, 1926302.57896744, 1926302.57896744, 1926302.57896744, 
    1926302.57896744, 1926302.57896744, 1926302.57896744, 1926302.57896744, 
    1926302.57896744, 1926302.57896744, 1926302.57896744, 1926302.57896744, 
    1926302.57896744, 1926302.57896744, 1926302.57896744, 1926302.57896744, 
    1926302.57896744, 1926302.57896744, 1926302.57896744, 1926302.57896744, 
    1926302.57896744, 1926302.57896744, 1926302.57896744,
  1963346.85933219, 1963346.85933219, 1963346.85933219, 1963346.85933219, 
    1963346.85933219, 1963346.85933219, 1963346.85933219, 1963346.85933219, 
    1963346.85933219, 1963346.85933219, 1963346.85933219, 1963346.85933219, 
    1963346.85933219, 1963346.85933219, 1963346.85933219, 1963346.85933219, 
    1963346.85933219, 1963346.85933219, 1963346.85933219, 1963346.85933219, 
    1963346.85933219, 1963346.85933219, 1963346.85933219, 1963346.85933219, 
    1963346.85933219, 1963346.85933219, 1963346.85933219, 1963346.85933219, 
    1963346.85933219, 1963346.85933219, 1963346.85933219, 1963346.85933219, 
    1963346.85933219, 1963346.85933219, 1963346.85933219, 1963346.85933219, 
    1963346.85933219, 1963346.85933219, 1963346.85933219, 1963346.85933219, 
    1963346.85933219, 1963346.85933219, 1963346.85933219, 1963346.85933219, 
    1963346.85933219, 1963346.85933219, 1963346.85933219, 1963346.85933219, 
    1963346.85933219, 1963346.85933219, 1963346.85933219, 1963346.85933219, 
    1963346.85933219, 1963346.85933219, 1963346.85933219,
  2000391.13969695, 2000391.13969695, 2000391.13969695, 2000391.13969695, 
    2000391.13969695, 2000391.13969695, 2000391.13969695, 2000391.13969695, 
    2000391.13969695, 2000391.13969695, 2000391.13969695, 2000391.13969695, 
    2000391.13969695, 2000391.13969695, 2000391.13969695, 2000391.13969695, 
    2000391.13969695, 2000391.13969695, 2000391.13969695, 2000391.13969695, 
    2000391.13969695, 2000391.13969695, 2000391.13969695, 2000391.13969695, 
    2000391.13969695, 2000391.13969695, 2000391.13969695, 2000391.13969695, 
    2000391.13969695, 2000391.13969695, 2000391.13969695, 2000391.13969695, 
    2000391.13969695, 2000391.13969695, 2000391.13969695, 2000391.13969695, 
    2000391.13969695, 2000391.13969695, 2000391.13969695, 2000391.13969695, 
    2000391.13969695, 2000391.13969695, 2000391.13969695, 2000391.13969695, 
    2000391.13969695, 2000391.13969695, 2000391.13969695, 2000391.13969695, 
    2000391.13969695, 2000391.13969695, 2000391.13969695, 2000391.13969695, 
    2000391.13969695, 2000391.13969695, 2000391.13969695 ;

 y_v =
  18522.1401823791, 18522.1401823791, 18522.1401823791, 18522.1401823791, 
    18522.1401823791, 18522.1401823791, 18522.1401823791, 18522.1401823791, 
    18522.1401823791, 18522.1401823791, 18522.1401823791, 18522.1401823791, 
    18522.1401823791, 18522.1401823791, 18522.1401823791, 18522.1401823791, 
    18522.1401823791, 18522.1401823791, 18522.1401823791, 18522.1401823791, 
    18522.1401823791, 18522.1401823791, 18522.1401823791, 18522.1401823791, 
    18522.1401823791, 18522.1401823791, 18522.1401823791, 18522.1401823791, 
    18522.1401823791, 18522.1401823791, 18522.1401823791, 18522.1401823791, 
    18522.1401823791, 18522.1401823791, 18522.1401823791, 18522.1401823791, 
    18522.1401823791, 18522.1401823791, 18522.1401823791, 18522.1401823791, 
    18522.1401823791, 18522.1401823791, 18522.1401823791, 18522.1401823791, 
    18522.1401823791, 18522.1401823791, 18522.1401823791, 18522.1401823791, 
    18522.1401823791, 18522.1401823791, 18522.1401823791, 18522.1401823791, 
    18522.1401823791, 18522.1401823791, 18522.1401823791, 18522.1401823791,
  55566.4205471374, 55566.4205471374, 55566.4205471374, 55566.4205471374, 
    55566.4205471374, 55566.4205471374, 55566.4205471374, 55566.4205471374, 
    55566.4205471374, 55566.4205471374, 55566.4205471374, 55566.4205471374, 
    55566.4205471374, 55566.4205471374, 55566.4205471374, 55566.4205471374, 
    55566.4205471374, 55566.4205471374, 55566.4205471374, 55566.4205471374, 
    55566.4205471374, 55566.4205471374, 55566.4205471374, 55566.4205471374, 
    55566.4205471374, 55566.4205471374, 55566.4205471374, 55566.4205471374, 
    55566.4205471374, 55566.4205471374, 55566.4205471374, 55566.4205471374, 
    55566.4205471374, 55566.4205471374, 55566.4205471374, 55566.4205471374, 
    55566.4205471374, 55566.4205471374, 55566.4205471374, 55566.4205471374, 
    55566.4205471374, 55566.4205471374, 55566.4205471374, 55566.4205471374, 
    55566.4205471374, 55566.4205471374, 55566.4205471374, 55566.4205471374, 
    55566.4205471374, 55566.4205471374, 55566.4205471374, 55566.4205471374, 
    55566.4205471374, 55566.4205471374, 55566.4205471374, 55566.4205471374,
  92610.7009118959, 92610.7009118959, 92610.7009118959, 92610.7009118959, 
    92610.7009118959, 92610.7009118959, 92610.7009118959, 92610.7009118959, 
    92610.7009118959, 92610.7009118959, 92610.7009118959, 92610.7009118959, 
    92610.7009118959, 92610.7009118959, 92610.7009118959, 92610.7009118959, 
    92610.7009118959, 92610.7009118959, 92610.7009118959, 92610.7009118959, 
    92610.7009118959, 92610.7009118959, 92610.7009118959, 92610.7009118959, 
    92610.7009118959, 92610.7009118959, 92610.7009118959, 92610.7009118959, 
    92610.7009118959, 92610.7009118959, 92610.7009118959, 92610.7009118959, 
    92610.7009118959, 92610.7009118959, 92610.7009118959, 92610.7009118959, 
    92610.7009118959, 92610.7009118959, 92610.7009118959, 92610.7009118959, 
    92610.7009118959, 92610.7009118959, 92610.7009118959, 92610.7009118959, 
    92610.7009118959, 92610.7009118959, 92610.7009118959, 92610.7009118959, 
    92610.7009118959, 92610.7009118959, 92610.7009118959, 92610.7009118959, 
    92610.7009118959, 92610.7009118959, 92610.7009118959, 92610.7009118959,
  129654.981276654, 129654.981276654, 129654.981276654, 129654.981276654, 
    129654.981276654, 129654.981276654, 129654.981276654, 129654.981276654, 
    129654.981276654, 129654.981276654, 129654.981276654, 129654.981276654, 
    129654.981276654, 129654.981276654, 129654.981276654, 129654.981276654, 
    129654.981276654, 129654.981276654, 129654.981276654, 129654.981276654, 
    129654.981276654, 129654.981276654, 129654.981276654, 129654.981276654, 
    129654.981276654, 129654.981276654, 129654.981276654, 129654.981276654, 
    129654.981276654, 129654.981276654, 129654.981276654, 129654.981276654, 
    129654.981276654, 129654.981276654, 129654.981276654, 129654.981276654, 
    129654.981276654, 129654.981276654, 129654.981276654, 129654.981276654, 
    129654.981276654, 129654.981276654, 129654.981276654, 129654.981276654, 
    129654.981276654, 129654.981276654, 129654.981276654, 129654.981276654, 
    129654.981276654, 129654.981276654, 129654.981276654, 129654.981276654, 
    129654.981276654, 129654.981276654, 129654.981276654, 129654.981276654,
  166699.261641412, 166699.261641412, 166699.261641412, 166699.261641412, 
    166699.261641412, 166699.261641412, 166699.261641412, 166699.261641412, 
    166699.261641412, 166699.261641412, 166699.261641412, 166699.261641412, 
    166699.261641412, 166699.261641412, 166699.261641412, 166699.261641412, 
    166699.261641412, 166699.261641412, 166699.261641412, 166699.261641412, 
    166699.261641412, 166699.261641412, 166699.261641412, 166699.261641412, 
    166699.261641412, 166699.261641412, 166699.261641412, 166699.261641412, 
    166699.261641412, 166699.261641412, 166699.261641412, 166699.261641412, 
    166699.261641412, 166699.261641412, 166699.261641412, 166699.261641412, 
    166699.261641412, 166699.261641412, 166699.261641412, 166699.261641412, 
    166699.261641412, 166699.261641412, 166699.261641412, 166699.261641412, 
    166699.261641412, 166699.261641412, 166699.261641412, 166699.261641412, 
    166699.261641412, 166699.261641412, 166699.261641412, 166699.261641412, 
    166699.261641412, 166699.261641412, 166699.261641412, 166699.261641412,
  203743.542006171, 203743.542006171, 203743.542006171, 203743.542006171, 
    203743.542006171, 203743.542006171, 203743.542006171, 203743.542006171, 
    203743.542006171, 203743.542006171, 203743.542006171, 203743.542006171, 
    203743.542006171, 203743.542006171, 203743.542006171, 203743.542006171, 
    203743.542006171, 203743.542006171, 203743.542006171, 203743.542006171, 
    203743.542006171, 203743.542006171, 203743.542006171, 203743.542006171, 
    203743.542006171, 203743.542006171, 203743.542006171, 203743.542006171, 
    203743.542006171, 203743.542006171, 203743.542006171, 203743.542006171, 
    203743.542006171, 203743.542006171, 203743.542006171, 203743.542006171, 
    203743.542006171, 203743.542006171, 203743.542006171, 203743.542006171, 
    203743.542006171, 203743.542006171, 203743.542006171, 203743.542006171, 
    203743.542006171, 203743.542006171, 203743.542006171, 203743.542006171, 
    203743.542006171, 203743.542006171, 203743.542006171, 203743.542006171, 
    203743.542006171, 203743.542006171, 203743.542006171, 203743.542006171,
  240787.82237093, 240787.82237093, 240787.82237093, 240787.82237093, 
    240787.82237093, 240787.82237093, 240787.82237093, 240787.82237093, 
    240787.82237093, 240787.82237093, 240787.82237093, 240787.82237093, 
    240787.82237093, 240787.82237093, 240787.82237093, 240787.82237093, 
    240787.82237093, 240787.82237093, 240787.82237093, 240787.82237093, 
    240787.82237093, 240787.82237093, 240787.82237093, 240787.82237093, 
    240787.82237093, 240787.82237093, 240787.82237093, 240787.82237093, 
    240787.82237093, 240787.82237093, 240787.82237093, 240787.82237093, 
    240787.82237093, 240787.82237093, 240787.82237093, 240787.82237093, 
    240787.82237093, 240787.82237093, 240787.82237093, 240787.82237093, 
    240787.82237093, 240787.82237093, 240787.82237093, 240787.82237093, 
    240787.82237093, 240787.82237093, 240787.82237093, 240787.82237093, 
    240787.82237093, 240787.82237093, 240787.82237093, 240787.82237093, 
    240787.82237093, 240787.82237093, 240787.82237093, 240787.82237093,
  277832.102735688, 277832.102735688, 277832.102735688, 277832.102735688, 
    277832.102735688, 277832.102735688, 277832.102735688, 277832.102735688, 
    277832.102735688, 277832.102735688, 277832.102735688, 277832.102735688, 
    277832.102735688, 277832.102735688, 277832.102735688, 277832.102735688, 
    277832.102735688, 277832.102735688, 277832.102735688, 277832.102735688, 
    277832.102735688, 277832.102735688, 277832.102735688, 277832.102735688, 
    277832.102735688, 277832.102735688, 277832.102735688, 277832.102735688, 
    277832.102735688, 277832.102735688, 277832.102735688, 277832.102735688, 
    277832.102735688, 277832.102735688, 277832.102735688, 277832.102735688, 
    277832.102735688, 277832.102735688, 277832.102735688, 277832.102735688, 
    277832.102735688, 277832.102735688, 277832.102735688, 277832.102735688, 
    277832.102735688, 277832.102735688, 277832.102735688, 277832.102735688, 
    277832.102735688, 277832.102735688, 277832.102735688, 277832.102735688, 
    277832.102735688, 277832.102735688, 277832.102735688, 277832.102735688,
  314876.383100447, 314876.383100447, 314876.383100447, 314876.383100447, 
    314876.383100447, 314876.383100447, 314876.383100447, 314876.383100447, 
    314876.383100447, 314876.383100447, 314876.383100447, 314876.383100447, 
    314876.383100447, 314876.383100447, 314876.383100447, 314876.383100447, 
    314876.383100447, 314876.383100447, 314876.383100447, 314876.383100447, 
    314876.383100447, 314876.383100447, 314876.383100447, 314876.383100447, 
    314876.383100447, 314876.383100447, 314876.383100447, 314876.383100447, 
    314876.383100447, 314876.383100447, 314876.383100447, 314876.383100447, 
    314876.383100447, 314876.383100447, 314876.383100447, 314876.383100447, 
    314876.383100447, 314876.383100447, 314876.383100447, 314876.383100447, 
    314876.383100447, 314876.383100447, 314876.383100447, 314876.383100447, 
    314876.383100447, 314876.383100447, 314876.383100447, 314876.383100447, 
    314876.383100447, 314876.383100447, 314876.383100447, 314876.383100447, 
    314876.383100447, 314876.383100447, 314876.383100447, 314876.383100447,
  351920.663465205, 351920.663465205, 351920.663465205, 351920.663465205, 
    351920.663465205, 351920.663465205, 351920.663465205, 351920.663465205, 
    351920.663465205, 351920.663465205, 351920.663465205, 351920.663465205, 
    351920.663465205, 351920.663465205, 351920.663465205, 351920.663465205, 
    351920.663465205, 351920.663465205, 351920.663465205, 351920.663465205, 
    351920.663465205, 351920.663465205, 351920.663465205, 351920.663465205, 
    351920.663465205, 351920.663465205, 351920.663465205, 351920.663465205, 
    351920.663465205, 351920.663465205, 351920.663465205, 351920.663465205, 
    351920.663465205, 351920.663465205, 351920.663465205, 351920.663465205, 
    351920.663465205, 351920.663465205, 351920.663465205, 351920.663465205, 
    351920.663465205, 351920.663465205, 351920.663465205, 351920.663465205, 
    351920.663465205, 351920.663465205, 351920.663465205, 351920.663465205, 
    351920.663465205, 351920.663465205, 351920.663465205, 351920.663465205, 
    351920.663465205, 351920.663465205, 351920.663465205, 351920.663465205,
  388964.943829963, 388964.943829963, 388964.943829963, 388964.943829963, 
    388964.943829963, 388964.943829963, 388964.943829963, 388964.943829963, 
    388964.943829963, 388964.943829963, 388964.943829963, 388964.943829963, 
    388964.943829963, 388964.943829963, 388964.943829963, 388964.943829963, 
    388964.943829963, 388964.943829963, 388964.943829963, 388964.943829963, 
    388964.943829963, 388964.943829963, 388964.943829963, 388964.943829963, 
    388964.943829963, 388964.943829963, 388964.943829963, 388964.943829963, 
    388964.943829963, 388964.943829963, 388964.943829963, 388964.943829963, 
    388964.943829963, 388964.943829963, 388964.943829963, 388964.943829963, 
    388964.943829963, 388964.943829963, 388964.943829963, 388964.943829963, 
    388964.943829963, 388964.943829963, 388964.943829963, 388964.943829963, 
    388964.943829963, 388964.943829963, 388964.943829963, 388964.943829963, 
    388964.943829963, 388964.943829963, 388964.943829963, 388964.943829963, 
    388964.943829963, 388964.943829963, 388964.943829963, 388964.943829963,
  426009.224194721, 426009.224194721, 426009.224194721, 426009.224194721, 
    426009.224194721, 426009.224194721, 426009.224194721, 426009.224194721, 
    426009.224194721, 426009.224194721, 426009.224194721, 426009.224194721, 
    426009.224194721, 426009.224194721, 426009.224194721, 426009.224194721, 
    426009.224194721, 426009.224194721, 426009.224194721, 426009.224194721, 
    426009.224194721, 426009.224194721, 426009.224194721, 426009.224194721, 
    426009.224194721, 426009.224194721, 426009.224194721, 426009.224194721, 
    426009.224194721, 426009.224194721, 426009.224194721, 426009.224194721, 
    426009.224194721, 426009.224194721, 426009.224194721, 426009.224194721, 
    426009.224194721, 426009.224194721, 426009.224194721, 426009.224194721, 
    426009.224194721, 426009.224194721, 426009.224194721, 426009.224194721, 
    426009.224194721, 426009.224194721, 426009.224194721, 426009.224194721, 
    426009.224194721, 426009.224194721, 426009.224194721, 426009.224194721, 
    426009.224194721, 426009.224194721, 426009.224194721, 426009.224194721,
  463053.50455948, 463053.50455948, 463053.50455948, 463053.50455948, 
    463053.50455948, 463053.50455948, 463053.50455948, 463053.50455948, 
    463053.50455948, 463053.50455948, 463053.50455948, 463053.50455948, 
    463053.50455948, 463053.50455948, 463053.50455948, 463053.50455948, 
    463053.50455948, 463053.50455948, 463053.50455948, 463053.50455948, 
    463053.50455948, 463053.50455948, 463053.50455948, 463053.50455948, 
    463053.50455948, 463053.50455948, 463053.50455948, 463053.50455948, 
    463053.50455948, 463053.50455948, 463053.50455948, 463053.50455948, 
    463053.50455948, 463053.50455948, 463053.50455948, 463053.50455948, 
    463053.50455948, 463053.50455948, 463053.50455948, 463053.50455948, 
    463053.50455948, 463053.50455948, 463053.50455948, 463053.50455948, 
    463053.50455948, 463053.50455948, 463053.50455948, 463053.50455948, 
    463053.50455948, 463053.50455948, 463053.50455948, 463053.50455948, 
    463053.50455948, 463053.50455948, 463053.50455948, 463053.50455948,
  500097.784924238, 500097.784924238, 500097.784924238, 500097.784924238, 
    500097.784924238, 500097.784924238, 500097.784924238, 500097.784924238, 
    500097.784924238, 500097.784924238, 500097.784924238, 500097.784924238, 
    500097.784924238, 500097.784924238, 500097.784924238, 500097.784924238, 
    500097.784924238, 500097.784924238, 500097.784924238, 500097.784924238, 
    500097.784924238, 500097.784924238, 500097.784924238, 500097.784924238, 
    500097.784924238, 500097.784924238, 500097.784924238, 500097.784924238, 
    500097.784924238, 500097.784924238, 500097.784924238, 500097.784924238, 
    500097.784924238, 500097.784924238, 500097.784924238, 500097.784924238, 
    500097.784924238, 500097.784924238, 500097.784924238, 500097.784924238, 
    500097.784924238, 500097.784924238, 500097.784924238, 500097.784924238, 
    500097.784924238, 500097.784924238, 500097.784924238, 500097.784924238, 
    500097.784924238, 500097.784924238, 500097.784924238, 500097.784924238, 
    500097.784924238, 500097.784924238, 500097.784924238, 500097.784924238,
  537142.065288996, 537142.065288996, 537142.065288996, 537142.065288996, 
    537142.065288996, 537142.065288996, 537142.065288996, 537142.065288996, 
    537142.065288996, 537142.065288996, 537142.065288996, 537142.065288996, 
    537142.065288996, 537142.065288996, 537142.065288996, 537142.065288996, 
    537142.065288996, 537142.065288996, 537142.065288996, 537142.065288996, 
    537142.065288996, 537142.065288996, 537142.065288996, 537142.065288996, 
    537142.065288996, 537142.065288996, 537142.065288996, 537142.065288996, 
    537142.065288996, 537142.065288996, 537142.065288996, 537142.065288996, 
    537142.065288996, 537142.065288996, 537142.065288996, 537142.065288996, 
    537142.065288996, 537142.065288996, 537142.065288996, 537142.065288996, 
    537142.065288996, 537142.065288996, 537142.065288996, 537142.065288996, 
    537142.065288996, 537142.065288996, 537142.065288996, 537142.065288996, 
    537142.065288996, 537142.065288996, 537142.065288996, 537142.065288996, 
    537142.065288996, 537142.065288996, 537142.065288996, 537142.065288996,
  574186.345653754, 574186.345653754, 574186.345653754, 574186.345653754, 
    574186.345653754, 574186.345653754, 574186.345653754, 574186.345653754, 
    574186.345653754, 574186.345653754, 574186.345653754, 574186.345653754, 
    574186.345653754, 574186.345653754, 574186.345653754, 574186.345653754, 
    574186.345653754, 574186.345653754, 574186.345653754, 574186.345653754, 
    574186.345653754, 574186.345653754, 574186.345653754, 574186.345653754, 
    574186.345653754, 574186.345653754, 574186.345653754, 574186.345653754, 
    574186.345653754, 574186.345653754, 574186.345653754, 574186.345653754, 
    574186.345653754, 574186.345653754, 574186.345653754, 574186.345653754, 
    574186.345653754, 574186.345653754, 574186.345653754, 574186.345653754, 
    574186.345653754, 574186.345653754, 574186.345653754, 574186.345653754, 
    574186.345653754, 574186.345653754, 574186.345653754, 574186.345653754, 
    574186.345653754, 574186.345653754, 574186.345653754, 574186.345653754, 
    574186.345653754, 574186.345653754, 574186.345653754, 574186.345653754,
  611230.626018513, 611230.626018513, 611230.626018513, 611230.626018513, 
    611230.626018513, 611230.626018513, 611230.626018513, 611230.626018513, 
    611230.626018513, 611230.626018513, 611230.626018513, 611230.626018513, 
    611230.626018513, 611230.626018513, 611230.626018513, 611230.626018513, 
    611230.626018513, 611230.626018513, 611230.626018513, 611230.626018513, 
    611230.626018513, 611230.626018513, 611230.626018513, 611230.626018513, 
    611230.626018513, 611230.626018513, 611230.626018513, 611230.626018513, 
    611230.626018513, 611230.626018513, 611230.626018513, 611230.626018513, 
    611230.626018513, 611230.626018513, 611230.626018513, 611230.626018513, 
    611230.626018513, 611230.626018513, 611230.626018513, 611230.626018513, 
    611230.626018513, 611230.626018513, 611230.626018513, 611230.626018513, 
    611230.626018513, 611230.626018513, 611230.626018513, 611230.626018513, 
    611230.626018513, 611230.626018513, 611230.626018513, 611230.626018513, 
    611230.626018513, 611230.626018513, 611230.626018513, 611230.626018513,
  648274.906383271, 648274.906383271, 648274.906383271, 648274.906383271, 
    648274.906383271, 648274.906383271, 648274.906383271, 648274.906383271, 
    648274.906383271, 648274.906383271, 648274.906383271, 648274.906383271, 
    648274.906383271, 648274.906383271, 648274.906383271, 648274.906383271, 
    648274.906383271, 648274.906383271, 648274.906383271, 648274.906383271, 
    648274.906383271, 648274.906383271, 648274.906383271, 648274.906383271, 
    648274.906383271, 648274.906383271, 648274.906383271, 648274.906383271, 
    648274.906383271, 648274.906383271, 648274.906383271, 648274.906383271, 
    648274.906383271, 648274.906383271, 648274.906383271, 648274.906383271, 
    648274.906383271, 648274.906383271, 648274.906383271, 648274.906383271, 
    648274.906383271, 648274.906383271, 648274.906383271, 648274.906383271, 
    648274.906383271, 648274.906383271, 648274.906383271, 648274.906383271, 
    648274.906383271, 648274.906383271, 648274.906383271, 648274.906383271, 
    648274.906383271, 648274.906383271, 648274.906383271, 648274.906383271,
  685319.18674803, 685319.18674803, 685319.18674803, 685319.18674803, 
    685319.18674803, 685319.18674803, 685319.18674803, 685319.18674803, 
    685319.18674803, 685319.18674803, 685319.18674803, 685319.18674803, 
    685319.18674803, 685319.18674803, 685319.18674803, 685319.18674803, 
    685319.18674803, 685319.18674803, 685319.18674803, 685319.18674803, 
    685319.18674803, 685319.18674803, 685319.18674803, 685319.18674803, 
    685319.18674803, 685319.18674803, 685319.18674803, 685319.18674803, 
    685319.18674803, 685319.18674803, 685319.18674803, 685319.18674803, 
    685319.18674803, 685319.18674803, 685319.18674803, 685319.18674803, 
    685319.18674803, 685319.18674803, 685319.18674803, 685319.18674803, 
    685319.18674803, 685319.18674803, 685319.18674803, 685319.18674803, 
    685319.18674803, 685319.18674803, 685319.18674803, 685319.18674803, 
    685319.18674803, 685319.18674803, 685319.18674803, 685319.18674803, 
    685319.18674803, 685319.18674803, 685319.18674803, 685319.18674803,
  722363.467112788, 722363.467112788, 722363.467112788, 722363.467112788, 
    722363.467112788, 722363.467112788, 722363.467112788, 722363.467112788, 
    722363.467112788, 722363.467112788, 722363.467112788, 722363.467112788, 
    722363.467112788, 722363.467112788, 722363.467112788, 722363.467112788, 
    722363.467112788, 722363.467112788, 722363.467112788, 722363.467112788, 
    722363.467112788, 722363.467112788, 722363.467112788, 722363.467112788, 
    722363.467112788, 722363.467112788, 722363.467112788, 722363.467112788, 
    722363.467112788, 722363.467112788, 722363.467112788, 722363.467112788, 
    722363.467112788, 722363.467112788, 722363.467112788, 722363.467112788, 
    722363.467112788, 722363.467112788, 722363.467112788, 722363.467112788, 
    722363.467112788, 722363.467112788, 722363.467112788, 722363.467112788, 
    722363.467112788, 722363.467112788, 722363.467112788, 722363.467112788, 
    722363.467112788, 722363.467112788, 722363.467112788, 722363.467112788, 
    722363.467112788, 722363.467112788, 722363.467112788, 722363.467112788,
  759407.747477546, 759407.747477546, 759407.747477546, 759407.747477546, 
    759407.747477546, 759407.747477546, 759407.747477546, 759407.747477546, 
    759407.747477546, 759407.747477546, 759407.747477546, 759407.747477546, 
    759407.747477546, 759407.747477546, 759407.747477546, 759407.747477546, 
    759407.747477546, 759407.747477546, 759407.747477546, 759407.747477546, 
    759407.747477546, 759407.747477546, 759407.747477546, 759407.747477546, 
    759407.747477546, 759407.747477546, 759407.747477546, 759407.747477546, 
    759407.747477546, 759407.747477546, 759407.747477546, 759407.747477546, 
    759407.747477546, 759407.747477546, 759407.747477546, 759407.747477546, 
    759407.747477546, 759407.747477546, 759407.747477546, 759407.747477546, 
    759407.747477546, 759407.747477546, 759407.747477546, 759407.747477546, 
    759407.747477546, 759407.747477546, 759407.747477546, 759407.747477546, 
    759407.747477546, 759407.747477546, 759407.747477546, 759407.747477546, 
    759407.747477546, 759407.747477546, 759407.747477546, 759407.747477546,
  796452.027842304, 796452.027842304, 796452.027842304, 796452.027842304, 
    796452.027842304, 796452.027842304, 796452.027842304, 796452.027842304, 
    796452.027842304, 796452.027842304, 796452.027842304, 796452.027842304, 
    796452.027842304, 796452.027842304, 796452.027842304, 796452.027842304, 
    796452.027842304, 796452.027842304, 796452.027842304, 796452.027842304, 
    796452.027842304, 796452.027842304, 796452.027842304, 796452.027842304, 
    796452.027842304, 796452.027842304, 796452.027842304, 796452.027842304, 
    796452.027842304, 796452.027842304, 796452.027842304, 796452.027842304, 
    796452.027842304, 796452.027842304, 796452.027842304, 796452.027842304, 
    796452.027842304, 796452.027842304, 796452.027842304, 796452.027842304, 
    796452.027842304, 796452.027842304, 796452.027842304, 796452.027842304, 
    796452.027842304, 796452.027842304, 796452.027842304, 796452.027842304, 
    796452.027842304, 796452.027842304, 796452.027842304, 796452.027842304, 
    796452.027842304, 796452.027842304, 796452.027842304, 796452.027842304,
  833496.308207063, 833496.308207063, 833496.308207063, 833496.308207063, 
    833496.308207063, 833496.308207063, 833496.308207063, 833496.308207063, 
    833496.308207063, 833496.308207063, 833496.308207063, 833496.308207063, 
    833496.308207063, 833496.308207063, 833496.308207063, 833496.308207063, 
    833496.308207063, 833496.308207063, 833496.308207063, 833496.308207063, 
    833496.308207063, 833496.308207063, 833496.308207063, 833496.308207063, 
    833496.308207063, 833496.308207063, 833496.308207063, 833496.308207063, 
    833496.308207063, 833496.308207063, 833496.308207063, 833496.308207063, 
    833496.308207063, 833496.308207063, 833496.308207063, 833496.308207063, 
    833496.308207063, 833496.308207063, 833496.308207063, 833496.308207063, 
    833496.308207063, 833496.308207063, 833496.308207063, 833496.308207063, 
    833496.308207063, 833496.308207063, 833496.308207063, 833496.308207063, 
    833496.308207063, 833496.308207063, 833496.308207063, 833496.308207063, 
    833496.308207063, 833496.308207063, 833496.308207063, 833496.308207063,
  870540.588571821, 870540.588571821, 870540.588571821, 870540.588571821, 
    870540.588571821, 870540.588571821, 870540.588571821, 870540.588571821, 
    870540.588571821, 870540.588571821, 870540.588571821, 870540.588571821, 
    870540.588571821, 870540.588571821, 870540.588571821, 870540.588571821, 
    870540.588571821, 870540.588571821, 870540.588571821, 870540.588571821, 
    870540.588571821, 870540.588571821, 870540.588571821, 870540.588571821, 
    870540.588571821, 870540.588571821, 870540.588571821, 870540.588571821, 
    870540.588571821, 870540.588571821, 870540.588571821, 870540.588571821, 
    870540.588571821, 870540.588571821, 870540.588571821, 870540.588571821, 
    870540.588571821, 870540.588571821, 870540.588571821, 870540.588571821, 
    870540.588571821, 870540.588571821, 870540.588571821, 870540.588571821, 
    870540.588571821, 870540.588571821, 870540.588571821, 870540.588571821, 
    870540.588571821, 870540.588571821, 870540.588571821, 870540.588571821, 
    870540.588571821, 870540.588571821, 870540.588571821, 870540.588571821,
  907584.868936579, 907584.868936579, 907584.868936579, 907584.868936579, 
    907584.868936579, 907584.868936579, 907584.868936579, 907584.868936579, 
    907584.868936579, 907584.868936579, 907584.868936579, 907584.868936579, 
    907584.868936579, 907584.868936579, 907584.868936579, 907584.868936579, 
    907584.868936579, 907584.868936579, 907584.868936579, 907584.868936579, 
    907584.868936579, 907584.868936579, 907584.868936579, 907584.868936579, 
    907584.868936579, 907584.868936579, 907584.868936579, 907584.868936579, 
    907584.868936579, 907584.868936579, 907584.868936579, 907584.868936579, 
    907584.868936579, 907584.868936579, 907584.868936579, 907584.868936579, 
    907584.868936579, 907584.868936579, 907584.868936579, 907584.868936579, 
    907584.868936579, 907584.868936579, 907584.868936579, 907584.868936579, 
    907584.868936579, 907584.868936579, 907584.868936579, 907584.868936579, 
    907584.868936579, 907584.868936579, 907584.868936579, 907584.868936579, 
    907584.868936579, 907584.868936579, 907584.868936579, 907584.868936579,
  944629.149301337, 944629.149301337, 944629.149301337, 944629.149301337, 
    944629.149301337, 944629.149301337, 944629.149301337, 944629.149301337, 
    944629.149301337, 944629.149301337, 944629.149301337, 944629.149301337, 
    944629.149301337, 944629.149301337, 944629.149301337, 944629.149301337, 
    944629.149301337, 944629.149301337, 944629.149301337, 944629.149301337, 
    944629.149301337, 944629.149301337, 944629.149301337, 944629.149301337, 
    944629.149301337, 944629.149301337, 944629.149301337, 944629.149301337, 
    944629.149301337, 944629.149301337, 944629.149301337, 944629.149301337, 
    944629.149301337, 944629.149301337, 944629.149301337, 944629.149301337, 
    944629.149301337, 944629.149301337, 944629.149301337, 944629.149301337, 
    944629.149301337, 944629.149301337, 944629.149301337, 944629.149301337, 
    944629.149301337, 944629.149301337, 944629.149301337, 944629.149301337, 
    944629.149301337, 944629.149301337, 944629.149301337, 944629.149301337, 
    944629.149301337, 944629.149301337, 944629.149301337, 944629.149301337,
  981673.429666096, 981673.429666096, 981673.429666096, 981673.429666096, 
    981673.429666096, 981673.429666096, 981673.429666096, 981673.429666096, 
    981673.429666096, 981673.429666096, 981673.429666096, 981673.429666096, 
    981673.429666096, 981673.429666096, 981673.429666096, 981673.429666096, 
    981673.429666096, 981673.429666096, 981673.429666096, 981673.429666096, 
    981673.429666096, 981673.429666096, 981673.429666096, 981673.429666096, 
    981673.429666096, 981673.429666096, 981673.429666096, 981673.429666096, 
    981673.429666096, 981673.429666096, 981673.429666096, 981673.429666096, 
    981673.429666096, 981673.429666096, 981673.429666096, 981673.429666096, 
    981673.429666096, 981673.429666096, 981673.429666096, 981673.429666096, 
    981673.429666096, 981673.429666096, 981673.429666096, 981673.429666096, 
    981673.429666096, 981673.429666096, 981673.429666096, 981673.429666096, 
    981673.429666096, 981673.429666096, 981673.429666096, 981673.429666096, 
    981673.429666096, 981673.429666096, 981673.429666096, 981673.429666096,
  1018717.71003085, 1018717.71003085, 1018717.71003085, 1018717.71003085, 
    1018717.71003085, 1018717.71003085, 1018717.71003085, 1018717.71003085, 
    1018717.71003085, 1018717.71003085, 1018717.71003085, 1018717.71003085, 
    1018717.71003085, 1018717.71003085, 1018717.71003085, 1018717.71003085, 
    1018717.71003085, 1018717.71003085, 1018717.71003085, 1018717.71003085, 
    1018717.71003085, 1018717.71003085, 1018717.71003085, 1018717.71003085, 
    1018717.71003085, 1018717.71003085, 1018717.71003085, 1018717.71003085, 
    1018717.71003085, 1018717.71003085, 1018717.71003085, 1018717.71003085, 
    1018717.71003085, 1018717.71003085, 1018717.71003085, 1018717.71003085, 
    1018717.71003085, 1018717.71003085, 1018717.71003085, 1018717.71003085, 
    1018717.71003085, 1018717.71003085, 1018717.71003085, 1018717.71003085, 
    1018717.71003085, 1018717.71003085, 1018717.71003085, 1018717.71003085, 
    1018717.71003085, 1018717.71003085, 1018717.71003085, 1018717.71003085, 
    1018717.71003085, 1018717.71003085, 1018717.71003085, 1018717.71003085,
  1055761.99039561, 1055761.99039561, 1055761.99039561, 1055761.99039561, 
    1055761.99039561, 1055761.99039561, 1055761.99039561, 1055761.99039561, 
    1055761.99039561, 1055761.99039561, 1055761.99039561, 1055761.99039561, 
    1055761.99039561, 1055761.99039561, 1055761.99039561, 1055761.99039561, 
    1055761.99039561, 1055761.99039561, 1055761.99039561, 1055761.99039561, 
    1055761.99039561, 1055761.99039561, 1055761.99039561, 1055761.99039561, 
    1055761.99039561, 1055761.99039561, 1055761.99039561, 1055761.99039561, 
    1055761.99039561, 1055761.99039561, 1055761.99039561, 1055761.99039561, 
    1055761.99039561, 1055761.99039561, 1055761.99039561, 1055761.99039561, 
    1055761.99039561, 1055761.99039561, 1055761.99039561, 1055761.99039561, 
    1055761.99039561, 1055761.99039561, 1055761.99039561, 1055761.99039561, 
    1055761.99039561, 1055761.99039561, 1055761.99039561, 1055761.99039561, 
    1055761.99039561, 1055761.99039561, 1055761.99039561, 1055761.99039561, 
    1055761.99039561, 1055761.99039561, 1055761.99039561, 1055761.99039561,
  1092806.27076037, 1092806.27076037, 1092806.27076037, 1092806.27076037, 
    1092806.27076037, 1092806.27076037, 1092806.27076037, 1092806.27076037, 
    1092806.27076037, 1092806.27076037, 1092806.27076037, 1092806.27076037, 
    1092806.27076037, 1092806.27076037, 1092806.27076037, 1092806.27076037, 
    1092806.27076037, 1092806.27076037, 1092806.27076037, 1092806.27076037, 
    1092806.27076037, 1092806.27076037, 1092806.27076037, 1092806.27076037, 
    1092806.27076037, 1092806.27076037, 1092806.27076037, 1092806.27076037, 
    1092806.27076037, 1092806.27076037, 1092806.27076037, 1092806.27076037, 
    1092806.27076037, 1092806.27076037, 1092806.27076037, 1092806.27076037, 
    1092806.27076037, 1092806.27076037, 1092806.27076037, 1092806.27076037, 
    1092806.27076037, 1092806.27076037, 1092806.27076037, 1092806.27076037, 
    1092806.27076037, 1092806.27076037, 1092806.27076037, 1092806.27076037, 
    1092806.27076037, 1092806.27076037, 1092806.27076037, 1092806.27076037, 
    1092806.27076037, 1092806.27076037, 1092806.27076037, 1092806.27076037,
  1129850.55112513, 1129850.55112513, 1129850.55112513, 1129850.55112513, 
    1129850.55112513, 1129850.55112513, 1129850.55112513, 1129850.55112513, 
    1129850.55112513, 1129850.55112513, 1129850.55112513, 1129850.55112513, 
    1129850.55112513, 1129850.55112513, 1129850.55112513, 1129850.55112513, 
    1129850.55112513, 1129850.55112513, 1129850.55112513, 1129850.55112513, 
    1129850.55112513, 1129850.55112513, 1129850.55112513, 1129850.55112513, 
    1129850.55112513, 1129850.55112513, 1129850.55112513, 1129850.55112513, 
    1129850.55112513, 1129850.55112513, 1129850.55112513, 1129850.55112513, 
    1129850.55112513, 1129850.55112513, 1129850.55112513, 1129850.55112513, 
    1129850.55112513, 1129850.55112513, 1129850.55112513, 1129850.55112513, 
    1129850.55112513, 1129850.55112513, 1129850.55112513, 1129850.55112513, 
    1129850.55112513, 1129850.55112513, 1129850.55112513, 1129850.55112513, 
    1129850.55112513, 1129850.55112513, 1129850.55112513, 1129850.55112513, 
    1129850.55112513, 1129850.55112513, 1129850.55112513, 1129850.55112513,
  1166894.83148989, 1166894.83148989, 1166894.83148989, 1166894.83148989, 
    1166894.83148989, 1166894.83148989, 1166894.83148989, 1166894.83148989, 
    1166894.83148989, 1166894.83148989, 1166894.83148989, 1166894.83148989, 
    1166894.83148989, 1166894.83148989, 1166894.83148989, 1166894.83148989, 
    1166894.83148989, 1166894.83148989, 1166894.83148989, 1166894.83148989, 
    1166894.83148989, 1166894.83148989, 1166894.83148989, 1166894.83148989, 
    1166894.83148989, 1166894.83148989, 1166894.83148989, 1166894.83148989, 
    1166894.83148989, 1166894.83148989, 1166894.83148989, 1166894.83148989, 
    1166894.83148989, 1166894.83148989, 1166894.83148989, 1166894.83148989, 
    1166894.83148989, 1166894.83148989, 1166894.83148989, 1166894.83148989, 
    1166894.83148989, 1166894.83148989, 1166894.83148989, 1166894.83148989, 
    1166894.83148989, 1166894.83148989, 1166894.83148989, 1166894.83148989, 
    1166894.83148989, 1166894.83148989, 1166894.83148989, 1166894.83148989, 
    1166894.83148989, 1166894.83148989, 1166894.83148989, 1166894.83148989,
  1203939.11185465, 1203939.11185465, 1203939.11185465, 1203939.11185465, 
    1203939.11185465, 1203939.11185465, 1203939.11185465, 1203939.11185465, 
    1203939.11185465, 1203939.11185465, 1203939.11185465, 1203939.11185465, 
    1203939.11185465, 1203939.11185465, 1203939.11185465, 1203939.11185465, 
    1203939.11185465, 1203939.11185465, 1203939.11185465, 1203939.11185465, 
    1203939.11185465, 1203939.11185465, 1203939.11185465, 1203939.11185465, 
    1203939.11185465, 1203939.11185465, 1203939.11185465, 1203939.11185465, 
    1203939.11185465, 1203939.11185465, 1203939.11185465, 1203939.11185465, 
    1203939.11185465, 1203939.11185465, 1203939.11185465, 1203939.11185465, 
    1203939.11185465, 1203939.11185465, 1203939.11185465, 1203939.11185465, 
    1203939.11185465, 1203939.11185465, 1203939.11185465, 1203939.11185465, 
    1203939.11185465, 1203939.11185465, 1203939.11185465, 1203939.11185465, 
    1203939.11185465, 1203939.11185465, 1203939.11185465, 1203939.11185465, 
    1203939.11185465, 1203939.11185465, 1203939.11185465, 1203939.11185465,
  1240983.3922194, 1240983.3922194, 1240983.3922194, 1240983.3922194, 
    1240983.3922194, 1240983.3922194, 1240983.3922194, 1240983.3922194, 
    1240983.3922194, 1240983.3922194, 1240983.3922194, 1240983.3922194, 
    1240983.3922194, 1240983.3922194, 1240983.3922194, 1240983.3922194, 
    1240983.3922194, 1240983.3922194, 1240983.3922194, 1240983.3922194, 
    1240983.3922194, 1240983.3922194, 1240983.3922194, 1240983.3922194, 
    1240983.3922194, 1240983.3922194, 1240983.3922194, 1240983.3922194, 
    1240983.3922194, 1240983.3922194, 1240983.3922194, 1240983.3922194, 
    1240983.3922194, 1240983.3922194, 1240983.3922194, 1240983.3922194, 
    1240983.3922194, 1240983.3922194, 1240983.3922194, 1240983.3922194, 
    1240983.3922194, 1240983.3922194, 1240983.3922194, 1240983.3922194, 
    1240983.3922194, 1240983.3922194, 1240983.3922194, 1240983.3922194, 
    1240983.3922194, 1240983.3922194, 1240983.3922194, 1240983.3922194, 
    1240983.3922194, 1240983.3922194, 1240983.3922194, 1240983.3922194,
  1278027.67258416, 1278027.67258416, 1278027.67258416, 1278027.67258416, 
    1278027.67258416, 1278027.67258416, 1278027.67258416, 1278027.67258416, 
    1278027.67258416, 1278027.67258416, 1278027.67258416, 1278027.67258416, 
    1278027.67258416, 1278027.67258416, 1278027.67258416, 1278027.67258416, 
    1278027.67258416, 1278027.67258416, 1278027.67258416, 1278027.67258416, 
    1278027.67258416, 1278027.67258416, 1278027.67258416, 1278027.67258416, 
    1278027.67258416, 1278027.67258416, 1278027.67258416, 1278027.67258416, 
    1278027.67258416, 1278027.67258416, 1278027.67258416, 1278027.67258416, 
    1278027.67258416, 1278027.67258416, 1278027.67258416, 1278027.67258416, 
    1278027.67258416, 1278027.67258416, 1278027.67258416, 1278027.67258416, 
    1278027.67258416, 1278027.67258416, 1278027.67258416, 1278027.67258416, 
    1278027.67258416, 1278027.67258416, 1278027.67258416, 1278027.67258416, 
    1278027.67258416, 1278027.67258416, 1278027.67258416, 1278027.67258416, 
    1278027.67258416, 1278027.67258416, 1278027.67258416, 1278027.67258416,
  1315071.95294892, 1315071.95294892, 1315071.95294892, 1315071.95294892, 
    1315071.95294892, 1315071.95294892, 1315071.95294892, 1315071.95294892, 
    1315071.95294892, 1315071.95294892, 1315071.95294892, 1315071.95294892, 
    1315071.95294892, 1315071.95294892, 1315071.95294892, 1315071.95294892, 
    1315071.95294892, 1315071.95294892, 1315071.95294892, 1315071.95294892, 
    1315071.95294892, 1315071.95294892, 1315071.95294892, 1315071.95294892, 
    1315071.95294892, 1315071.95294892, 1315071.95294892, 1315071.95294892, 
    1315071.95294892, 1315071.95294892, 1315071.95294892, 1315071.95294892, 
    1315071.95294892, 1315071.95294892, 1315071.95294892, 1315071.95294892, 
    1315071.95294892, 1315071.95294892, 1315071.95294892, 1315071.95294892, 
    1315071.95294892, 1315071.95294892, 1315071.95294892, 1315071.95294892, 
    1315071.95294892, 1315071.95294892, 1315071.95294892, 1315071.95294892, 
    1315071.95294892, 1315071.95294892, 1315071.95294892, 1315071.95294892, 
    1315071.95294892, 1315071.95294892, 1315071.95294892, 1315071.95294892,
  1352116.23331368, 1352116.23331368, 1352116.23331368, 1352116.23331368, 
    1352116.23331368, 1352116.23331368, 1352116.23331368, 1352116.23331368, 
    1352116.23331368, 1352116.23331368, 1352116.23331368, 1352116.23331368, 
    1352116.23331368, 1352116.23331368, 1352116.23331368, 1352116.23331368, 
    1352116.23331368, 1352116.23331368, 1352116.23331368, 1352116.23331368, 
    1352116.23331368, 1352116.23331368, 1352116.23331368, 1352116.23331368, 
    1352116.23331368, 1352116.23331368, 1352116.23331368, 1352116.23331368, 
    1352116.23331368, 1352116.23331368, 1352116.23331368, 1352116.23331368, 
    1352116.23331368, 1352116.23331368, 1352116.23331368, 1352116.23331368, 
    1352116.23331368, 1352116.23331368, 1352116.23331368, 1352116.23331368, 
    1352116.23331368, 1352116.23331368, 1352116.23331368, 1352116.23331368, 
    1352116.23331368, 1352116.23331368, 1352116.23331368, 1352116.23331368, 
    1352116.23331368, 1352116.23331368, 1352116.23331368, 1352116.23331368, 
    1352116.23331368, 1352116.23331368, 1352116.23331368, 1352116.23331368,
  1389160.51367844, 1389160.51367844, 1389160.51367844, 1389160.51367844, 
    1389160.51367844, 1389160.51367844, 1389160.51367844, 1389160.51367844, 
    1389160.51367844, 1389160.51367844, 1389160.51367844, 1389160.51367844, 
    1389160.51367844, 1389160.51367844, 1389160.51367844, 1389160.51367844, 
    1389160.51367844, 1389160.51367844, 1389160.51367844, 1389160.51367844, 
    1389160.51367844, 1389160.51367844, 1389160.51367844, 1389160.51367844, 
    1389160.51367844, 1389160.51367844, 1389160.51367844, 1389160.51367844, 
    1389160.51367844, 1389160.51367844, 1389160.51367844, 1389160.51367844, 
    1389160.51367844, 1389160.51367844, 1389160.51367844, 1389160.51367844, 
    1389160.51367844, 1389160.51367844, 1389160.51367844, 1389160.51367844, 
    1389160.51367844, 1389160.51367844, 1389160.51367844, 1389160.51367844, 
    1389160.51367844, 1389160.51367844, 1389160.51367844, 1389160.51367844, 
    1389160.51367844, 1389160.51367844, 1389160.51367844, 1389160.51367844, 
    1389160.51367844, 1389160.51367844, 1389160.51367844, 1389160.51367844,
  1426204.7940432, 1426204.7940432, 1426204.7940432, 1426204.7940432, 
    1426204.7940432, 1426204.7940432, 1426204.7940432, 1426204.7940432, 
    1426204.7940432, 1426204.7940432, 1426204.7940432, 1426204.7940432, 
    1426204.7940432, 1426204.7940432, 1426204.7940432, 1426204.7940432, 
    1426204.7940432, 1426204.7940432, 1426204.7940432, 1426204.7940432, 
    1426204.7940432, 1426204.7940432, 1426204.7940432, 1426204.7940432, 
    1426204.7940432, 1426204.7940432, 1426204.7940432, 1426204.7940432, 
    1426204.7940432, 1426204.7940432, 1426204.7940432, 1426204.7940432, 
    1426204.7940432, 1426204.7940432, 1426204.7940432, 1426204.7940432, 
    1426204.7940432, 1426204.7940432, 1426204.7940432, 1426204.7940432, 
    1426204.7940432, 1426204.7940432, 1426204.7940432, 1426204.7940432, 
    1426204.7940432, 1426204.7940432, 1426204.7940432, 1426204.7940432, 
    1426204.7940432, 1426204.7940432, 1426204.7940432, 1426204.7940432, 
    1426204.7940432, 1426204.7940432, 1426204.7940432, 1426204.7940432,
  1463249.07440796, 1463249.07440796, 1463249.07440796, 1463249.07440796, 
    1463249.07440796, 1463249.07440796, 1463249.07440796, 1463249.07440796, 
    1463249.07440796, 1463249.07440796, 1463249.07440796, 1463249.07440796, 
    1463249.07440796, 1463249.07440796, 1463249.07440796, 1463249.07440796, 
    1463249.07440796, 1463249.07440796, 1463249.07440796, 1463249.07440796, 
    1463249.07440796, 1463249.07440796, 1463249.07440796, 1463249.07440796, 
    1463249.07440796, 1463249.07440796, 1463249.07440796, 1463249.07440796, 
    1463249.07440796, 1463249.07440796, 1463249.07440796, 1463249.07440796, 
    1463249.07440796, 1463249.07440796, 1463249.07440796, 1463249.07440796, 
    1463249.07440796, 1463249.07440796, 1463249.07440796, 1463249.07440796, 
    1463249.07440796, 1463249.07440796, 1463249.07440796, 1463249.07440796, 
    1463249.07440796, 1463249.07440796, 1463249.07440796, 1463249.07440796, 
    1463249.07440796, 1463249.07440796, 1463249.07440796, 1463249.07440796, 
    1463249.07440796, 1463249.07440796, 1463249.07440796, 1463249.07440796,
  1500293.35477271, 1500293.35477271, 1500293.35477271, 1500293.35477271, 
    1500293.35477271, 1500293.35477271, 1500293.35477271, 1500293.35477271, 
    1500293.35477271, 1500293.35477271, 1500293.35477271, 1500293.35477271, 
    1500293.35477271, 1500293.35477271, 1500293.35477271, 1500293.35477271, 
    1500293.35477271, 1500293.35477271, 1500293.35477271, 1500293.35477271, 
    1500293.35477271, 1500293.35477271, 1500293.35477271, 1500293.35477271, 
    1500293.35477271, 1500293.35477271, 1500293.35477271, 1500293.35477271, 
    1500293.35477271, 1500293.35477271, 1500293.35477271, 1500293.35477271, 
    1500293.35477271, 1500293.35477271, 1500293.35477271, 1500293.35477271, 
    1500293.35477271, 1500293.35477271, 1500293.35477271, 1500293.35477271, 
    1500293.35477271, 1500293.35477271, 1500293.35477271, 1500293.35477271, 
    1500293.35477271, 1500293.35477271, 1500293.35477271, 1500293.35477271, 
    1500293.35477271, 1500293.35477271, 1500293.35477271, 1500293.35477271, 
    1500293.35477271, 1500293.35477271, 1500293.35477271, 1500293.35477271,
  1537337.63513747, 1537337.63513747, 1537337.63513747, 1537337.63513747, 
    1537337.63513747, 1537337.63513747, 1537337.63513747, 1537337.63513747, 
    1537337.63513747, 1537337.63513747, 1537337.63513747, 1537337.63513747, 
    1537337.63513747, 1537337.63513747, 1537337.63513747, 1537337.63513747, 
    1537337.63513747, 1537337.63513747, 1537337.63513747, 1537337.63513747, 
    1537337.63513747, 1537337.63513747, 1537337.63513747, 1537337.63513747, 
    1537337.63513747, 1537337.63513747, 1537337.63513747, 1537337.63513747, 
    1537337.63513747, 1537337.63513747, 1537337.63513747, 1537337.63513747, 
    1537337.63513747, 1537337.63513747, 1537337.63513747, 1537337.63513747, 
    1537337.63513747, 1537337.63513747, 1537337.63513747, 1537337.63513747, 
    1537337.63513747, 1537337.63513747, 1537337.63513747, 1537337.63513747, 
    1537337.63513747, 1537337.63513747, 1537337.63513747, 1537337.63513747, 
    1537337.63513747, 1537337.63513747, 1537337.63513747, 1537337.63513747, 
    1537337.63513747, 1537337.63513747, 1537337.63513747, 1537337.63513747,
  1574381.91550223, 1574381.91550223, 1574381.91550223, 1574381.91550223, 
    1574381.91550223, 1574381.91550223, 1574381.91550223, 1574381.91550223, 
    1574381.91550223, 1574381.91550223, 1574381.91550223, 1574381.91550223, 
    1574381.91550223, 1574381.91550223, 1574381.91550223, 1574381.91550223, 
    1574381.91550223, 1574381.91550223, 1574381.91550223, 1574381.91550223, 
    1574381.91550223, 1574381.91550223, 1574381.91550223, 1574381.91550223, 
    1574381.91550223, 1574381.91550223, 1574381.91550223, 1574381.91550223, 
    1574381.91550223, 1574381.91550223, 1574381.91550223, 1574381.91550223, 
    1574381.91550223, 1574381.91550223, 1574381.91550223, 1574381.91550223, 
    1574381.91550223, 1574381.91550223, 1574381.91550223, 1574381.91550223, 
    1574381.91550223, 1574381.91550223, 1574381.91550223, 1574381.91550223, 
    1574381.91550223, 1574381.91550223, 1574381.91550223, 1574381.91550223, 
    1574381.91550223, 1574381.91550223, 1574381.91550223, 1574381.91550223, 
    1574381.91550223, 1574381.91550223, 1574381.91550223, 1574381.91550223,
  1611426.19586699, 1611426.19586699, 1611426.19586699, 1611426.19586699, 
    1611426.19586699, 1611426.19586699, 1611426.19586699, 1611426.19586699, 
    1611426.19586699, 1611426.19586699, 1611426.19586699, 1611426.19586699, 
    1611426.19586699, 1611426.19586699, 1611426.19586699, 1611426.19586699, 
    1611426.19586699, 1611426.19586699, 1611426.19586699, 1611426.19586699, 
    1611426.19586699, 1611426.19586699, 1611426.19586699, 1611426.19586699, 
    1611426.19586699, 1611426.19586699, 1611426.19586699, 1611426.19586699, 
    1611426.19586699, 1611426.19586699, 1611426.19586699, 1611426.19586699, 
    1611426.19586699, 1611426.19586699, 1611426.19586699, 1611426.19586699, 
    1611426.19586699, 1611426.19586699, 1611426.19586699, 1611426.19586699, 
    1611426.19586699, 1611426.19586699, 1611426.19586699, 1611426.19586699, 
    1611426.19586699, 1611426.19586699, 1611426.19586699, 1611426.19586699, 
    1611426.19586699, 1611426.19586699, 1611426.19586699, 1611426.19586699, 
    1611426.19586699, 1611426.19586699, 1611426.19586699, 1611426.19586699,
  1648470.47623175, 1648470.47623175, 1648470.47623175, 1648470.47623175, 
    1648470.47623175, 1648470.47623175, 1648470.47623175, 1648470.47623175, 
    1648470.47623175, 1648470.47623175, 1648470.47623175, 1648470.47623175, 
    1648470.47623175, 1648470.47623175, 1648470.47623175, 1648470.47623175, 
    1648470.47623175, 1648470.47623175, 1648470.47623175, 1648470.47623175, 
    1648470.47623175, 1648470.47623175, 1648470.47623175, 1648470.47623175, 
    1648470.47623175, 1648470.47623175, 1648470.47623175, 1648470.47623175, 
    1648470.47623175, 1648470.47623175, 1648470.47623175, 1648470.47623175, 
    1648470.47623175, 1648470.47623175, 1648470.47623175, 1648470.47623175, 
    1648470.47623175, 1648470.47623175, 1648470.47623175, 1648470.47623175, 
    1648470.47623175, 1648470.47623175, 1648470.47623175, 1648470.47623175, 
    1648470.47623175, 1648470.47623175, 1648470.47623175, 1648470.47623175, 
    1648470.47623175, 1648470.47623175, 1648470.47623175, 1648470.47623175, 
    1648470.47623175, 1648470.47623175, 1648470.47623175, 1648470.47623175,
  1685514.75659651, 1685514.75659651, 1685514.75659651, 1685514.75659651, 
    1685514.75659651, 1685514.75659651, 1685514.75659651, 1685514.75659651, 
    1685514.75659651, 1685514.75659651, 1685514.75659651, 1685514.75659651, 
    1685514.75659651, 1685514.75659651, 1685514.75659651, 1685514.75659651, 
    1685514.75659651, 1685514.75659651, 1685514.75659651, 1685514.75659651, 
    1685514.75659651, 1685514.75659651, 1685514.75659651, 1685514.75659651, 
    1685514.75659651, 1685514.75659651, 1685514.75659651, 1685514.75659651, 
    1685514.75659651, 1685514.75659651, 1685514.75659651, 1685514.75659651, 
    1685514.75659651, 1685514.75659651, 1685514.75659651, 1685514.75659651, 
    1685514.75659651, 1685514.75659651, 1685514.75659651, 1685514.75659651, 
    1685514.75659651, 1685514.75659651, 1685514.75659651, 1685514.75659651, 
    1685514.75659651, 1685514.75659651, 1685514.75659651, 1685514.75659651, 
    1685514.75659651, 1685514.75659651, 1685514.75659651, 1685514.75659651, 
    1685514.75659651, 1685514.75659651, 1685514.75659651, 1685514.75659651,
  1722559.03696126, 1722559.03696126, 1722559.03696126, 1722559.03696126, 
    1722559.03696126, 1722559.03696126, 1722559.03696126, 1722559.03696126, 
    1722559.03696126, 1722559.03696126, 1722559.03696126, 1722559.03696126, 
    1722559.03696126, 1722559.03696126, 1722559.03696126, 1722559.03696126, 
    1722559.03696126, 1722559.03696126, 1722559.03696126, 1722559.03696126, 
    1722559.03696126, 1722559.03696126, 1722559.03696126, 1722559.03696126, 
    1722559.03696126, 1722559.03696126, 1722559.03696126, 1722559.03696126, 
    1722559.03696126, 1722559.03696126, 1722559.03696126, 1722559.03696126, 
    1722559.03696126, 1722559.03696126, 1722559.03696126, 1722559.03696126, 
    1722559.03696126, 1722559.03696126, 1722559.03696126, 1722559.03696126, 
    1722559.03696126, 1722559.03696126, 1722559.03696126, 1722559.03696126, 
    1722559.03696126, 1722559.03696126, 1722559.03696126, 1722559.03696126, 
    1722559.03696126, 1722559.03696126, 1722559.03696126, 1722559.03696126, 
    1722559.03696126, 1722559.03696126, 1722559.03696126, 1722559.03696126,
  1759603.31732602, 1759603.31732602, 1759603.31732602, 1759603.31732602, 
    1759603.31732602, 1759603.31732602, 1759603.31732602, 1759603.31732602, 
    1759603.31732602, 1759603.31732602, 1759603.31732602, 1759603.31732602, 
    1759603.31732602, 1759603.31732602, 1759603.31732602, 1759603.31732602, 
    1759603.31732602, 1759603.31732602, 1759603.31732602, 1759603.31732602, 
    1759603.31732602, 1759603.31732602, 1759603.31732602, 1759603.31732602, 
    1759603.31732602, 1759603.31732602, 1759603.31732602, 1759603.31732602, 
    1759603.31732602, 1759603.31732602, 1759603.31732602, 1759603.31732602, 
    1759603.31732602, 1759603.31732602, 1759603.31732602, 1759603.31732602, 
    1759603.31732602, 1759603.31732602, 1759603.31732602, 1759603.31732602, 
    1759603.31732602, 1759603.31732602, 1759603.31732602, 1759603.31732602, 
    1759603.31732602, 1759603.31732602, 1759603.31732602, 1759603.31732602, 
    1759603.31732602, 1759603.31732602, 1759603.31732602, 1759603.31732602, 
    1759603.31732602, 1759603.31732602, 1759603.31732602, 1759603.31732602,
  1796647.59769078, 1796647.59769078, 1796647.59769078, 1796647.59769078, 
    1796647.59769078, 1796647.59769078, 1796647.59769078, 1796647.59769078, 
    1796647.59769078, 1796647.59769078, 1796647.59769078, 1796647.59769078, 
    1796647.59769078, 1796647.59769078, 1796647.59769078, 1796647.59769078, 
    1796647.59769078, 1796647.59769078, 1796647.59769078, 1796647.59769078, 
    1796647.59769078, 1796647.59769078, 1796647.59769078, 1796647.59769078, 
    1796647.59769078, 1796647.59769078, 1796647.59769078, 1796647.59769078, 
    1796647.59769078, 1796647.59769078, 1796647.59769078, 1796647.59769078, 
    1796647.59769078, 1796647.59769078, 1796647.59769078, 1796647.59769078, 
    1796647.59769078, 1796647.59769078, 1796647.59769078, 1796647.59769078, 
    1796647.59769078, 1796647.59769078, 1796647.59769078, 1796647.59769078, 
    1796647.59769078, 1796647.59769078, 1796647.59769078, 1796647.59769078, 
    1796647.59769078, 1796647.59769078, 1796647.59769078, 1796647.59769078, 
    1796647.59769078, 1796647.59769078, 1796647.59769078, 1796647.59769078,
  1833691.87805554, 1833691.87805554, 1833691.87805554, 1833691.87805554, 
    1833691.87805554, 1833691.87805554, 1833691.87805554, 1833691.87805554, 
    1833691.87805554, 1833691.87805554, 1833691.87805554, 1833691.87805554, 
    1833691.87805554, 1833691.87805554, 1833691.87805554, 1833691.87805554, 
    1833691.87805554, 1833691.87805554, 1833691.87805554, 1833691.87805554, 
    1833691.87805554, 1833691.87805554, 1833691.87805554, 1833691.87805554, 
    1833691.87805554, 1833691.87805554, 1833691.87805554, 1833691.87805554, 
    1833691.87805554, 1833691.87805554, 1833691.87805554, 1833691.87805554, 
    1833691.87805554, 1833691.87805554, 1833691.87805554, 1833691.87805554, 
    1833691.87805554, 1833691.87805554, 1833691.87805554, 1833691.87805554, 
    1833691.87805554, 1833691.87805554, 1833691.87805554, 1833691.87805554, 
    1833691.87805554, 1833691.87805554, 1833691.87805554, 1833691.87805554, 
    1833691.87805554, 1833691.87805554, 1833691.87805554, 1833691.87805554, 
    1833691.87805554, 1833691.87805554, 1833691.87805554, 1833691.87805554,
  1870736.1584203, 1870736.1584203, 1870736.1584203, 1870736.1584203, 
    1870736.1584203, 1870736.1584203, 1870736.1584203, 1870736.1584203, 
    1870736.1584203, 1870736.1584203, 1870736.1584203, 1870736.1584203, 
    1870736.1584203, 1870736.1584203, 1870736.1584203, 1870736.1584203, 
    1870736.1584203, 1870736.1584203, 1870736.1584203, 1870736.1584203, 
    1870736.1584203, 1870736.1584203, 1870736.1584203, 1870736.1584203, 
    1870736.1584203, 1870736.1584203, 1870736.1584203, 1870736.1584203, 
    1870736.1584203, 1870736.1584203, 1870736.1584203, 1870736.1584203, 
    1870736.1584203, 1870736.1584203, 1870736.1584203, 1870736.1584203, 
    1870736.1584203, 1870736.1584203, 1870736.1584203, 1870736.1584203, 
    1870736.1584203, 1870736.1584203, 1870736.1584203, 1870736.1584203, 
    1870736.1584203, 1870736.1584203, 1870736.1584203, 1870736.1584203, 
    1870736.1584203, 1870736.1584203, 1870736.1584203, 1870736.1584203, 
    1870736.1584203, 1870736.1584203, 1870736.1584203, 1870736.1584203,
  1907780.43878506, 1907780.43878506, 1907780.43878506, 1907780.43878506, 
    1907780.43878506, 1907780.43878506, 1907780.43878506, 1907780.43878506, 
    1907780.43878506, 1907780.43878506, 1907780.43878506, 1907780.43878506, 
    1907780.43878506, 1907780.43878506, 1907780.43878506, 1907780.43878506, 
    1907780.43878506, 1907780.43878506, 1907780.43878506, 1907780.43878506, 
    1907780.43878506, 1907780.43878506, 1907780.43878506, 1907780.43878506, 
    1907780.43878506, 1907780.43878506, 1907780.43878506, 1907780.43878506, 
    1907780.43878506, 1907780.43878506, 1907780.43878506, 1907780.43878506, 
    1907780.43878506, 1907780.43878506, 1907780.43878506, 1907780.43878506, 
    1907780.43878506, 1907780.43878506, 1907780.43878506, 1907780.43878506, 
    1907780.43878506, 1907780.43878506, 1907780.43878506, 1907780.43878506, 
    1907780.43878506, 1907780.43878506, 1907780.43878506, 1907780.43878506, 
    1907780.43878506, 1907780.43878506, 1907780.43878506, 1907780.43878506, 
    1907780.43878506, 1907780.43878506, 1907780.43878506, 1907780.43878506,
  1944824.71914981, 1944824.71914981, 1944824.71914981, 1944824.71914981, 
    1944824.71914981, 1944824.71914981, 1944824.71914981, 1944824.71914981, 
    1944824.71914981, 1944824.71914981, 1944824.71914981, 1944824.71914981, 
    1944824.71914981, 1944824.71914981, 1944824.71914981, 1944824.71914981, 
    1944824.71914981, 1944824.71914981, 1944824.71914981, 1944824.71914981, 
    1944824.71914981, 1944824.71914981, 1944824.71914981, 1944824.71914981, 
    1944824.71914981, 1944824.71914981, 1944824.71914981, 1944824.71914981, 
    1944824.71914981, 1944824.71914981, 1944824.71914981, 1944824.71914981, 
    1944824.71914981, 1944824.71914981, 1944824.71914981, 1944824.71914981, 
    1944824.71914981, 1944824.71914981, 1944824.71914981, 1944824.71914981, 
    1944824.71914981, 1944824.71914981, 1944824.71914981, 1944824.71914981, 
    1944824.71914981, 1944824.71914981, 1944824.71914981, 1944824.71914981, 
    1944824.71914981, 1944824.71914981, 1944824.71914981, 1944824.71914981, 
    1944824.71914981, 1944824.71914981, 1944824.71914981, 1944824.71914981,
  1981868.99951457, 1981868.99951457, 1981868.99951457, 1981868.99951457, 
    1981868.99951457, 1981868.99951457, 1981868.99951457, 1981868.99951457, 
    1981868.99951457, 1981868.99951457, 1981868.99951457, 1981868.99951457, 
    1981868.99951457, 1981868.99951457, 1981868.99951457, 1981868.99951457, 
    1981868.99951457, 1981868.99951457, 1981868.99951457, 1981868.99951457, 
    1981868.99951457, 1981868.99951457, 1981868.99951457, 1981868.99951457, 
    1981868.99951457, 1981868.99951457, 1981868.99951457, 1981868.99951457, 
    1981868.99951457, 1981868.99951457, 1981868.99951457, 1981868.99951457, 
    1981868.99951457, 1981868.99951457, 1981868.99951457, 1981868.99951457, 
    1981868.99951457, 1981868.99951457, 1981868.99951457, 1981868.99951457, 
    1981868.99951457, 1981868.99951457, 1981868.99951457, 1981868.99951457, 
    1981868.99951457, 1981868.99951457, 1981868.99951457, 1981868.99951457, 
    1981868.99951457, 1981868.99951457, 1981868.99951457, 1981868.99951457, 
    1981868.99951457, 1981868.99951457, 1981868.99951457, 1981868.99951457 ;

 y_psi =
  18522.1401823791, 18522.1401823791, 18522.1401823791, 18522.1401823791, 
    18522.1401823791, 18522.1401823791, 18522.1401823791, 18522.1401823791, 
    18522.1401823791, 18522.1401823791, 18522.1401823791, 18522.1401823791, 
    18522.1401823791, 18522.1401823791, 18522.1401823791, 18522.1401823791, 
    18522.1401823791, 18522.1401823791, 18522.1401823791, 18522.1401823791, 
    18522.1401823791, 18522.1401823791, 18522.1401823791, 18522.1401823791, 
    18522.1401823791, 18522.1401823791, 18522.1401823791, 18522.1401823791, 
    18522.1401823791, 18522.1401823791, 18522.1401823791, 18522.1401823791, 
    18522.1401823791, 18522.1401823791, 18522.1401823791, 18522.1401823791, 
    18522.1401823791, 18522.1401823791, 18522.1401823791, 18522.1401823791, 
    18522.1401823791, 18522.1401823791, 18522.1401823791, 18522.1401823791, 
    18522.1401823791, 18522.1401823791, 18522.1401823791, 18522.1401823791, 
    18522.1401823791, 18522.1401823791, 18522.1401823791, 18522.1401823791, 
    18522.1401823791, 18522.1401823791, 18522.1401823791,
  55566.4205471374, 55566.4205471374, 55566.4205471374, 55566.4205471374, 
    55566.4205471374, 55566.4205471374, 55566.4205471374, 55566.4205471374, 
    55566.4205471374, 55566.4205471374, 55566.4205471374, 55566.4205471374, 
    55566.4205471374, 55566.4205471374, 55566.4205471374, 55566.4205471374, 
    55566.4205471374, 55566.4205471374, 55566.4205471374, 55566.4205471374, 
    55566.4205471374, 55566.4205471374, 55566.4205471374, 55566.4205471374, 
    55566.4205471374, 55566.4205471374, 55566.4205471374, 55566.4205471374, 
    55566.4205471374, 55566.4205471374, 55566.4205471374, 55566.4205471374, 
    55566.4205471374, 55566.4205471374, 55566.4205471374, 55566.4205471374, 
    55566.4205471374, 55566.4205471374, 55566.4205471374, 55566.4205471374, 
    55566.4205471374, 55566.4205471374, 55566.4205471374, 55566.4205471374, 
    55566.4205471374, 55566.4205471374, 55566.4205471374, 55566.4205471374, 
    55566.4205471374, 55566.4205471374, 55566.4205471374, 55566.4205471374, 
    55566.4205471374, 55566.4205471374, 55566.4205471374,
  92610.7009118959, 92610.7009118959, 92610.7009118959, 92610.7009118959, 
    92610.7009118959, 92610.7009118959, 92610.7009118959, 92610.7009118959, 
    92610.7009118959, 92610.7009118959, 92610.7009118959, 92610.7009118959, 
    92610.7009118959, 92610.7009118959, 92610.7009118959, 92610.7009118959, 
    92610.7009118959, 92610.7009118959, 92610.7009118959, 92610.7009118959, 
    92610.7009118959, 92610.7009118959, 92610.7009118959, 92610.7009118959, 
    92610.7009118959, 92610.7009118959, 92610.7009118959, 92610.7009118959, 
    92610.7009118959, 92610.7009118959, 92610.7009118959, 92610.7009118959, 
    92610.7009118959, 92610.7009118959, 92610.7009118959, 92610.7009118959, 
    92610.7009118959, 92610.7009118959, 92610.7009118959, 92610.7009118959, 
    92610.7009118959, 92610.7009118959, 92610.7009118959, 92610.7009118959, 
    92610.7009118959, 92610.7009118959, 92610.7009118959, 92610.7009118959, 
    92610.7009118959, 92610.7009118959, 92610.7009118959, 92610.7009118959, 
    92610.7009118959, 92610.7009118959, 92610.7009118959,
  129654.981276654, 129654.981276654, 129654.981276654, 129654.981276654, 
    129654.981276654, 129654.981276654, 129654.981276654, 129654.981276654, 
    129654.981276654, 129654.981276654, 129654.981276654, 129654.981276654, 
    129654.981276654, 129654.981276654, 129654.981276654, 129654.981276654, 
    129654.981276654, 129654.981276654, 129654.981276654, 129654.981276654, 
    129654.981276654, 129654.981276654, 129654.981276654, 129654.981276654, 
    129654.981276654, 129654.981276654, 129654.981276654, 129654.981276654, 
    129654.981276654, 129654.981276654, 129654.981276654, 129654.981276654, 
    129654.981276654, 129654.981276654, 129654.981276654, 129654.981276654, 
    129654.981276654, 129654.981276654, 129654.981276654, 129654.981276654, 
    129654.981276654, 129654.981276654, 129654.981276654, 129654.981276654, 
    129654.981276654, 129654.981276654, 129654.981276654, 129654.981276654, 
    129654.981276654, 129654.981276654, 129654.981276654, 129654.981276654, 
    129654.981276654, 129654.981276654, 129654.981276654,
  166699.261641412, 166699.261641412, 166699.261641412, 166699.261641412, 
    166699.261641412, 166699.261641412, 166699.261641412, 166699.261641412, 
    166699.261641412, 166699.261641412, 166699.261641412, 166699.261641412, 
    166699.261641412, 166699.261641412, 166699.261641412, 166699.261641412, 
    166699.261641412, 166699.261641412, 166699.261641412, 166699.261641412, 
    166699.261641412, 166699.261641412, 166699.261641412, 166699.261641412, 
    166699.261641412, 166699.261641412, 166699.261641412, 166699.261641412, 
    166699.261641412, 166699.261641412, 166699.261641412, 166699.261641412, 
    166699.261641412, 166699.261641412, 166699.261641412, 166699.261641412, 
    166699.261641412, 166699.261641412, 166699.261641412, 166699.261641412, 
    166699.261641412, 166699.261641412, 166699.261641412, 166699.261641412, 
    166699.261641412, 166699.261641412, 166699.261641412, 166699.261641412, 
    166699.261641412, 166699.261641412, 166699.261641412, 166699.261641412, 
    166699.261641412, 166699.261641412, 166699.261641412,
  203743.542006171, 203743.542006171, 203743.542006171, 203743.542006171, 
    203743.542006171, 203743.542006171, 203743.542006171, 203743.542006171, 
    203743.542006171, 203743.542006171, 203743.542006171, 203743.542006171, 
    203743.542006171, 203743.542006171, 203743.542006171, 203743.542006171, 
    203743.542006171, 203743.542006171, 203743.542006171, 203743.542006171, 
    203743.542006171, 203743.542006171, 203743.542006171, 203743.542006171, 
    203743.542006171, 203743.542006171, 203743.542006171, 203743.542006171, 
    203743.542006171, 203743.542006171, 203743.542006171, 203743.542006171, 
    203743.542006171, 203743.542006171, 203743.542006171, 203743.542006171, 
    203743.542006171, 203743.542006171, 203743.542006171, 203743.542006171, 
    203743.542006171, 203743.542006171, 203743.542006171, 203743.542006171, 
    203743.542006171, 203743.542006171, 203743.542006171, 203743.542006171, 
    203743.542006171, 203743.542006171, 203743.542006171, 203743.542006171, 
    203743.542006171, 203743.542006171, 203743.542006171,
  240787.82237093, 240787.82237093, 240787.82237093, 240787.82237093, 
    240787.82237093, 240787.82237093, 240787.82237093, 240787.82237093, 
    240787.82237093, 240787.82237093, 240787.82237093, 240787.82237093, 
    240787.82237093, 240787.82237093, 240787.82237093, 240787.82237093, 
    240787.82237093, 240787.82237093, 240787.82237093, 240787.82237093, 
    240787.82237093, 240787.82237093, 240787.82237093, 240787.82237093, 
    240787.82237093, 240787.82237093, 240787.82237093, 240787.82237093, 
    240787.82237093, 240787.82237093, 240787.82237093, 240787.82237093, 
    240787.82237093, 240787.82237093, 240787.82237093, 240787.82237093, 
    240787.82237093, 240787.82237093, 240787.82237093, 240787.82237093, 
    240787.82237093, 240787.82237093, 240787.82237093, 240787.82237093, 
    240787.82237093, 240787.82237093, 240787.82237093, 240787.82237093, 
    240787.82237093, 240787.82237093, 240787.82237093, 240787.82237093, 
    240787.82237093, 240787.82237093, 240787.82237093,
  277832.102735688, 277832.102735688, 277832.102735688, 277832.102735688, 
    277832.102735688, 277832.102735688, 277832.102735688, 277832.102735688, 
    277832.102735688, 277832.102735688, 277832.102735688, 277832.102735688, 
    277832.102735688, 277832.102735688, 277832.102735688, 277832.102735688, 
    277832.102735688, 277832.102735688, 277832.102735688, 277832.102735688, 
    277832.102735688, 277832.102735688, 277832.102735688, 277832.102735688, 
    277832.102735688, 277832.102735688, 277832.102735688, 277832.102735688, 
    277832.102735688, 277832.102735688, 277832.102735688, 277832.102735688, 
    277832.102735688, 277832.102735688, 277832.102735688, 277832.102735688, 
    277832.102735688, 277832.102735688, 277832.102735688, 277832.102735688, 
    277832.102735688, 277832.102735688, 277832.102735688, 277832.102735688, 
    277832.102735688, 277832.102735688, 277832.102735688, 277832.102735688, 
    277832.102735688, 277832.102735688, 277832.102735688, 277832.102735688, 
    277832.102735688, 277832.102735688, 277832.102735688,
  314876.383100447, 314876.383100447, 314876.383100447, 314876.383100447, 
    314876.383100447, 314876.383100447, 314876.383100447, 314876.383100447, 
    314876.383100447, 314876.383100447, 314876.383100447, 314876.383100447, 
    314876.383100447, 314876.383100447, 314876.383100447, 314876.383100447, 
    314876.383100447, 314876.383100447, 314876.383100447, 314876.383100447, 
    314876.383100447, 314876.383100447, 314876.383100447, 314876.383100447, 
    314876.383100447, 314876.383100447, 314876.383100447, 314876.383100447, 
    314876.383100447, 314876.383100447, 314876.383100447, 314876.383100447, 
    314876.383100447, 314876.383100447, 314876.383100447, 314876.383100447, 
    314876.383100447, 314876.383100447, 314876.383100447, 314876.383100447, 
    314876.383100447, 314876.383100447, 314876.383100447, 314876.383100447, 
    314876.383100447, 314876.383100447, 314876.383100447, 314876.383100447, 
    314876.383100447, 314876.383100447, 314876.383100447, 314876.383100447, 
    314876.383100447, 314876.383100447, 314876.383100447,
  351920.663465205, 351920.663465205, 351920.663465205, 351920.663465205, 
    351920.663465205, 351920.663465205, 351920.663465205, 351920.663465205, 
    351920.663465205, 351920.663465205, 351920.663465205, 351920.663465205, 
    351920.663465205, 351920.663465205, 351920.663465205, 351920.663465205, 
    351920.663465205, 351920.663465205, 351920.663465205, 351920.663465205, 
    351920.663465205, 351920.663465205, 351920.663465205, 351920.663465205, 
    351920.663465205, 351920.663465205, 351920.663465205, 351920.663465205, 
    351920.663465205, 351920.663465205, 351920.663465205, 351920.663465205, 
    351920.663465205, 351920.663465205, 351920.663465205, 351920.663465205, 
    351920.663465205, 351920.663465205, 351920.663465205, 351920.663465205, 
    351920.663465205, 351920.663465205, 351920.663465205, 351920.663465205, 
    351920.663465205, 351920.663465205, 351920.663465205, 351920.663465205, 
    351920.663465205, 351920.663465205, 351920.663465205, 351920.663465205, 
    351920.663465205, 351920.663465205, 351920.663465205,
  388964.943829963, 388964.943829963, 388964.943829963, 388964.943829963, 
    388964.943829963, 388964.943829963, 388964.943829963, 388964.943829963, 
    388964.943829963, 388964.943829963, 388964.943829963, 388964.943829963, 
    388964.943829963, 388964.943829963, 388964.943829963, 388964.943829963, 
    388964.943829963, 388964.943829963, 388964.943829963, 388964.943829963, 
    388964.943829963, 388964.943829963, 388964.943829963, 388964.943829963, 
    388964.943829963, 388964.943829963, 388964.943829963, 388964.943829963, 
    388964.943829963, 388964.943829963, 388964.943829963, 388964.943829963, 
    388964.943829963, 388964.943829963, 388964.943829963, 388964.943829963, 
    388964.943829963, 388964.943829963, 388964.943829963, 388964.943829963, 
    388964.943829963, 388964.943829963, 388964.943829963, 388964.943829963, 
    388964.943829963, 388964.943829963, 388964.943829963, 388964.943829963, 
    388964.943829963, 388964.943829963, 388964.943829963, 388964.943829963, 
    388964.943829963, 388964.943829963, 388964.943829963,
  426009.224194721, 426009.224194721, 426009.224194721, 426009.224194721, 
    426009.224194721, 426009.224194721, 426009.224194721, 426009.224194721, 
    426009.224194721, 426009.224194721, 426009.224194721, 426009.224194721, 
    426009.224194721, 426009.224194721, 426009.224194721, 426009.224194721, 
    426009.224194721, 426009.224194721, 426009.224194721, 426009.224194721, 
    426009.224194721, 426009.224194721, 426009.224194721, 426009.224194721, 
    426009.224194721, 426009.224194721, 426009.224194721, 426009.224194721, 
    426009.224194721, 426009.224194721, 426009.224194721, 426009.224194721, 
    426009.224194721, 426009.224194721, 426009.224194721, 426009.224194721, 
    426009.224194721, 426009.224194721, 426009.224194721, 426009.224194721, 
    426009.224194721, 426009.224194721, 426009.224194721, 426009.224194721, 
    426009.224194721, 426009.224194721, 426009.224194721, 426009.224194721, 
    426009.224194721, 426009.224194721, 426009.224194721, 426009.224194721, 
    426009.224194721, 426009.224194721, 426009.224194721,
  463053.50455948, 463053.50455948, 463053.50455948, 463053.50455948, 
    463053.50455948, 463053.50455948, 463053.50455948, 463053.50455948, 
    463053.50455948, 463053.50455948, 463053.50455948, 463053.50455948, 
    463053.50455948, 463053.50455948, 463053.50455948, 463053.50455948, 
    463053.50455948, 463053.50455948, 463053.50455948, 463053.50455948, 
    463053.50455948, 463053.50455948, 463053.50455948, 463053.50455948, 
    463053.50455948, 463053.50455948, 463053.50455948, 463053.50455948, 
    463053.50455948, 463053.50455948, 463053.50455948, 463053.50455948, 
    463053.50455948, 463053.50455948, 463053.50455948, 463053.50455948, 
    463053.50455948, 463053.50455948, 463053.50455948, 463053.50455948, 
    463053.50455948, 463053.50455948, 463053.50455948, 463053.50455948, 
    463053.50455948, 463053.50455948, 463053.50455948, 463053.50455948, 
    463053.50455948, 463053.50455948, 463053.50455948, 463053.50455948, 
    463053.50455948, 463053.50455948, 463053.50455948,
  500097.784924238, 500097.784924238, 500097.784924238, 500097.784924238, 
    500097.784924238, 500097.784924238, 500097.784924238, 500097.784924238, 
    500097.784924238, 500097.784924238, 500097.784924238, 500097.784924238, 
    500097.784924238, 500097.784924238, 500097.784924238, 500097.784924238, 
    500097.784924238, 500097.784924238, 500097.784924238, 500097.784924238, 
    500097.784924238, 500097.784924238, 500097.784924238, 500097.784924238, 
    500097.784924238, 500097.784924238, 500097.784924238, 500097.784924238, 
    500097.784924238, 500097.784924238, 500097.784924238, 500097.784924238, 
    500097.784924238, 500097.784924238, 500097.784924238, 500097.784924238, 
    500097.784924238, 500097.784924238, 500097.784924238, 500097.784924238, 
    500097.784924238, 500097.784924238, 500097.784924238, 500097.784924238, 
    500097.784924238, 500097.784924238, 500097.784924238, 500097.784924238, 
    500097.784924238, 500097.784924238, 500097.784924238, 500097.784924238, 
    500097.784924238, 500097.784924238, 500097.784924238,
  537142.065288996, 537142.065288996, 537142.065288996, 537142.065288996, 
    537142.065288996, 537142.065288996, 537142.065288996, 537142.065288996, 
    537142.065288996, 537142.065288996, 537142.065288996, 537142.065288996, 
    537142.065288996, 537142.065288996, 537142.065288996, 537142.065288996, 
    537142.065288996, 537142.065288996, 537142.065288996, 537142.065288996, 
    537142.065288996, 537142.065288996, 537142.065288996, 537142.065288996, 
    537142.065288996, 537142.065288996, 537142.065288996, 537142.065288996, 
    537142.065288996, 537142.065288996, 537142.065288996, 537142.065288996, 
    537142.065288996, 537142.065288996, 537142.065288996, 537142.065288996, 
    537142.065288996, 537142.065288996, 537142.065288996, 537142.065288996, 
    537142.065288996, 537142.065288996, 537142.065288996, 537142.065288996, 
    537142.065288996, 537142.065288996, 537142.065288996, 537142.065288996, 
    537142.065288996, 537142.065288996, 537142.065288996, 537142.065288996, 
    537142.065288996, 537142.065288996, 537142.065288996,
  574186.345653754, 574186.345653754, 574186.345653754, 574186.345653754, 
    574186.345653754, 574186.345653754, 574186.345653754, 574186.345653754, 
    574186.345653754, 574186.345653754, 574186.345653754, 574186.345653754, 
    574186.345653754, 574186.345653754, 574186.345653754, 574186.345653754, 
    574186.345653754, 574186.345653754, 574186.345653754, 574186.345653754, 
    574186.345653754, 574186.345653754, 574186.345653754, 574186.345653754, 
    574186.345653754, 574186.345653754, 574186.345653754, 574186.345653754, 
    574186.345653754, 574186.345653754, 574186.345653754, 574186.345653754, 
    574186.345653754, 574186.345653754, 574186.345653754, 574186.345653754, 
    574186.345653754, 574186.345653754, 574186.345653754, 574186.345653754, 
    574186.345653754, 574186.345653754, 574186.345653754, 574186.345653754, 
    574186.345653754, 574186.345653754, 574186.345653754, 574186.345653754, 
    574186.345653754, 574186.345653754, 574186.345653754, 574186.345653754, 
    574186.345653754, 574186.345653754, 574186.345653754,
  611230.626018513, 611230.626018513, 611230.626018513, 611230.626018513, 
    611230.626018513, 611230.626018513, 611230.626018513, 611230.626018513, 
    611230.626018513, 611230.626018513, 611230.626018513, 611230.626018513, 
    611230.626018513, 611230.626018513, 611230.626018513, 611230.626018513, 
    611230.626018513, 611230.626018513, 611230.626018513, 611230.626018513, 
    611230.626018513, 611230.626018513, 611230.626018513, 611230.626018513, 
    611230.626018513, 611230.626018513, 611230.626018513, 611230.626018513, 
    611230.626018513, 611230.626018513, 611230.626018513, 611230.626018513, 
    611230.626018513, 611230.626018513, 611230.626018513, 611230.626018513, 
    611230.626018513, 611230.626018513, 611230.626018513, 611230.626018513, 
    611230.626018513, 611230.626018513, 611230.626018513, 611230.626018513, 
    611230.626018513, 611230.626018513, 611230.626018513, 611230.626018513, 
    611230.626018513, 611230.626018513, 611230.626018513, 611230.626018513, 
    611230.626018513, 611230.626018513, 611230.626018513,
  648274.906383271, 648274.906383271, 648274.906383271, 648274.906383271, 
    648274.906383271, 648274.906383271, 648274.906383271, 648274.906383271, 
    648274.906383271, 648274.906383271, 648274.906383271, 648274.906383271, 
    648274.906383271, 648274.906383271, 648274.906383271, 648274.906383271, 
    648274.906383271, 648274.906383271, 648274.906383271, 648274.906383271, 
    648274.906383271, 648274.906383271, 648274.906383271, 648274.906383271, 
    648274.906383271, 648274.906383271, 648274.906383271, 648274.906383271, 
    648274.906383271, 648274.906383271, 648274.906383271, 648274.906383271, 
    648274.906383271, 648274.906383271, 648274.906383271, 648274.906383271, 
    648274.906383271, 648274.906383271, 648274.906383271, 648274.906383271, 
    648274.906383271, 648274.906383271, 648274.906383271, 648274.906383271, 
    648274.906383271, 648274.906383271, 648274.906383271, 648274.906383271, 
    648274.906383271, 648274.906383271, 648274.906383271, 648274.906383271, 
    648274.906383271, 648274.906383271, 648274.906383271,
  685319.18674803, 685319.18674803, 685319.18674803, 685319.18674803, 
    685319.18674803, 685319.18674803, 685319.18674803, 685319.18674803, 
    685319.18674803, 685319.18674803, 685319.18674803, 685319.18674803, 
    685319.18674803, 685319.18674803, 685319.18674803, 685319.18674803, 
    685319.18674803, 685319.18674803, 685319.18674803, 685319.18674803, 
    685319.18674803, 685319.18674803, 685319.18674803, 685319.18674803, 
    685319.18674803, 685319.18674803, 685319.18674803, 685319.18674803, 
    685319.18674803, 685319.18674803, 685319.18674803, 685319.18674803, 
    685319.18674803, 685319.18674803, 685319.18674803, 685319.18674803, 
    685319.18674803, 685319.18674803, 685319.18674803, 685319.18674803, 
    685319.18674803, 685319.18674803, 685319.18674803, 685319.18674803, 
    685319.18674803, 685319.18674803, 685319.18674803, 685319.18674803, 
    685319.18674803, 685319.18674803, 685319.18674803, 685319.18674803, 
    685319.18674803, 685319.18674803, 685319.18674803,
  722363.467112788, 722363.467112788, 722363.467112788, 722363.467112788, 
    722363.467112788, 722363.467112788, 722363.467112788, 722363.467112788, 
    722363.467112788, 722363.467112788, 722363.467112788, 722363.467112788, 
    722363.467112788, 722363.467112788, 722363.467112788, 722363.467112788, 
    722363.467112788, 722363.467112788, 722363.467112788, 722363.467112788, 
    722363.467112788, 722363.467112788, 722363.467112788, 722363.467112788, 
    722363.467112788, 722363.467112788, 722363.467112788, 722363.467112788, 
    722363.467112788, 722363.467112788, 722363.467112788, 722363.467112788, 
    722363.467112788, 722363.467112788, 722363.467112788, 722363.467112788, 
    722363.467112788, 722363.467112788, 722363.467112788, 722363.467112788, 
    722363.467112788, 722363.467112788, 722363.467112788, 722363.467112788, 
    722363.467112788, 722363.467112788, 722363.467112788, 722363.467112788, 
    722363.467112788, 722363.467112788, 722363.467112788, 722363.467112788, 
    722363.467112788, 722363.467112788, 722363.467112788,
  759407.747477546, 759407.747477546, 759407.747477546, 759407.747477546, 
    759407.747477546, 759407.747477546, 759407.747477546, 759407.747477546, 
    759407.747477546, 759407.747477546, 759407.747477546, 759407.747477546, 
    759407.747477546, 759407.747477546, 759407.747477546, 759407.747477546, 
    759407.747477546, 759407.747477546, 759407.747477546, 759407.747477546, 
    759407.747477546, 759407.747477546, 759407.747477546, 759407.747477546, 
    759407.747477546, 759407.747477546, 759407.747477546, 759407.747477546, 
    759407.747477546, 759407.747477546, 759407.747477546, 759407.747477546, 
    759407.747477546, 759407.747477546, 759407.747477546, 759407.747477546, 
    759407.747477546, 759407.747477546, 759407.747477546, 759407.747477546, 
    759407.747477546, 759407.747477546, 759407.747477546, 759407.747477546, 
    759407.747477546, 759407.747477546, 759407.747477546, 759407.747477546, 
    759407.747477546, 759407.747477546, 759407.747477546, 759407.747477546, 
    759407.747477546, 759407.747477546, 759407.747477546,
  796452.027842304, 796452.027842304, 796452.027842304, 796452.027842304, 
    796452.027842304, 796452.027842304, 796452.027842304, 796452.027842304, 
    796452.027842304, 796452.027842304, 796452.027842304, 796452.027842304, 
    796452.027842304, 796452.027842304, 796452.027842304, 796452.027842304, 
    796452.027842304, 796452.027842304, 796452.027842304, 796452.027842304, 
    796452.027842304, 796452.027842304, 796452.027842304, 796452.027842304, 
    796452.027842304, 796452.027842304, 796452.027842304, 796452.027842304, 
    796452.027842304, 796452.027842304, 796452.027842304, 796452.027842304, 
    796452.027842304, 796452.027842304, 796452.027842304, 796452.027842304, 
    796452.027842304, 796452.027842304, 796452.027842304, 796452.027842304, 
    796452.027842304, 796452.027842304, 796452.027842304, 796452.027842304, 
    796452.027842304, 796452.027842304, 796452.027842304, 796452.027842304, 
    796452.027842304, 796452.027842304, 796452.027842304, 796452.027842304, 
    796452.027842304, 796452.027842304, 796452.027842304,
  833496.308207063, 833496.308207063, 833496.308207063, 833496.308207063, 
    833496.308207063, 833496.308207063, 833496.308207063, 833496.308207063, 
    833496.308207063, 833496.308207063, 833496.308207063, 833496.308207063, 
    833496.308207063, 833496.308207063, 833496.308207063, 833496.308207063, 
    833496.308207063, 833496.308207063, 833496.308207063, 833496.308207063, 
    833496.308207063, 833496.308207063, 833496.308207063, 833496.308207063, 
    833496.308207063, 833496.308207063, 833496.308207063, 833496.308207063, 
    833496.308207063, 833496.308207063, 833496.308207063, 833496.308207063, 
    833496.308207063, 833496.308207063, 833496.308207063, 833496.308207063, 
    833496.308207063, 833496.308207063, 833496.308207063, 833496.308207063, 
    833496.308207063, 833496.308207063, 833496.308207063, 833496.308207063, 
    833496.308207063, 833496.308207063, 833496.308207063, 833496.308207063, 
    833496.308207063, 833496.308207063, 833496.308207063, 833496.308207063, 
    833496.308207063, 833496.308207063, 833496.308207063,
  870540.588571821, 870540.588571821, 870540.588571821, 870540.588571821, 
    870540.588571821, 870540.588571821, 870540.588571821, 870540.588571821, 
    870540.588571821, 870540.588571821, 870540.588571821, 870540.588571821, 
    870540.588571821, 870540.588571821, 870540.588571821, 870540.588571821, 
    870540.588571821, 870540.588571821, 870540.588571821, 870540.588571821, 
    870540.588571821, 870540.588571821, 870540.588571821, 870540.588571821, 
    870540.588571821, 870540.588571821, 870540.588571821, 870540.588571821, 
    870540.588571821, 870540.588571821, 870540.588571821, 870540.588571821, 
    870540.588571821, 870540.588571821, 870540.588571821, 870540.588571821, 
    870540.588571821, 870540.588571821, 870540.588571821, 870540.588571821, 
    870540.588571821, 870540.588571821, 870540.588571821, 870540.588571821, 
    870540.588571821, 870540.588571821, 870540.588571821, 870540.588571821, 
    870540.588571821, 870540.588571821, 870540.588571821, 870540.588571821, 
    870540.588571821, 870540.588571821, 870540.588571821,
  907584.868936579, 907584.868936579, 907584.868936579, 907584.868936579, 
    907584.868936579, 907584.868936579, 907584.868936579, 907584.868936579, 
    907584.868936579, 907584.868936579, 907584.868936579, 907584.868936579, 
    907584.868936579, 907584.868936579, 907584.868936579, 907584.868936579, 
    907584.868936579, 907584.868936579, 907584.868936579, 907584.868936579, 
    907584.868936579, 907584.868936579, 907584.868936579, 907584.868936579, 
    907584.868936579, 907584.868936579, 907584.868936579, 907584.868936579, 
    907584.868936579, 907584.868936579, 907584.868936579, 907584.868936579, 
    907584.868936579, 907584.868936579, 907584.868936579, 907584.868936579, 
    907584.868936579, 907584.868936579, 907584.868936579, 907584.868936579, 
    907584.868936579, 907584.868936579, 907584.868936579, 907584.868936579, 
    907584.868936579, 907584.868936579, 907584.868936579, 907584.868936579, 
    907584.868936579, 907584.868936579, 907584.868936579, 907584.868936579, 
    907584.868936579, 907584.868936579, 907584.868936579,
  944629.149301337, 944629.149301337, 944629.149301337, 944629.149301337, 
    944629.149301337, 944629.149301337, 944629.149301337, 944629.149301337, 
    944629.149301337, 944629.149301337, 944629.149301337, 944629.149301337, 
    944629.149301337, 944629.149301337, 944629.149301337, 944629.149301337, 
    944629.149301337, 944629.149301337, 944629.149301337, 944629.149301337, 
    944629.149301337, 944629.149301337, 944629.149301337, 944629.149301337, 
    944629.149301337, 944629.149301337, 944629.149301337, 944629.149301337, 
    944629.149301337, 944629.149301337, 944629.149301337, 944629.149301337, 
    944629.149301337, 944629.149301337, 944629.149301337, 944629.149301337, 
    944629.149301337, 944629.149301337, 944629.149301337, 944629.149301337, 
    944629.149301337, 944629.149301337, 944629.149301337, 944629.149301337, 
    944629.149301337, 944629.149301337, 944629.149301337, 944629.149301337, 
    944629.149301337, 944629.149301337, 944629.149301337, 944629.149301337, 
    944629.149301337, 944629.149301337, 944629.149301337,
  981673.429666096, 981673.429666096, 981673.429666096, 981673.429666096, 
    981673.429666096, 981673.429666096, 981673.429666096, 981673.429666096, 
    981673.429666096, 981673.429666096, 981673.429666096, 981673.429666096, 
    981673.429666096, 981673.429666096, 981673.429666096, 981673.429666096, 
    981673.429666096, 981673.429666096, 981673.429666096, 981673.429666096, 
    981673.429666096, 981673.429666096, 981673.429666096, 981673.429666096, 
    981673.429666096, 981673.429666096, 981673.429666096, 981673.429666096, 
    981673.429666096, 981673.429666096, 981673.429666096, 981673.429666096, 
    981673.429666096, 981673.429666096, 981673.429666096, 981673.429666096, 
    981673.429666096, 981673.429666096, 981673.429666096, 981673.429666096, 
    981673.429666096, 981673.429666096, 981673.429666096, 981673.429666096, 
    981673.429666096, 981673.429666096, 981673.429666096, 981673.429666096, 
    981673.429666096, 981673.429666096, 981673.429666096, 981673.429666096, 
    981673.429666096, 981673.429666096, 981673.429666096,
  1018717.71003085, 1018717.71003085, 1018717.71003085, 1018717.71003085, 
    1018717.71003085, 1018717.71003085, 1018717.71003085, 1018717.71003085, 
    1018717.71003085, 1018717.71003085, 1018717.71003085, 1018717.71003085, 
    1018717.71003085, 1018717.71003085, 1018717.71003085, 1018717.71003085, 
    1018717.71003085, 1018717.71003085, 1018717.71003085, 1018717.71003085, 
    1018717.71003085, 1018717.71003085, 1018717.71003085, 1018717.71003085, 
    1018717.71003085, 1018717.71003085, 1018717.71003085, 1018717.71003085, 
    1018717.71003085, 1018717.71003085, 1018717.71003085, 1018717.71003085, 
    1018717.71003085, 1018717.71003085, 1018717.71003085, 1018717.71003085, 
    1018717.71003085, 1018717.71003085, 1018717.71003085, 1018717.71003085, 
    1018717.71003085, 1018717.71003085, 1018717.71003085, 1018717.71003085, 
    1018717.71003085, 1018717.71003085, 1018717.71003085, 1018717.71003085, 
    1018717.71003085, 1018717.71003085, 1018717.71003085, 1018717.71003085, 
    1018717.71003085, 1018717.71003085, 1018717.71003085,
  1055761.99039561, 1055761.99039561, 1055761.99039561, 1055761.99039561, 
    1055761.99039561, 1055761.99039561, 1055761.99039561, 1055761.99039561, 
    1055761.99039561, 1055761.99039561, 1055761.99039561, 1055761.99039561, 
    1055761.99039561, 1055761.99039561, 1055761.99039561, 1055761.99039561, 
    1055761.99039561, 1055761.99039561, 1055761.99039561, 1055761.99039561, 
    1055761.99039561, 1055761.99039561, 1055761.99039561, 1055761.99039561, 
    1055761.99039561, 1055761.99039561, 1055761.99039561, 1055761.99039561, 
    1055761.99039561, 1055761.99039561, 1055761.99039561, 1055761.99039561, 
    1055761.99039561, 1055761.99039561, 1055761.99039561, 1055761.99039561, 
    1055761.99039561, 1055761.99039561, 1055761.99039561, 1055761.99039561, 
    1055761.99039561, 1055761.99039561, 1055761.99039561, 1055761.99039561, 
    1055761.99039561, 1055761.99039561, 1055761.99039561, 1055761.99039561, 
    1055761.99039561, 1055761.99039561, 1055761.99039561, 1055761.99039561, 
    1055761.99039561, 1055761.99039561, 1055761.99039561,
  1092806.27076037, 1092806.27076037, 1092806.27076037, 1092806.27076037, 
    1092806.27076037, 1092806.27076037, 1092806.27076037, 1092806.27076037, 
    1092806.27076037, 1092806.27076037, 1092806.27076037, 1092806.27076037, 
    1092806.27076037, 1092806.27076037, 1092806.27076037, 1092806.27076037, 
    1092806.27076037, 1092806.27076037, 1092806.27076037, 1092806.27076037, 
    1092806.27076037, 1092806.27076037, 1092806.27076037, 1092806.27076037, 
    1092806.27076037, 1092806.27076037, 1092806.27076037, 1092806.27076037, 
    1092806.27076037, 1092806.27076037, 1092806.27076037, 1092806.27076037, 
    1092806.27076037, 1092806.27076037, 1092806.27076037, 1092806.27076037, 
    1092806.27076037, 1092806.27076037, 1092806.27076037, 1092806.27076037, 
    1092806.27076037, 1092806.27076037, 1092806.27076037, 1092806.27076037, 
    1092806.27076037, 1092806.27076037, 1092806.27076037, 1092806.27076037, 
    1092806.27076037, 1092806.27076037, 1092806.27076037, 1092806.27076037, 
    1092806.27076037, 1092806.27076037, 1092806.27076037,
  1129850.55112513, 1129850.55112513, 1129850.55112513, 1129850.55112513, 
    1129850.55112513, 1129850.55112513, 1129850.55112513, 1129850.55112513, 
    1129850.55112513, 1129850.55112513, 1129850.55112513, 1129850.55112513, 
    1129850.55112513, 1129850.55112513, 1129850.55112513, 1129850.55112513, 
    1129850.55112513, 1129850.55112513, 1129850.55112513, 1129850.55112513, 
    1129850.55112513, 1129850.55112513, 1129850.55112513, 1129850.55112513, 
    1129850.55112513, 1129850.55112513, 1129850.55112513, 1129850.55112513, 
    1129850.55112513, 1129850.55112513, 1129850.55112513, 1129850.55112513, 
    1129850.55112513, 1129850.55112513, 1129850.55112513, 1129850.55112513, 
    1129850.55112513, 1129850.55112513, 1129850.55112513, 1129850.55112513, 
    1129850.55112513, 1129850.55112513, 1129850.55112513, 1129850.55112513, 
    1129850.55112513, 1129850.55112513, 1129850.55112513, 1129850.55112513, 
    1129850.55112513, 1129850.55112513, 1129850.55112513, 1129850.55112513, 
    1129850.55112513, 1129850.55112513, 1129850.55112513,
  1166894.83148989, 1166894.83148989, 1166894.83148989, 1166894.83148989, 
    1166894.83148989, 1166894.83148989, 1166894.83148989, 1166894.83148989, 
    1166894.83148989, 1166894.83148989, 1166894.83148989, 1166894.83148989, 
    1166894.83148989, 1166894.83148989, 1166894.83148989, 1166894.83148989, 
    1166894.83148989, 1166894.83148989, 1166894.83148989, 1166894.83148989, 
    1166894.83148989, 1166894.83148989, 1166894.83148989, 1166894.83148989, 
    1166894.83148989, 1166894.83148989, 1166894.83148989, 1166894.83148989, 
    1166894.83148989, 1166894.83148989, 1166894.83148989, 1166894.83148989, 
    1166894.83148989, 1166894.83148989, 1166894.83148989, 1166894.83148989, 
    1166894.83148989, 1166894.83148989, 1166894.83148989, 1166894.83148989, 
    1166894.83148989, 1166894.83148989, 1166894.83148989, 1166894.83148989, 
    1166894.83148989, 1166894.83148989, 1166894.83148989, 1166894.83148989, 
    1166894.83148989, 1166894.83148989, 1166894.83148989, 1166894.83148989, 
    1166894.83148989, 1166894.83148989, 1166894.83148989,
  1203939.11185465, 1203939.11185465, 1203939.11185465, 1203939.11185465, 
    1203939.11185465, 1203939.11185465, 1203939.11185465, 1203939.11185465, 
    1203939.11185465, 1203939.11185465, 1203939.11185465, 1203939.11185465, 
    1203939.11185465, 1203939.11185465, 1203939.11185465, 1203939.11185465, 
    1203939.11185465, 1203939.11185465, 1203939.11185465, 1203939.11185465, 
    1203939.11185465, 1203939.11185465, 1203939.11185465, 1203939.11185465, 
    1203939.11185465, 1203939.11185465, 1203939.11185465, 1203939.11185465, 
    1203939.11185465, 1203939.11185465, 1203939.11185465, 1203939.11185465, 
    1203939.11185465, 1203939.11185465, 1203939.11185465, 1203939.11185465, 
    1203939.11185465, 1203939.11185465, 1203939.11185465, 1203939.11185465, 
    1203939.11185465, 1203939.11185465, 1203939.11185465, 1203939.11185465, 
    1203939.11185465, 1203939.11185465, 1203939.11185465, 1203939.11185465, 
    1203939.11185465, 1203939.11185465, 1203939.11185465, 1203939.11185465, 
    1203939.11185465, 1203939.11185465, 1203939.11185465,
  1240983.3922194, 1240983.3922194, 1240983.3922194, 1240983.3922194, 
    1240983.3922194, 1240983.3922194, 1240983.3922194, 1240983.3922194, 
    1240983.3922194, 1240983.3922194, 1240983.3922194, 1240983.3922194, 
    1240983.3922194, 1240983.3922194, 1240983.3922194, 1240983.3922194, 
    1240983.3922194, 1240983.3922194, 1240983.3922194, 1240983.3922194, 
    1240983.3922194, 1240983.3922194, 1240983.3922194, 1240983.3922194, 
    1240983.3922194, 1240983.3922194, 1240983.3922194, 1240983.3922194, 
    1240983.3922194, 1240983.3922194, 1240983.3922194, 1240983.3922194, 
    1240983.3922194, 1240983.3922194, 1240983.3922194, 1240983.3922194, 
    1240983.3922194, 1240983.3922194, 1240983.3922194, 1240983.3922194, 
    1240983.3922194, 1240983.3922194, 1240983.3922194, 1240983.3922194, 
    1240983.3922194, 1240983.3922194, 1240983.3922194, 1240983.3922194, 
    1240983.3922194, 1240983.3922194, 1240983.3922194, 1240983.3922194, 
    1240983.3922194, 1240983.3922194, 1240983.3922194,
  1278027.67258416, 1278027.67258416, 1278027.67258416, 1278027.67258416, 
    1278027.67258416, 1278027.67258416, 1278027.67258416, 1278027.67258416, 
    1278027.67258416, 1278027.67258416, 1278027.67258416, 1278027.67258416, 
    1278027.67258416, 1278027.67258416, 1278027.67258416, 1278027.67258416, 
    1278027.67258416, 1278027.67258416, 1278027.67258416, 1278027.67258416, 
    1278027.67258416, 1278027.67258416, 1278027.67258416, 1278027.67258416, 
    1278027.67258416, 1278027.67258416, 1278027.67258416, 1278027.67258416, 
    1278027.67258416, 1278027.67258416, 1278027.67258416, 1278027.67258416, 
    1278027.67258416, 1278027.67258416, 1278027.67258416, 1278027.67258416, 
    1278027.67258416, 1278027.67258416, 1278027.67258416, 1278027.67258416, 
    1278027.67258416, 1278027.67258416, 1278027.67258416, 1278027.67258416, 
    1278027.67258416, 1278027.67258416, 1278027.67258416, 1278027.67258416, 
    1278027.67258416, 1278027.67258416, 1278027.67258416, 1278027.67258416, 
    1278027.67258416, 1278027.67258416, 1278027.67258416,
  1315071.95294892, 1315071.95294892, 1315071.95294892, 1315071.95294892, 
    1315071.95294892, 1315071.95294892, 1315071.95294892, 1315071.95294892, 
    1315071.95294892, 1315071.95294892, 1315071.95294892, 1315071.95294892, 
    1315071.95294892, 1315071.95294892, 1315071.95294892, 1315071.95294892, 
    1315071.95294892, 1315071.95294892, 1315071.95294892, 1315071.95294892, 
    1315071.95294892, 1315071.95294892, 1315071.95294892, 1315071.95294892, 
    1315071.95294892, 1315071.95294892, 1315071.95294892, 1315071.95294892, 
    1315071.95294892, 1315071.95294892, 1315071.95294892, 1315071.95294892, 
    1315071.95294892, 1315071.95294892, 1315071.95294892, 1315071.95294892, 
    1315071.95294892, 1315071.95294892, 1315071.95294892, 1315071.95294892, 
    1315071.95294892, 1315071.95294892, 1315071.95294892, 1315071.95294892, 
    1315071.95294892, 1315071.95294892, 1315071.95294892, 1315071.95294892, 
    1315071.95294892, 1315071.95294892, 1315071.95294892, 1315071.95294892, 
    1315071.95294892, 1315071.95294892, 1315071.95294892,
  1352116.23331368, 1352116.23331368, 1352116.23331368, 1352116.23331368, 
    1352116.23331368, 1352116.23331368, 1352116.23331368, 1352116.23331368, 
    1352116.23331368, 1352116.23331368, 1352116.23331368, 1352116.23331368, 
    1352116.23331368, 1352116.23331368, 1352116.23331368, 1352116.23331368, 
    1352116.23331368, 1352116.23331368, 1352116.23331368, 1352116.23331368, 
    1352116.23331368, 1352116.23331368, 1352116.23331368, 1352116.23331368, 
    1352116.23331368, 1352116.23331368, 1352116.23331368, 1352116.23331368, 
    1352116.23331368, 1352116.23331368, 1352116.23331368, 1352116.23331368, 
    1352116.23331368, 1352116.23331368, 1352116.23331368, 1352116.23331368, 
    1352116.23331368, 1352116.23331368, 1352116.23331368, 1352116.23331368, 
    1352116.23331368, 1352116.23331368, 1352116.23331368, 1352116.23331368, 
    1352116.23331368, 1352116.23331368, 1352116.23331368, 1352116.23331368, 
    1352116.23331368, 1352116.23331368, 1352116.23331368, 1352116.23331368, 
    1352116.23331368, 1352116.23331368, 1352116.23331368,
  1389160.51367844, 1389160.51367844, 1389160.51367844, 1389160.51367844, 
    1389160.51367844, 1389160.51367844, 1389160.51367844, 1389160.51367844, 
    1389160.51367844, 1389160.51367844, 1389160.51367844, 1389160.51367844, 
    1389160.51367844, 1389160.51367844, 1389160.51367844, 1389160.51367844, 
    1389160.51367844, 1389160.51367844, 1389160.51367844, 1389160.51367844, 
    1389160.51367844, 1389160.51367844, 1389160.51367844, 1389160.51367844, 
    1389160.51367844, 1389160.51367844, 1389160.51367844, 1389160.51367844, 
    1389160.51367844, 1389160.51367844, 1389160.51367844, 1389160.51367844, 
    1389160.51367844, 1389160.51367844, 1389160.51367844, 1389160.51367844, 
    1389160.51367844, 1389160.51367844, 1389160.51367844, 1389160.51367844, 
    1389160.51367844, 1389160.51367844, 1389160.51367844, 1389160.51367844, 
    1389160.51367844, 1389160.51367844, 1389160.51367844, 1389160.51367844, 
    1389160.51367844, 1389160.51367844, 1389160.51367844, 1389160.51367844, 
    1389160.51367844, 1389160.51367844, 1389160.51367844,
  1426204.7940432, 1426204.7940432, 1426204.7940432, 1426204.7940432, 
    1426204.7940432, 1426204.7940432, 1426204.7940432, 1426204.7940432, 
    1426204.7940432, 1426204.7940432, 1426204.7940432, 1426204.7940432, 
    1426204.7940432, 1426204.7940432, 1426204.7940432, 1426204.7940432, 
    1426204.7940432, 1426204.7940432, 1426204.7940432, 1426204.7940432, 
    1426204.7940432, 1426204.7940432, 1426204.7940432, 1426204.7940432, 
    1426204.7940432, 1426204.7940432, 1426204.7940432, 1426204.7940432, 
    1426204.7940432, 1426204.7940432, 1426204.7940432, 1426204.7940432, 
    1426204.7940432, 1426204.7940432, 1426204.7940432, 1426204.7940432, 
    1426204.7940432, 1426204.7940432, 1426204.7940432, 1426204.7940432, 
    1426204.7940432, 1426204.7940432, 1426204.7940432, 1426204.7940432, 
    1426204.7940432, 1426204.7940432, 1426204.7940432, 1426204.7940432, 
    1426204.7940432, 1426204.7940432, 1426204.7940432, 1426204.7940432, 
    1426204.7940432, 1426204.7940432, 1426204.7940432,
  1463249.07440796, 1463249.07440796, 1463249.07440796, 1463249.07440796, 
    1463249.07440796, 1463249.07440796, 1463249.07440796, 1463249.07440796, 
    1463249.07440796, 1463249.07440796, 1463249.07440796, 1463249.07440796, 
    1463249.07440796, 1463249.07440796, 1463249.07440796, 1463249.07440796, 
    1463249.07440796, 1463249.07440796, 1463249.07440796, 1463249.07440796, 
    1463249.07440796, 1463249.07440796, 1463249.07440796, 1463249.07440796, 
    1463249.07440796, 1463249.07440796, 1463249.07440796, 1463249.07440796, 
    1463249.07440796, 1463249.07440796, 1463249.07440796, 1463249.07440796, 
    1463249.07440796, 1463249.07440796, 1463249.07440796, 1463249.07440796, 
    1463249.07440796, 1463249.07440796, 1463249.07440796, 1463249.07440796, 
    1463249.07440796, 1463249.07440796, 1463249.07440796, 1463249.07440796, 
    1463249.07440796, 1463249.07440796, 1463249.07440796, 1463249.07440796, 
    1463249.07440796, 1463249.07440796, 1463249.07440796, 1463249.07440796, 
    1463249.07440796, 1463249.07440796, 1463249.07440796,
  1500293.35477271, 1500293.35477271, 1500293.35477271, 1500293.35477271, 
    1500293.35477271, 1500293.35477271, 1500293.35477271, 1500293.35477271, 
    1500293.35477271, 1500293.35477271, 1500293.35477271, 1500293.35477271, 
    1500293.35477271, 1500293.35477271, 1500293.35477271, 1500293.35477271, 
    1500293.35477271, 1500293.35477271, 1500293.35477271, 1500293.35477271, 
    1500293.35477271, 1500293.35477271, 1500293.35477271, 1500293.35477271, 
    1500293.35477271, 1500293.35477271, 1500293.35477271, 1500293.35477271, 
    1500293.35477271, 1500293.35477271, 1500293.35477271, 1500293.35477271, 
    1500293.35477271, 1500293.35477271, 1500293.35477271, 1500293.35477271, 
    1500293.35477271, 1500293.35477271, 1500293.35477271, 1500293.35477271, 
    1500293.35477271, 1500293.35477271, 1500293.35477271, 1500293.35477271, 
    1500293.35477271, 1500293.35477271, 1500293.35477271, 1500293.35477271, 
    1500293.35477271, 1500293.35477271, 1500293.35477271, 1500293.35477271, 
    1500293.35477271, 1500293.35477271, 1500293.35477271,
  1537337.63513747, 1537337.63513747, 1537337.63513747, 1537337.63513747, 
    1537337.63513747, 1537337.63513747, 1537337.63513747, 1537337.63513747, 
    1537337.63513747, 1537337.63513747, 1537337.63513747, 1537337.63513747, 
    1537337.63513747, 1537337.63513747, 1537337.63513747, 1537337.63513747, 
    1537337.63513747, 1537337.63513747, 1537337.63513747, 1537337.63513747, 
    1537337.63513747, 1537337.63513747, 1537337.63513747, 1537337.63513747, 
    1537337.63513747, 1537337.63513747, 1537337.63513747, 1537337.63513747, 
    1537337.63513747, 1537337.63513747, 1537337.63513747, 1537337.63513747, 
    1537337.63513747, 1537337.63513747, 1537337.63513747, 1537337.63513747, 
    1537337.63513747, 1537337.63513747, 1537337.63513747, 1537337.63513747, 
    1537337.63513747, 1537337.63513747, 1537337.63513747, 1537337.63513747, 
    1537337.63513747, 1537337.63513747, 1537337.63513747, 1537337.63513747, 
    1537337.63513747, 1537337.63513747, 1537337.63513747, 1537337.63513747, 
    1537337.63513747, 1537337.63513747, 1537337.63513747,
  1574381.91550223, 1574381.91550223, 1574381.91550223, 1574381.91550223, 
    1574381.91550223, 1574381.91550223, 1574381.91550223, 1574381.91550223, 
    1574381.91550223, 1574381.91550223, 1574381.91550223, 1574381.91550223, 
    1574381.91550223, 1574381.91550223, 1574381.91550223, 1574381.91550223, 
    1574381.91550223, 1574381.91550223, 1574381.91550223, 1574381.91550223, 
    1574381.91550223, 1574381.91550223, 1574381.91550223, 1574381.91550223, 
    1574381.91550223, 1574381.91550223, 1574381.91550223, 1574381.91550223, 
    1574381.91550223, 1574381.91550223, 1574381.91550223, 1574381.91550223, 
    1574381.91550223, 1574381.91550223, 1574381.91550223, 1574381.91550223, 
    1574381.91550223, 1574381.91550223, 1574381.91550223, 1574381.91550223, 
    1574381.91550223, 1574381.91550223, 1574381.91550223, 1574381.91550223, 
    1574381.91550223, 1574381.91550223, 1574381.91550223, 1574381.91550223, 
    1574381.91550223, 1574381.91550223, 1574381.91550223, 1574381.91550223, 
    1574381.91550223, 1574381.91550223, 1574381.91550223,
  1611426.19586699, 1611426.19586699, 1611426.19586699, 1611426.19586699, 
    1611426.19586699, 1611426.19586699, 1611426.19586699, 1611426.19586699, 
    1611426.19586699, 1611426.19586699, 1611426.19586699, 1611426.19586699, 
    1611426.19586699, 1611426.19586699, 1611426.19586699, 1611426.19586699, 
    1611426.19586699, 1611426.19586699, 1611426.19586699, 1611426.19586699, 
    1611426.19586699, 1611426.19586699, 1611426.19586699, 1611426.19586699, 
    1611426.19586699, 1611426.19586699, 1611426.19586699, 1611426.19586699, 
    1611426.19586699, 1611426.19586699, 1611426.19586699, 1611426.19586699, 
    1611426.19586699, 1611426.19586699, 1611426.19586699, 1611426.19586699, 
    1611426.19586699, 1611426.19586699, 1611426.19586699, 1611426.19586699, 
    1611426.19586699, 1611426.19586699, 1611426.19586699, 1611426.19586699, 
    1611426.19586699, 1611426.19586699, 1611426.19586699, 1611426.19586699, 
    1611426.19586699, 1611426.19586699, 1611426.19586699, 1611426.19586699, 
    1611426.19586699, 1611426.19586699, 1611426.19586699,
  1648470.47623175, 1648470.47623175, 1648470.47623175, 1648470.47623175, 
    1648470.47623175, 1648470.47623175, 1648470.47623175, 1648470.47623175, 
    1648470.47623175, 1648470.47623175, 1648470.47623175, 1648470.47623175, 
    1648470.47623175, 1648470.47623175, 1648470.47623175, 1648470.47623175, 
    1648470.47623175, 1648470.47623175, 1648470.47623175, 1648470.47623175, 
    1648470.47623175, 1648470.47623175, 1648470.47623175, 1648470.47623175, 
    1648470.47623175, 1648470.47623175, 1648470.47623175, 1648470.47623175, 
    1648470.47623175, 1648470.47623175, 1648470.47623175, 1648470.47623175, 
    1648470.47623175, 1648470.47623175, 1648470.47623175, 1648470.47623175, 
    1648470.47623175, 1648470.47623175, 1648470.47623175, 1648470.47623175, 
    1648470.47623175, 1648470.47623175, 1648470.47623175, 1648470.47623175, 
    1648470.47623175, 1648470.47623175, 1648470.47623175, 1648470.47623175, 
    1648470.47623175, 1648470.47623175, 1648470.47623175, 1648470.47623175, 
    1648470.47623175, 1648470.47623175, 1648470.47623175,
  1685514.75659651, 1685514.75659651, 1685514.75659651, 1685514.75659651, 
    1685514.75659651, 1685514.75659651, 1685514.75659651, 1685514.75659651, 
    1685514.75659651, 1685514.75659651, 1685514.75659651, 1685514.75659651, 
    1685514.75659651, 1685514.75659651, 1685514.75659651, 1685514.75659651, 
    1685514.75659651, 1685514.75659651, 1685514.75659651, 1685514.75659651, 
    1685514.75659651, 1685514.75659651, 1685514.75659651, 1685514.75659651, 
    1685514.75659651, 1685514.75659651, 1685514.75659651, 1685514.75659651, 
    1685514.75659651, 1685514.75659651, 1685514.75659651, 1685514.75659651, 
    1685514.75659651, 1685514.75659651, 1685514.75659651, 1685514.75659651, 
    1685514.75659651, 1685514.75659651, 1685514.75659651, 1685514.75659651, 
    1685514.75659651, 1685514.75659651, 1685514.75659651, 1685514.75659651, 
    1685514.75659651, 1685514.75659651, 1685514.75659651, 1685514.75659651, 
    1685514.75659651, 1685514.75659651, 1685514.75659651, 1685514.75659651, 
    1685514.75659651, 1685514.75659651, 1685514.75659651,
  1722559.03696126, 1722559.03696126, 1722559.03696126, 1722559.03696126, 
    1722559.03696126, 1722559.03696126, 1722559.03696126, 1722559.03696126, 
    1722559.03696126, 1722559.03696126, 1722559.03696126, 1722559.03696126, 
    1722559.03696126, 1722559.03696126, 1722559.03696126, 1722559.03696126, 
    1722559.03696126, 1722559.03696126, 1722559.03696126, 1722559.03696126, 
    1722559.03696126, 1722559.03696126, 1722559.03696126, 1722559.03696126, 
    1722559.03696126, 1722559.03696126, 1722559.03696126, 1722559.03696126, 
    1722559.03696126, 1722559.03696126, 1722559.03696126, 1722559.03696126, 
    1722559.03696126, 1722559.03696126, 1722559.03696126, 1722559.03696126, 
    1722559.03696126, 1722559.03696126, 1722559.03696126, 1722559.03696126, 
    1722559.03696126, 1722559.03696126, 1722559.03696126, 1722559.03696126, 
    1722559.03696126, 1722559.03696126, 1722559.03696126, 1722559.03696126, 
    1722559.03696126, 1722559.03696126, 1722559.03696126, 1722559.03696126, 
    1722559.03696126, 1722559.03696126, 1722559.03696126,
  1759603.31732602, 1759603.31732602, 1759603.31732602, 1759603.31732602, 
    1759603.31732602, 1759603.31732602, 1759603.31732602, 1759603.31732602, 
    1759603.31732602, 1759603.31732602, 1759603.31732602, 1759603.31732602, 
    1759603.31732602, 1759603.31732602, 1759603.31732602, 1759603.31732602, 
    1759603.31732602, 1759603.31732602, 1759603.31732602, 1759603.31732602, 
    1759603.31732602, 1759603.31732602, 1759603.31732602, 1759603.31732602, 
    1759603.31732602, 1759603.31732602, 1759603.31732602, 1759603.31732602, 
    1759603.31732602, 1759603.31732602, 1759603.31732602, 1759603.31732602, 
    1759603.31732602, 1759603.31732602, 1759603.31732602, 1759603.31732602, 
    1759603.31732602, 1759603.31732602, 1759603.31732602, 1759603.31732602, 
    1759603.31732602, 1759603.31732602, 1759603.31732602, 1759603.31732602, 
    1759603.31732602, 1759603.31732602, 1759603.31732602, 1759603.31732602, 
    1759603.31732602, 1759603.31732602, 1759603.31732602, 1759603.31732602, 
    1759603.31732602, 1759603.31732602, 1759603.31732602,
  1796647.59769078, 1796647.59769078, 1796647.59769078, 1796647.59769078, 
    1796647.59769078, 1796647.59769078, 1796647.59769078, 1796647.59769078, 
    1796647.59769078, 1796647.59769078, 1796647.59769078, 1796647.59769078, 
    1796647.59769078, 1796647.59769078, 1796647.59769078, 1796647.59769078, 
    1796647.59769078, 1796647.59769078, 1796647.59769078, 1796647.59769078, 
    1796647.59769078, 1796647.59769078, 1796647.59769078, 1796647.59769078, 
    1796647.59769078, 1796647.59769078, 1796647.59769078, 1796647.59769078, 
    1796647.59769078, 1796647.59769078, 1796647.59769078, 1796647.59769078, 
    1796647.59769078, 1796647.59769078, 1796647.59769078, 1796647.59769078, 
    1796647.59769078, 1796647.59769078, 1796647.59769078, 1796647.59769078, 
    1796647.59769078, 1796647.59769078, 1796647.59769078, 1796647.59769078, 
    1796647.59769078, 1796647.59769078, 1796647.59769078, 1796647.59769078, 
    1796647.59769078, 1796647.59769078, 1796647.59769078, 1796647.59769078, 
    1796647.59769078, 1796647.59769078, 1796647.59769078,
  1833691.87805554, 1833691.87805554, 1833691.87805554, 1833691.87805554, 
    1833691.87805554, 1833691.87805554, 1833691.87805554, 1833691.87805554, 
    1833691.87805554, 1833691.87805554, 1833691.87805554, 1833691.87805554, 
    1833691.87805554, 1833691.87805554, 1833691.87805554, 1833691.87805554, 
    1833691.87805554, 1833691.87805554, 1833691.87805554, 1833691.87805554, 
    1833691.87805554, 1833691.87805554, 1833691.87805554, 1833691.87805554, 
    1833691.87805554, 1833691.87805554, 1833691.87805554, 1833691.87805554, 
    1833691.87805554, 1833691.87805554, 1833691.87805554, 1833691.87805554, 
    1833691.87805554, 1833691.87805554, 1833691.87805554, 1833691.87805554, 
    1833691.87805554, 1833691.87805554, 1833691.87805554, 1833691.87805554, 
    1833691.87805554, 1833691.87805554, 1833691.87805554, 1833691.87805554, 
    1833691.87805554, 1833691.87805554, 1833691.87805554, 1833691.87805554, 
    1833691.87805554, 1833691.87805554, 1833691.87805554, 1833691.87805554, 
    1833691.87805554, 1833691.87805554, 1833691.87805554,
  1870736.1584203, 1870736.1584203, 1870736.1584203, 1870736.1584203, 
    1870736.1584203, 1870736.1584203, 1870736.1584203, 1870736.1584203, 
    1870736.1584203, 1870736.1584203, 1870736.1584203, 1870736.1584203, 
    1870736.1584203, 1870736.1584203, 1870736.1584203, 1870736.1584203, 
    1870736.1584203, 1870736.1584203, 1870736.1584203, 1870736.1584203, 
    1870736.1584203, 1870736.1584203, 1870736.1584203, 1870736.1584203, 
    1870736.1584203, 1870736.1584203, 1870736.1584203, 1870736.1584203, 
    1870736.1584203, 1870736.1584203, 1870736.1584203, 1870736.1584203, 
    1870736.1584203, 1870736.1584203, 1870736.1584203, 1870736.1584203, 
    1870736.1584203, 1870736.1584203, 1870736.1584203, 1870736.1584203, 
    1870736.1584203, 1870736.1584203, 1870736.1584203, 1870736.1584203, 
    1870736.1584203, 1870736.1584203, 1870736.1584203, 1870736.1584203, 
    1870736.1584203, 1870736.1584203, 1870736.1584203, 1870736.1584203, 
    1870736.1584203, 1870736.1584203, 1870736.1584203,
  1907780.43878506, 1907780.43878506, 1907780.43878506, 1907780.43878506, 
    1907780.43878506, 1907780.43878506, 1907780.43878506, 1907780.43878506, 
    1907780.43878506, 1907780.43878506, 1907780.43878506, 1907780.43878506, 
    1907780.43878506, 1907780.43878506, 1907780.43878506, 1907780.43878506, 
    1907780.43878506, 1907780.43878506, 1907780.43878506, 1907780.43878506, 
    1907780.43878506, 1907780.43878506, 1907780.43878506, 1907780.43878506, 
    1907780.43878506, 1907780.43878506, 1907780.43878506, 1907780.43878506, 
    1907780.43878506, 1907780.43878506, 1907780.43878506, 1907780.43878506, 
    1907780.43878506, 1907780.43878506, 1907780.43878506, 1907780.43878506, 
    1907780.43878506, 1907780.43878506, 1907780.43878506, 1907780.43878506, 
    1907780.43878506, 1907780.43878506, 1907780.43878506, 1907780.43878506, 
    1907780.43878506, 1907780.43878506, 1907780.43878506, 1907780.43878506, 
    1907780.43878506, 1907780.43878506, 1907780.43878506, 1907780.43878506, 
    1907780.43878506, 1907780.43878506, 1907780.43878506,
  1944824.71914981, 1944824.71914981, 1944824.71914981, 1944824.71914981, 
    1944824.71914981, 1944824.71914981, 1944824.71914981, 1944824.71914981, 
    1944824.71914981, 1944824.71914981, 1944824.71914981, 1944824.71914981, 
    1944824.71914981, 1944824.71914981, 1944824.71914981, 1944824.71914981, 
    1944824.71914981, 1944824.71914981, 1944824.71914981, 1944824.71914981, 
    1944824.71914981, 1944824.71914981, 1944824.71914981, 1944824.71914981, 
    1944824.71914981, 1944824.71914981, 1944824.71914981, 1944824.71914981, 
    1944824.71914981, 1944824.71914981, 1944824.71914981, 1944824.71914981, 
    1944824.71914981, 1944824.71914981, 1944824.71914981, 1944824.71914981, 
    1944824.71914981, 1944824.71914981, 1944824.71914981, 1944824.71914981, 
    1944824.71914981, 1944824.71914981, 1944824.71914981, 1944824.71914981, 
    1944824.71914981, 1944824.71914981, 1944824.71914981, 1944824.71914981, 
    1944824.71914981, 1944824.71914981, 1944824.71914981, 1944824.71914981, 
    1944824.71914981, 1944824.71914981, 1944824.71914981,
  1981868.99951457, 1981868.99951457, 1981868.99951457, 1981868.99951457, 
    1981868.99951457, 1981868.99951457, 1981868.99951457, 1981868.99951457, 
    1981868.99951457, 1981868.99951457, 1981868.99951457, 1981868.99951457, 
    1981868.99951457, 1981868.99951457, 1981868.99951457, 1981868.99951457, 
    1981868.99951457, 1981868.99951457, 1981868.99951457, 1981868.99951457, 
    1981868.99951457, 1981868.99951457, 1981868.99951457, 1981868.99951457, 
    1981868.99951457, 1981868.99951457, 1981868.99951457, 1981868.99951457, 
    1981868.99951457, 1981868.99951457, 1981868.99951457, 1981868.99951457, 
    1981868.99951457, 1981868.99951457, 1981868.99951457, 1981868.99951457, 
    1981868.99951457, 1981868.99951457, 1981868.99951457, 1981868.99951457, 
    1981868.99951457, 1981868.99951457, 1981868.99951457, 1981868.99951457, 
    1981868.99951457, 1981868.99951457, 1981868.99951457, 1981868.99951457, 
    1981868.99951457, 1981868.99951457, 1981868.99951457, 1981868.99951457, 
    1981868.99951457, 1981868.99951457, 1981868.99951457 ;

 lon_rho =
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667 ;

 lon_u =
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333 ;

 lon_v =
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667 ;

 lon_psi =
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333 ;

 lat_rho =
  30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30,
  30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333,
  30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667,
  31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 
    31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 
    31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31,
  31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333,
  31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667,
  32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 
    32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 
    32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32,
  32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333,
  32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667,
  33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 
    33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 
    33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33,
  33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333,
  33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667,
  34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 
    34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 
    34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34,
  34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333,
  34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333,
  35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667,
  36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 
    36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 
    36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36,
  36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333,
  36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667,
  37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 
    37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 
    37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37,
  37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333,
  37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667,
  38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 
    38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 
    38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38,
  38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333,
  38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667,
  39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 
    39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 
    39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39,
  39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333,
  39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667,
  40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 
    40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 
    40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40,
  40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333,
  40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667,
  41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 
    41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 
    41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41,
  41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333,
  41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667,
  42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 
    42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 
    42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42,
  42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333,
  42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667,
  43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 
    43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 
    43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43,
  43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333,
  43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667,
  44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 
    44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 
    44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44,
  44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333,
  44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667,
  45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 
    45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 
    45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45,
  45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333,
  45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667,
  46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 
    46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 
    46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46,
  46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333,
  46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667,
  47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 
    47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 
    47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47,
  47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333,
  47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667,
  48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 
    48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 
    48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48 ;

 lat_u =
  30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30,
  30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333,
  30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667,
  31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 
    31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 
    31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31,
  31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333,
  31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667,
  32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 
    32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 
    32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32,
  32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333,
  32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667,
  33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 
    33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 
    33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33,
  33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333,
  33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667,
  34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 
    34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 
    34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34,
  34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333,
  34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333,
  35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667,
  36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 
    36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 
    36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36,
  36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333,
  36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667,
  37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 
    37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 
    37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37,
  37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333,
  37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667,
  38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 
    38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 
    38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38,
  38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333,
  38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667,
  39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 
    39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 
    39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39,
  39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333,
  39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667,
  40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 
    40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 
    40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40,
  40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333,
  40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667,
  41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 
    41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 
    41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41,
  41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333,
  41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667,
  42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 
    42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 
    42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42,
  42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333,
  42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667,
  43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 
    43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 
    43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43,
  43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333,
  43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667,
  44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 
    44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 
    44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44,
  44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333,
  44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667,
  45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 
    45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 
    45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45,
  45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333,
  45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667,
  46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 
    46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 
    46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46,
  46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333,
  46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667,
  47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 
    47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 
    47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47,
  47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333,
  47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667,
  48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 
    48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 
    48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48 ;

 lat_v =
  30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667,
  30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 
    30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 
    30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 
    30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 
    30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5,
  30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333,
  31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667,
  31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 
    31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 
    31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 
    31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 
    31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5,
  31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333,
  32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667,
  32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 
    32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 
    32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 
    32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 
    32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5,
  32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333,
  33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667,
  33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 
    33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 
    33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 
    33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 
    33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5,
  33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333,
  34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667,
  34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 
    34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 
    34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 
    34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 
    34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5,
  34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333,
  35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667,
  35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 
    35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 
    35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 
    35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 
    35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5,
  35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333,
  36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667,
  36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 
    36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 
    36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 
    36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 
    36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5,
  36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333,
  37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667,
  37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 
    37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 
    37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 
    37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 
    37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5,
  37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333,
  38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667,
  38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 
    38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 
    38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 
    38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 
    38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5,
  38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333,
  39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667,
  39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 
    39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 
    39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 
    39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 
    39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5,
  39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333,
  40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667,
  40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 
    40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 
    40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 
    40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 
    40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5,
  40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333,
  41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667,
  41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 
    41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 
    41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 
    41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 
    41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5,
  41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333,
  42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667,
  42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 
    42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 
    42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 
    42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 
    42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5,
  42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333,
  43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667,
  43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 
    43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 
    43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 
    43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 
    43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5,
  43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333,
  44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667,
  44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 
    44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 
    44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 
    44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 
    44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5,
  44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333,
  45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667,
  45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 
    45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 
    45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 
    45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 
    45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5,
  45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333,
  46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667,
  46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 
    46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 
    46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 
    46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 
    46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5,
  46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333,
  47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667,
  47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 
    47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 
    47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 
    47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 
    47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5,
  47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333 ;

 lat_psi =
  30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667,
  30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 
    30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 
    30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 
    30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 
    30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5,
  30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333,
  31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667,
  31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 
    31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 
    31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 
    31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 
    31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5,
  31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333,
  32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667,
  32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 
    32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 
    32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 
    32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 
    32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5,
  32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333,
  33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667,
  33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 
    33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 
    33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 
    33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 
    33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5,
  33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333,
  34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667,
  34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 
    34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 
    34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 
    34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 
    34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5,
  34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333,
  35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667,
  35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 
    35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 
    35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 
    35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 
    35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5,
  35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333,
  36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667,
  36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 
    36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 
    36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 
    36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 
    36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5,
  36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333,
  37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667,
  37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 
    37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 
    37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 
    37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 
    37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5,
  37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333,
  38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667,
  38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 
    38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 
    38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 
    38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 
    38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5,
  38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333,
  39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667,
  39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 
    39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 
    39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 
    39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 
    39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5,
  39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333,
  40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667,
  40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 
    40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 
    40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 
    40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 
    40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5,
  40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333,
  41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667,
  41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 
    41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 
    41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 
    41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 
    41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5,
  41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333,
  42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667,
  42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 
    42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 
    42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 
    42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 
    42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5,
  42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333,
  43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667,
  43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 
    43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 
    43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 
    43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 
    43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5,
  43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333,
  44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667,
  44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 
    44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 
    44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 
    44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 
    44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5,
  44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333,
  45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667,
  45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 
    45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 
    45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 
    45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 
    45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5,
  45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333,
  46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667,
  46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 
    46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 
    46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 
    46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 
    46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5,
  46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333,
  47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667,
  47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 
    47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 
    47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 
    47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 
    47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5,
  47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333 ;

 mask_rho =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0 ;

 mask_u =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0 ;

 mask_v =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0 ;

 mask_psi =
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 
    1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0 ;

 lon_coast = NaN, -114, NaN, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114.002389, -114.01, -114.009444, -114.014639, -114.02925, 
    -114.030083, -114.032222, -114.035583, -114.031361, -114.014333, 
    -114.021833, -114.028667, -114.023667, -114.024611, -114.028417, 
    -114.032361, -114.026333, -114.034167, -114.033444, -114.025361, 
    -114.022028, -114.014972, -114.010333, -114.017139, -114.023111, 
    -114.022556, -114.0285, -114.044778, -114.06925, -114.132444, -114.15875, 
    -114.199361, -114.228722, -114.275833, -114.301694, -114.316361, 
    -114.327528, -114.329, -114.335694, -114.362222, -114.392444, 
    -114.416611, -114.432444, -114.446889, -114.45075, -114.451417, -114.466, 
    -114.495556, -114.496778, -114.513167, -114.510611, -114.532194, 
    -114.547028, -114.555056, -114.583333, -114.584722, -114.586833, 
    -114.617889, -114.676667, -114.689889, -114.709694, -114.755028, 
    -114.776111, -114.782694, -114.778402, -114.778972, -114.811361, 
    -114.830389, -114.840722, -114.85425, -114.902278, -114.915417, 
    -114.932528, -114.923917, -114.914556, -114.924639, -114.937444, 
    -114.95475, -114.9455, -114.931361, -114.9195, -114.907694, -114.896889, 
    -114.859778, -114.850917, -114.83925, -114.8485, -114.837972, 
    -114.828556, -114.838056, -114.846528, -114.851694, -114.887139, 
    -114.852917, -114.845806, -114.839361, -114.825389, -114.820917, 
    -114.823944, -114.790083, -114.784278, -114.782722, -114.785333, 
    -114.798083, -114.80925, -114.808722, -114.822111, -114.820222, 
    -114.830472, -114.832722, -114.843722, -114.851167, -114.858611, 
    -114.855111, -114.857833, -114.861306, -114.869611, -114.871861, 
    -114.881111, -114.882778, -114.88, -114.88325, -114.886278, -114.881972, 
    -114.883444, -114.887167, -114.88825, -114.900667, -114.888944, 
    -114.888611, -114.906806, -114.915389, -114.908639, -114.911806, 
    -114.897202, -114.887639, -114.898583, -114.892917, -114.886944, 
    -114.889333, -114.892139, -114.891889, -114.896194, -114.902694, 
    -114.906806, -114.904556, -114.893944, -114.894694, -114.915611, 
    -114.899528, -114.905833, -114.904472, -114.895139, -114.897639, 
    -114.903639, -114.900278, -114.913972, -114.909083, -114.919389, 
    -114.914222, -114.906778, -114.90925, -114.905333, -114.899556, 
    -114.907444, -114.899528, -114.899, -114.909, -114.898667, -114.909306, 
    -114.9, -114.908611, -114.902306, -114.897417, -114.896028, -114.900917, 
    -114.894833, -114.897667, -114.885111, -114.888556, -114.88775, 
    -114.891167, -114.890333, -114.890056, -114.886083, -114.88775, 
    -114.885361, -114.88325, -114.886806, -114.895667, -114.896722, 
    -114.899917, -114.903639, -114.90075, -114.893444, -114.885806, 
    -114.893444, -114.886583, -114.871306, -114.86375, -114.861028, 
    -114.849917, -114.834806, -114.824583, -114.817139, -114.8135, 
    -114.814333, -114.827139, -114.836056, -114.837556, -114.834667, 
    -114.827306, -114.811306, -114.721722, -114.712083, -114.707111, 
    -114.710639, -114.706639, -114.703167, -114.710056, -114.700556, 
    -114.701833, -114.699806, -114.696472, -114.70025, -114.697583, 
    -114.699917, -114.694028, -114.699028, -114.693972, -114.706111, 
    -114.694889, -114.698389, -114.677472, -114.665111, -114.660861, 
    -114.652361, -114.6525, -114.649028, -114.650806, -114.6315, -114.629806, 
    -114.632306, -114.638583, -114.637556, -114.630167, -114.642806, 
    -114.634972, -114.635889, -114.638528, -114.6425, -114.640028, 
    -114.645333, -114.645556, -114.652639, -114.6525, -114.656972, 
    -114.656639, -114.640861, -114.64, -114.652583, -114.650833, -114.653333, 
    -114.669111, -114.664083, -114.652583, -114.651111, -114.635639, 
    -114.634306, -114.629472, -114.607889, -114.596611, -114.586306, 
    -114.582444, -114.583722, -114.575833, -114.566889, -114.565694, 
    -114.552611, -114.538278, -114.532944, -114.508, -114.493194, 
    -114.486194, -114.471639, -114.447, -114.433611, -114.413639, 
    -114.410556, -114.414667, -114.400139, -114.394694, -114.397389, 
    -114.404056, -114.409056, -114.40875, -114.400139, -114.403278, 
    -114.400389, -114.397806, -114.393861, -114.393167, -114.397389, 
    -114.384194, -114.376111, -114.358861, -114.348111, -114.34175, 
    -114.331222, -114.309556, -114.303861, -114.302778, -114.297528, 
    -114.283028, -114.287083, -114.287722, -114.292222, -114.295083, 
    -114.294639, -114.286722, -114.284194, -114.273389, -114.265472, 
    -114.263639, -114.261306, -114.258972, -114.258833, -114.244833, 
    -114.228333, -114.207472, -114.200722, -114.179583, -114.166139, 
    -114.159889, -114.153306, -114.145083, -114.133111, -114.117667, 
    -114.109639, -114.080667, -114.064444, -114.046389, -114.031222, 
    -114.021778, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -115.048667, -115.054306, -115.083667, -115.078861, -115.058611, 
    -115.037444, -115.017583, -115.008528, -114.972806, -114.914944, 
    -114.879694, -114.866583, -114.852583, -114.85175, -114.844972, 
    -114.835417, -114.799056, -114.790472, -114.77225, -114.766694, 
    -114.727639, -114.717583, -114.718083, -114.438778, -114.4005, 
    -114.349417, -114.333361, -114.31925, -114.296, -114.292528, -114.294306, 
    -114.3035, -114.307667, -114.295111, -114.293556, -114.296944, 
    -114.302917, -114.30575, -114.305611, -114.300111, -114.29875, 
    -114.302556, -114.303778, -114.059694, -114.069139, -114.071944, 
    -114.069944, -114.176583, -114.179056, -114.169306, -114.167306, 
    -114.176556, -114.179694, -114.179861, -114.171444, -114.169556, 
    -114.143333, -114.141694, -114.135444, -114.134917, -114.132333, 
    -114.134139, -114.137167, -114.138361, -114.141806, -114.139972, 
    -114.155833, -114.15175, -114.133389, -114.160472, -114.177278, 
    -114.190083, -114.186611, -114.179778, -114.185083, -114.178556, 
    -114.174167, -114.173583, -114.178111, -114.171583, -114.175306, 
    -114.167306, -114.155833, -114.157333, -114.162556, -114.169056, 
    -114.168361, -114.160944, -114.164222, -114.169333, -114.166083, 
    -114.166306, -114.15775, -114.161861, -114.152694, -114.149167, 
    -114.152556, -114.147833, -114.147639, -114.151361, -114.150417, 
    -114.15425, -114.154583, -114.146944, -114.133833, -114.131472, 
    -114.135722, -114.140278, -114.143083, -114.139111, -114.144778, 
    -114.149389, -114.141306, -114.133417, -114.1275, -114.140111, 
    -114.163167, -114.158778, -114.166361, -114.165889, -114.162, 
    -114.156139, -114.154111, -114.161667, -114.170083, -114.181333, 
    -114.173722, -114.195972, -114.200056, -114.22025, -114.234278, 
    -114.244167, -114.257528, -114.266278, -114.272861, -114.277556, 
    -114.268972, -114.248472, -114.228556, -114.214389, -114.20944658715, 
    -114.18875, -114.139417, -114.132556, -114.121778, -114.115083, 
    -114.119167, -114.130417, -114.146028, -114.150972, -114.149194, 
    -114.148563156947, -114.128194, -114.128278, -114.135722, -114.139917, 
    -114.132611, -114.123944, -114.115694, -114.111167, -114.098611, 
    -114.098333, -114.093944, -114.096833, -114.087472, -114.089, 
    -114.098306, -114.096361, -114.10175, -114.092694, -114.0965, 
    -114.103917, -114.103917, -114.098361, -114.104722, -114.106889, 
    -114.117, -114.124972, -114.125861, -114.116694, -114.124278, 
    -114.120417, -114.094167, -114.093778, -114.09775, -114.102694, 
    -114.097583, -114.087389, -114.087667, -114.080889, -114.083944, -114.08, 
    -114.076008846858, -114.085833, -114.076889, -114.077611, -114.081722, 
    -114.078306, -114.078056, -114.073083, -114.066271379796, -114.040889, 
    -114.036167, -114.054778, -114.068361, -114.093861, -114.106389, 
    -114.104139, -114.116028, -114.113361, -114.087167, -114.072778, 
    -114.064028, -114.060056, -114.063556, -114.060972, -114.075278, 
    -114.075972, -114.075028, -114.068861, -114.066222, -114.067278, 
    -114.059083, -114.064417, -114.065222, -114.062778, -114.059333, 
    -114.056917, -114.067833, -114.064639, -114.067889, -114.063889, 
    -114.067056, -114.062944, -114.064056, -114.0605, -114.061167, 
    -114.054528, -114.050222, -114.045806, -114.051056, -114.051889, -114.06, 
    -114.065028, -114.070222, -114.073222, -114.076139, -114.076, -114.07275, 
    -114.076139, -114.073833, -114.080917, -114.086833, -114.08925, 
    -114.084778, -114.085583, -114.101528, -114.110694, -114.118611, 
    -114.127194, -114.083611, -114.063417, -114.052833, -114.0475, 
    -114.053417, -114.071389, -114.071722, -114.0675, -114.075361, 
    -114.086528, -114.097444, -114.116611, -114.131389, -114.147306, 
    -114.160833, -114.154861, -114.157611, -114.162694, -114.177389, 
    -114.224528, -114.243861, -114.246056, -114.259917, -114.270306, 
    -114.270111, -114.285056, -114.287889, -114.291167, -114.302028, 
    -114.307722, -114.314278, -114.346833, -114.349917, -114.346028, 
    -114.343583, -114.344417, -114.349028, -114.354222, -114.349056, 
    -114.350028, -114.361111, -114.362528, -114.376028, -114.379722, 
    -114.388056, -114.399389, -114.399444, -114.405, -114.407639, 
    -114.415528, -114.427861, -114.439194, -114.44175, -114.452222, 
    -114.462694, -114.473861, -114.491139, -114.504889, -114.51275, 
    -114.526389, -114.529194, -114.52775, -114.532222, -114.537083, 
    -114.5475, -114.545222, -114.552722, -114.568111, -114.582972, -114.585, 
    -114.580889, -114.581806, -114.592083, -114.598556, -114.601861, 
    -114.59925, -114.605, -114.602389, -114.604806, -114.608278, -114.605556, 
    -114.611444, -114.619806, -114.623222, -114.631444, -114.638389, 
    -114.653667, -114.667278, -114.674861, -114.697583, -114.700111, 
    -114.703583, -114.711583, -114.717611, -114.71825, -114.724083, 
    -114.728444, -114.734667, -114.737333, -114.73575, -114.739972, 
    -114.745611, -114.750972, -114.755861, -114.768917, -114.778111, 
    -114.785806, -114.797417, -114.809917, -114.824028, -114.830722, 
    -114.836556, -114.845028, -114.850861, -114.861444, -114.86225, 
    -114.873944, -114.879778, -114.886694, -114.900306, -114.90325, 
    -114.912556, -114.949778, -114.965472, -114.979972, -114.992278, 
    -115.014111, -115.028556, -115.054306, -115.07125, -115.096222, 
    -115.102778, -115.13075, -115.139639, -115.15525, -115.168639, 
    -115.179583, -115.189167, -115.196167, -115.213556, -115.218222, 
    -115.222333, -115.22875, -115.235556, -115.247778, -115.279528, 
    -115.29725, -115.314306, -115.341306, -115.367056, -115.378611, 
    -115.385028, -115.390111, -115.407167, -115.415111, -115.453306, 
    -115.463083, -115.477861, -115.493028, -115.504583, -115.514111, 
    -115.523333, -115.54025, -115.5525, -115.564167, -115.572806, -115.58475, 
    -115.602917, -115.621139, -115.678972, -115.696222, -115.699972, 
    -115.687556, -115.685833, -115.702583, -115.723389, -115.744056, 
    -115.787472, -115.803278, -115.8115, -115.81425, -115.79875, -115.781389, 
    -115.790667, -115.788583, -115.801444, -115.803056, -115.794806, 
    -115.795611, -115.803, -115.810833, -115.816528, -115.824694, 
    -115.834972, -115.845083, -115.863833, -115.900972, -115.919056, 
    -115.935861, -115.95475, -115.9815, -115.986694, -115.971167, 
    -115.968028, -115.964361, -115.950889, -115.940278, -115.943444, 
    -115.935861, -115.929667, -115.937972, -115.945472, -115.951194, 
    -115.967889, -115.97775, -115.982722, -115.97775, -115.993806, 
    -115.993222, -115.998222, -115.998194, -115.987194, -115.979056, 
    -115.973056, -115.976639, -115.967778, -115.961833, -115.962389, 
    -115.955889, -115.959222, -115.956417, -115.965639, -115.969028, 
    -115.979472, -115.993222, -115.996083, -116.005056, -116.015806, 
    -116.020833, -116.025417, -116.014639, -116.014583, -116.010417, 
    -115.994222, -115.995917, -115.99225, -115.9905, -115.991444, 
    -115.986944, -115.985389, -115.978917, -115.986222, -116, -116.006278, 
    -116.008, -116.004583, -116.004667, -116.01375, -116.02, -116.030444, 
    -116.034583, -116.043778, -116.047944, -116.048778, -116.044611, 
    -116.032111, -116.027139, -116.032917, -116.047111, -116.049639, 
    -116.060417, -116.078389, -116.086722, -116.096722, -116.105833, 
    -116.148333, -116.156667, -116.165861, -116.175889, -116.189167, 
    -116.205417, -116.214583, -116.222528, -116.235833, -116.245, 
    -116.268389, -116.284194, -116.295833, -116.32, -116.3275, -116.335444, 
    -116.340389, -116.31475, -116.310528, -116.33625, -116.341667, 
    -116.354083, -116.354028, -116.361111, -116.372111, -116.373139, 
    -116.388028, -116.396028, -116.403306, -116.408611, -116.416472, -116.42, 
    -116.432917, -116.441444, -116.449, -116.451889, -116.459694, 
    -116.457194, -116.458806, -116.471528, -116.473222, -116.480667, 
    -116.490306, -116.489278, -116.504889, -116.503722, -116.514111, 
    -116.525972, -116.547444, -116.553639, -116.573833, -116.583056, 
    -116.599028, -116.606111, -116.611528, -116.632972, -116.637333, 
    -116.648222, -116.648611, -116.661417, -116.661944, -116.666222, 
    -116.668444, -116.678389, -116.684556, -116.693639, -116.690472, 
    -116.694139, -116.683083, -116.674472, -116.655806, -116.652528, 
    -116.655444, -116.666389, -116.669278, -116.653972, -116.652222, 
    -116.68025, -116.679111, -116.693361, -116.691333, -116.698611, 
    -116.70975, -116.716306, -116.719056, -116.717417, -116.726139, 
    -116.728306, -116.735833, -116.738361, -116.749, -116.743917, 
    -116.743083, -116.72825, -116.697667, -116.682944, -116.672194, 
    -116.663194, -116.652472, -116.640611, -116.627361, -116.622722, 
    -116.626306, -116.625861, -116.632389, -116.640806, -116.659, -116.639, 
    -116.635472, -116.631444, -116.632944, -116.63875, -116.63975, 
    -116.623194, -116.620667, -116.614139, -116.611583, -116.622333, 
    -116.611444, -116.614778, -116.622861, -116.6215, -116.629, -116.631639, 
    -116.629917, -116.640611, -116.663306, -116.668667, -116.703194, 
    -116.714667, -116.720694, -116.750861, -116.757278, -116.762333, 
    -116.778278, -116.791389, -116.798972, -116.833917, -116.860583, 
    -116.866222, -116.882389, -116.888306, -116.884, -116.888306, 
    -116.889194, -116.903556, -116.909417, -116.915111, -116.922556, 
    -116.934694, -116.948472, -116.974444, -117.006083, -117.011806, 
    -117.024833, -117.038444, -117.054667, -117.066, -117.076778, 
    -117.090139, -117.1025, -117.111694, -117.120833, -117.125056, 
    -117.124167, -117.134917, -117.132528, -117.138306, -117.161722, 
    -117.180861, -117.196528, -117.206472, -117.223417, -117.228361, 
    -117.229139, -117.223528, -117.209444, -117.191778, -117.186944, 
    -117.188361, -117.16375, -117.167444, -117.164111, -117.157917, 
    -117.154167, -117.160056, -117.145056, -117.1375, -117.130944, 
    -117.130778, -117.126861, -117.129361, -117.121778, -117.114111, 
    -117.098222, -117.100889, -117.116139, -117.120694, -117.124972, 
    -117.120083, -117.134139, -117.140611, -117.139417, -117.174139, 
    -117.175861, -117.178778, -117.206917, -117.216528, -117.225806, 
    -117.225056, -117.220111, -117.221389, -117.236722, -117.240222, 
    -117.238694, -117.233444, -117.236944, -117.23725, -117.240139, -117.247, 
    -117.246472, -117.256833, -117.259417, -117.257111, -117.249222, 
    -117.253778, -117.254222, -117.259444, -117.281778, -117.28325, 
    -117.283444, -117.280139, -117.272, -117.265278, -117.259333, 
    -117.252472, -117.255111, -117.260389, -117.260611, -117.27, -117.281778, 
    -117.298833, -117.332444, -117.337278, -117.362278, -117.399778, 
    -117.405861, -117.435028, -117.507889, -117.551889, -117.579083, 
    -117.599389, -117.606111, -117.616583, -117.6555, -117.687444, 
    -117.69975, -117.707889, -117.710194, -117.717167, -117.728444, 
    -117.737944, -117.742361, -117.753556, -117.761778, -117.786528, 
    -117.806667, -117.809722, -117.820889, -117.823556, -117.834, 
    -117.842583, -117.860583, -117.87425, -117.9285, -117.941028, -117.9905, 
    -118.032528, -118.062556, -118.090861, -118.094611, -118.087528, 
    -118.08925, -118.096667, -118.097528, -118.101694, -118.105028, 
    -118.115861, -118.116667, -118.132472, -118.163333, -118.181722, 
    -118.186667, -118.190861, -118.191639, -118.1975, -118.206722, -118.2025, 
    -118.187139, -118.189639, -118.185833, -118.205028, -118.20425, 
    -118.194611, -118.199167, -118.200861, -118.207111, -118.2075, 
    -118.212111, -118.206694, -118.214167, -118.215417, -118.208778, 
    -118.208806, -118.210889, -118.214194, -118.215028, -118.221667, 
    -118.227556, -118.243722, -118.241722, -118.230056, -118.222556, 
    -118.222583, -118.230833, -118.239222, -118.244611, -118.2475, 
    -118.253778, -118.2625, -118.265444, -118.267528, -118.26875, 
    -118.264583, -118.268333, -118.276278, -118.269194, -118.248417, 
    -118.230028, -118.224194, -118.221667, -118.212972, -118.220833, 
    -118.222528, -118.249222, -118.254194, -118.259194, -118.263361, 
    -118.261278, -118.2675, -118.269972, -118.270861, -118.275417, 
    -118.273333, -118.277917, -118.278389, -118.287944, -118.280028, 
    -118.272972, -118.277139, -118.278778, -118.270444, -118.274611, 
    -118.272944, -118.275889, -118.282556, -118.281306, -118.285417, 
    -118.281306, -118.289194, -118.295833, -118.300861, -118.320028, 
    -118.324194, -118.352556, -118.356722, -118.364194, -118.375917, 
    -118.380861, -118.3875, -118.400028, -118.405861, -118.413333, 
    -118.416278, -118.429583, -118.425889, -118.410472, -118.407528, 
    -118.395472, -118.392917, -118.400444, -118.412917, -118.457083, 
    -118.4475, -118.442917, -118.446222, -118.445833, -118.454194, 
    -118.449611, -118.452944, -118.448778, -118.452139, -118.448778, 
    -118.452944, -118.449222, -118.44875, -118.458361, -118.477083, 
    -118.478778, -118.48625, -118.486778, -118.494333, -118.499278, 
    -118.501361, -118.523722, -118.534556, -118.545417, -118.573611, 
    -118.586, -118.600889, -118.611556, -118.673167, -118.683139, 
    -118.699583, -118.709833, -118.74275, -118.757306, -118.786417, 
    -118.794278, -118.803861, -118.807917, -118.851333, -118.877778, 
    -118.918139, -118.927278, -118.940472, -118.956389, -118.98, -119.002806, 
    -119.009944, -119.038194, -119.063639, -119.090056, -119.098972, 
    -119.109306, -119.133111, -119.195611, -119.215778, -119.223028, 
    -119.23575, -119.264861, -119.270694, -119.267306, -119.264972, 
    -119.259694, -119.267806, -119.272167, -119.276361, -119.28875, 
    -119.305139, -119.318389, -119.322389, -119.341, -119.350111, 
    -119.372667, -119.392333, -119.431417, -119.444528, -119.458972, 
    -119.472278, -119.4795, -119.490361, -119.516, -119.528333, -119.538472, 
    -119.565861, -119.579917, -119.597667, -119.615278, -119.6355, 
    -119.673417, -119.687889, -119.692778, -119.692278, -119.699417, 
    -119.704972, -119.713833, -119.728, -119.744333, -119.796278, 
    -119.838278, -119.845361, -119.863889, -119.880972, -119.88925, -119.921, 
    -119.929722, -119.957944, -119.980861, -119.990861, -120.005972, 
    -120.016833, -120.023472, -120.034, -120.06075, -120.069222, -120.07925, 
    -120.09325, -120.117361, -120.140889, -120.172444, -120.218806, 
    -120.277056, -120.297, -120.304472, -120.334389, -120.337528, 
    -120.409389, -120.418139, -120.421, -120.444722, -120.455167, 
    -120.464361, -120.473222, -120.477389, -120.481222, -120.492472, 
    -120.492917, -120.498056, -120.503444, -120.512167, -120.541528, 
    -120.555194, -120.567944, -120.581694, -120.60175, -120.617722, 
    -120.624611, -120.633667, -120.638694, -120.642028, -120.641389, 
    -120.652528, -120.646861, -120.647806, -120.642528, -120.645056, 
    -120.638111, -120.620139, -120.606722, -120.599222, -120.604472, 
    -120.602472, -120.608611, -120.61675, -120.629389, -120.632583, -120.631, 
    -120.639583, -120.620028, -120.611861, -120.613139, -120.641972, 
    -120.640861, -120.648361, -120.672694, -120.674222, -120.664917, 
    -120.669111, -120.661833, -120.645972, -120.632361, -120.631472, 
    -120.641444, -120.647333, -120.657972, -120.672861, -120.684611, 
    -120.705972, -120.726, -120.735694, -120.749111, -120.756389, 
    -120.754222, -120.769556, -120.779917, -120.786972, -120.814556, 
    -120.859222, -120.863222, -120.862028, -120.869972, -120.879917, 
    -120.887361, -120.899806, -120.8975, -120.900889, -120.8965, -120.896444, 
    -120.891694, -120.891611, -120.881694, -120.872583, -120.864167, 
    -120.863361, -120.859194, -120.858028, -120.860889, -120.867333, 
    -120.86175, -120.844889, -120.844806, -120.835222, -120.828056, 
    -120.833639, -120.835861, -120.843417, -120.857889, -120.863111, 
    -120.868389, -120.871611, -120.871833, -120.865361, -120.863278, 
    -120.866639, -120.885806, -120.907, -120.949833, -120.954056, 
    -120.969806, -121.005556, -121.025694, -121.039528, -121.048361, 
    -121.06125, -121.105139, -121.106944, -121.115139, -121.123306, 
    -121.125917, -121.133, -121.144944, -121.168833, -121.190694, 
    -121.194389, -121.192972, -121.19575, -121.220111, -121.242639, 
    -121.249917, -121.261361, -121.27225, -121.280583, -121.285194, 
    -121.293167, -121.318472, -121.314389, -121.319444, -121.317111, 
    -121.320556, -121.316028, -121.317944, -121.328028, -121.326083, 
    -121.333222, -121.358083, -121.372667, -121.375778, -121.387806, 
    -121.414556, -121.426111, -121.447194, -121.465278, -121.462556, 
    -121.476417, -121.469583, -121.470222, -121.478667, -121.476, 
    -121.484556, -121.487972, -121.505222, -121.535889, -121.552972, 
    -121.567306, -121.573667, -121.58425, -121.593833, -121.590861, 
    -121.594278, -121.607056, -121.621861, -121.625278, -121.63525, 
    -121.646306, -121.676944, -121.699472, -121.718417, -121.748361, 
    -121.754417, -121.77975, -121.787028, -121.797167, -121.806056, 
    -121.814444, -121.816917, -121.835611, -121.839583, -121.851694, 
    -121.861917, -121.875667, -121.887611, -121.903056, -121.904333, 
    -121.900111, -121.897056, -121.893472, -121.907556, -121.903667, 
    -121.907889, -121.903667, -121.904444, -121.907083, -121.915194, 
    -121.91875, -121.916083, -121.930222, -121.927889, -121.936583, 
    -121.942667, -121.946639, -121.938722, -121.941139, -121.956028, 
    -121.955056, -121.939556, -121.937861, -121.927194, -121.929361, 
    -121.934389, -121.930917, -121.935861, -121.941722, -121.942806, 
    -121.949306, -121.952889, -121.972056, -121.980361, -121.973528, 
    -121.967806, -121.96125, -121.957083, -121.949306, -121.943528, 
    -121.939417, -121.939556, -121.935333, -121.924444, -121.912889, 
    -121.902528, -121.888056, -121.874583, -121.859972, -121.831583, 
    -121.816139, -121.80875, -121.808028, -121.803583, -121.805444, 
    -121.790278, -121.809778, -121.814806, -121.863556, -121.89775, 
    -121.930278, -121.940417, -121.953806, -121.972556, -122.013472, 
    -122.025139, -122.026833, -122.04075, -122.051194, -122.058944, 
    -122.068306, -122.075944, -122.078111, -122.103583, -122.123194, 
    -122.136, -122.141444, -122.153583, -122.163583, -122.168444, 
    -122.171611, -122.186722, -122.195056, -122.207583, -122.218361, 
    -122.225861, -122.234583, -122.255472, -122.28, -122.294222, -122.313333, 
    -122.321694, -122.333361, -122.334639, -122.340472, -122.340472, 
    -122.347556, -122.364639, -122.362139, -122.367972, -122.385056, 
    -122.396667, -122.400444, -122.407111, -122.409583, -122.412111, 
    -122.418833, -122.422083, -122.420028, -122.4155, -122.41125, 
    -122.412917, -122.403, -122.400417, -122.407917, -122.409667, 
    -122.423778, -122.427917, -122.444583, -122.445444, -122.456278, 
    -122.478389, -122.491722, -122.49625, -122.496722, -122.502528, 
    -122.501278, -122.507167, -122.518778, -122.52125, -122.515472, 
    -122.515444, -122.519639, -122.518, -122.522111, -122.515917, 
    -122.507556, -122.500472, -122.502944, -122.497972, -122.499611, 
    -122.495444, -122.494639, -122.499667, -122.509583, -122.515472, 
    -122.5075, -122.488389, -122.478389, -122.455028, -122.436722, 
    -122.423389, -122.415889, -122.403361, -122.387111, -122.387083, 
    -122.381278, -122.385417, -122.384639, -122.380472, -122.382944, 
    -122.374611, -122.375861, -122.384667, -122.375861, -122.369583, 
    -122.375444, -122.373389, -122.365028, -122.356278, -122.361306, 
    -122.35875, -122.364167, -122.374167, -122.37675, -122.382556, 
    -122.377139, -122.378778, -122.375472, -122.392139, -122.386306, 
    -122.3805, -122.380389, -122.389222, -122.393778, -122.378389, 
    -122.373778, -122.378778, -122.375528, -122.377139, -122.390056, 
    -122.392083, -122.381278, -122.389222, -122.388361, -122.363778, 
    -122.368028, -122.35625, -122.357972, -122.372583, -122.377917, 
    -122.362528, -122.35425, -122.335917, -122.333444, -122.321722, 
    -122.315889, -122.314639, -122.306694, -122.296694, -122.295, 
    -122.286722, -122.275028, -122.261694, -122.256694, -122.247917, 
    -122.248361, -122.233361, -122.227972, -122.226306, -122.237528, 
    -122.220889, -122.218806, -122.2275, -122.206722, -122.196306, 
    -122.197944, -122.212889, -122.215861, -122.211306, -122.20375, 
    -122.204639, -122.200028, -122.187583, -122.182528, -122.177972, 
    -122.167972, -122.166667, -122.157556, -122.158389, -122.144222, 
    -122.136694, -122.130472, -122.1205, -122.113361, -122.101722, 
    -122.102944, -122.096667, -122.092528, -122.082583, -122.078361, 
    -122.075889, -122.0675, -122.065028, -122.043361, -122.031778, 
    -122.040472, -122.035861, -122.02675, -122.021722, -122.022556, 
    -122.008944, -122.027472, -122.040056, -122.050861, -122.057944, 
    -122.047556, -122.054194, -122.059222, -122.071722, -122.083389, 
    -122.085833, -122.096694, -122.108806, -122.112917, -122.111306, 
    -122.121333, -122.131306, -122.130417, -122.135417, -122.149583, 
    -122.148028, -122.1505, -122.155417, -122.152083, -122.155528, 
    -122.154611, -122.158778, -122.156306, -122.16375, -122.192917, 
    -122.190889, -122.185917, -122.189167, -122.194667, -122.189556, 
    -122.190444, -122.198389, -122.202972, -122.200889, -122.208389, 
    -122.214194, -122.243333, -122.243361, -122.239611, -122.262111, 
    -122.252528, -122.239222, -122.240083, -122.274278, -122.2775, 
    -122.280917, -122.282528, -122.286333, -122.283389, -122.289222, 
    -122.289194, -122.294222, -122.300444, -122.299167, -122.307528, 
    -122.308389, -122.315889, -122.317583, -122.332111, -122.334639, 
    -122.330833, -122.322556, -122.322083, -122.327556, -122.337528, 
    -122.342917, -122.337528, -122.322528, -122.312083, -122.330028, 
    -122.331278, -122.297944, -122.29925, -122.313778, -122.313333, 
    -122.299639, -122.30625, -122.310083, -122.315889, -122.317917, 
    -122.313361, -122.313778, -122.318361, -122.322139, -122.317583, 
    -122.314167, -122.30875, -122.317917, -122.325417, -122.31425, 
    -122.314639, -122.316694, -122.322556, -122.324694, -122.322139, 
    -122.329222, -122.351694, -122.346306, -122.3525, -122.355028, -122.36, 
    -122.363833, -122.370833, -122.375472, -122.367944, -122.363444, 
    -122.368417, -122.381722, -122.395861, -122.387139, -122.398333, 
    -122.414194, -122.414611, -122.422972, -122.421306, -122.429194, 
    -122.412583, -122.410028, -122.398361, -122.39625, -122.399194, 
    -122.393778, -122.400889, -122.389167, -122.383417, -122.371722, 
    -122.367167, -122.359611, -122.366306, -122.366694, -122.337472, 
    -122.33175, -122.316278, -122.299333, -122.291167, -122.290361, 
    -122.282722, -122.273806, -122.267167, -122.264833, -122.256389, 
    -122.256972, -122.274972, -122.2765, -122.298583, -122.322694, 
    -122.349833, -122.358972, -122.37475, -122.399583, -122.409083, 
    -122.406611, -122.411028, -122.446528, -122.454889, -122.456028, 
    -122.46025, -122.500056, -122.510864, -122.51575, -122.508556, 
    -122.491556, -122.491556, -122.488139, -122.485778, -122.486444, 
    -122.499056, -122.496667, -122.499889, -122.488139, -122.478028, 
    -122.462472, -122.448, -122.456694, -122.466722, -122.472528, 
    -122.476694, -122.481722, -122.479583, -122.482583, -122.502139, 
    -122.489611, -122.486278, -122.479194, -122.479167, -122.489167, 
    -122.505028, -122.512917, -122.505861, -122.502167, -122.492556, 
    -122.485083, -122.475444, -122.472139, -122.476306, -122.475028, 
    -122.460861, -122.449167, -122.438778, -122.452556, -122.463, 
    -122.458361, -122.472944, -122.475028, -122.489222, -122.503778, 
    -122.499611, -122.497528, -122.510917, -122.51175, -122.517528, 
    -122.519222, -122.523361, -122.519639, -122.522556, -122.513361, 
    -122.508361, -122.497972, -122.496722, -122.478806, -122.479639, 
    -122.472083, -122.472139, -122.477556, -122.4825, -122.491694, 
    -122.504194, -122.510028, -122.522556, -122.529611, -122.528389, 
    -122.537944, -122.537111, -122.540833, -122.551722, -122.554583, 
    -122.560028, -122.565889, -122.572528, -122.577556, -122.587528, 
    -122.604167, -122.620889, -122.630083, -122.65175, -122.666667, 
    -122.684222, -122.703333, -122.728333, -122.740028, -122.754167, 
    -122.766694, -122.774222, -122.778361, -122.780861, -122.785056, 
    -122.792083, -122.804194, -122.815028, -122.834083, -122.859972, 
    -122.899361, -122.930694, -122.933306, -122.937556, -122.94175, 
    -122.953028, -122.965722, -122.979889, -122.983806, -122.967528, 
    -122.965861, -122.991694, -123, -123.023028, -123.024278, -123.014528, 
    -123.010028, -122.983194, -122.956806, -122.95175, -122.956889, 
    -122.969972, -122.967528, -122.969417, -122.983194, -122.983194, 
    -122.996667, -122.995889, -122.989833, -122.9825, -122.974917, 
    -122.969889, -122.979889, -122.988306, -123.001778, -123.026917, 
    -123.046806, -123.054083, -123.052806, -123.062361, -123.066722, 
    -123.072028, -123.080806, -123.075944, -123.069833, -123.072528, 
    -123.088028, -123.100833, -123.103111, -123.122917, -123.132639, 
    -123.145472, -123.154917, -123.155444, -123.163889, -123.168139, 
    -123.202417, -123.230667, -123.237972, -123.246806, -123.25525, 
    -123.273972, -123.278444, -123.286333, -123.305361, -123.306639, 
    -123.323722, -123.33075, -123.335333, -123.3425, -123.3395, -123.345222, 
    -123.352111, -123.360444, -123.371194, -123.373389, -123.369333, 
    -123.369556, -123.376222, -123.390139, -123.390444, -123.39675, 
    -123.39525, -123.401889, -123.399722, -123.404389, -123.410417, 
    -123.408472, -123.420222, -123.434, -123.436639, -123.434222, 
    -123.447694, -123.453861, -123.461611, -123.485472, -123.49525, 
    -123.515222, -123.528472, -123.529167, -123.535111, -123.535806, 
    -123.546167, -123.563333, -123.56425, -123.579056, -123.588389, 
    -123.599306, -123.604583, -123.605944, -123.602417, -123.605028, 
    -123.614139, -123.627833, -123.641694, -123.648056, -123.657528, 
    -123.665972, -123.681694, -123.689361, -123.703556, -123.71425, 
    -123.714083, -123.727389, -123.731667, -123.730083, -123.744278, 
    -123.730667, -123.702639, -123.697472, -123.69075, -123.695083, 
    -123.695639, -123.692306, -123.695556, -123.707583, -123.709056, 
    -123.715028, -123.714944, -123.720972, -123.721056, -123.729944, 
    -123.734972, -123.739083, -123.735583, -123.75275, -123.757556, 
    -123.766028, -123.771028, -123.773972, -123.770694, -123.776583, 
    -123.770861, -123.778222, -123.771778, -123.780694, -123.775972, 
    -123.787278, -123.785028, -123.792583, -123.799639, -123.805194, 
    -123.804056, -123.797472, -123.798389, -123.795417, -123.80175, 
    -123.805667, -123.812361, -123.809611, -123.802639, -123.801806, 
    -123.809139, -123.807139, -123.813417, -123.819833, -123.818083, 
    -123.829194, -123.823694, -123.826333, -123.817583, -123.827556, 
    -123.819278, -123.824167, -123.820667, -123.823222, -123.813417, 
    -123.821083, -123.810083, -123.818889, -123.822611, -123.815972, 
    -123.816611, -123.805833, -123.804083, -123.807472, -123.798972, 
    -123.789028, -123.768, -123.772333, -123.778556, -123.779056, 
    -123.787333, -123.790972, -123.784778, -123.783972, -123.788722, 
    -123.787333, -123.789111, -123.795083, -123.796639, -123.809861, 
    -123.833278, -123.831889, -123.838222, -123.834917, -123.839889, 
    -123.840806, -123.847139, -123.852472, -123.886056, -123.906861, 
    -123.930556, -123.940556, -123.956444, -123.98025, -123.991694, 
    -124.006806, -124.01475, -124.019472, -124.038972, -124.060083, 
    -124.070361, -124.075639, -124.081833, -124.080806, -124.088472, 
    -124.110972, -124.140611, -124.173944, -124.189028, -124.214167, 
    -124.236667, -124.259889, -124.278306, -124.291611, -124.325944, 
    -124.330333, -124.35325, -124.364917, -124.365, -124.349944, -124.351528, 
    -124.363139, -124.366583, -124.366556, -124.3715, -124.383028, -124.395, 
    -124.4125, -124.410417, -124.394944, -124.3865, -124.385722, -124.390917, 
    -124.375, -124.365139, -124.325556, -124.322389, -124.308528, 
    -124.309639, -124.318583, -124.319972, -124.272556, -124.235667, 
    -124.225611, -124.227472, -124.223528, -124.210444, -124.201861, 
    -124.199389, -124.205889, -124.2035, -124.198694, -124.189444, 
    -124.180889, -124.18075, -124.186472, -124.200194, -124.218361, 
    -124.222861, -124.228, -124.234833, -124.218056, -124.167972, 
    -124.138167, -124.11725, -124.113056, -124.124861, -124.139694, 
    -124.145889, -124.146722, -124.15375, -124.15075, -124.160111, 
    -124.156528, -124.159556, -124.156, -124.165056, -124.160806, 
    -124.159861, -124.164972, -124.164278, -124.158167, -124.149722, 
    -124.143806, -124.106889, -124.1065, -124.110861, -124.10625, 
    -124.098444, -124.085139, -124.086778, -124.069139, -124.064028, 
    -124.068194, -124.083361, -124.074722, -124.092861, -124.101306, 
    -124.097139, -124.104083, -124.100778, -124.115778, -124.120944, 
    -124.135611, -124.140944, -124.137667, -124.142528, -124.142611, 
    -124.149306, -124.165889, -124.181639, -124.184917, -124.194278, 
    -124.197528, -124.195361, -124.198306, -124.21625, -124.243028, 
    -124.255778, -124.250833, -124.255861, -124.240861, -124.228389, 
    -124.207361, -124.204028, -124.209833, -124.205028, -124.209917, 
    -124.221667, -124.232972, -124.238778, -124.255, -124.270778, 
    -124.282167, -124.287806, -124.29175, -124.291056, -124.299778, 
    -124.308417, -124.320778, -124.32725, -124.338472, -124.344972, 
    -124.349444, -124.354861, -124.353333, -124.359194, -124.355111, 
    -124.353944, -124.357333, -124.362444, -124.368722, -124.362361, 
    -124.366, -124.362528, -124.367333, -124.372278, -124.377778, 
    -124.375611, -124.379889, -124.381333, -124.414, -124.409778, 
    -124.422639, -124.430139, -124.434389, -124.429194, -124.425889, 
    -124.426639, -124.431639, -124.4155, -124.416278, -124.422694, 
    -124.433917, -124.437556, -124.422083, -124.427583, -124.423389, 
    -124.423028, -124.426889, -124.421083, -124.424056, -124.406694, 
    -124.391222, -124.391444, -124.398028, -124.395389, -124.399889, 
    -124.404528, -124.410083, -124.404056, -124.40275, -124.408167, 
    -124.407167, -124.4155, -124.4135, -124.416667, -124.412333, -124.417917, 
    -124.452556, -124.449111, -124.455194, -124.475694, -124.492028, 
    -124.504694, -124.510028, -124.515389, -124.5255, -124.534778, 
    -124.553222, -124.565972, -124.568444, -124.565889, -124.55775, 
    -124.550722, -124.534639, -124.535861, -124.523833, -124.496639, -124.45, 
    -124.436694, -124.431583, -124.436722, -124.42425, -124.401667, 
    -124.394861, -124.395944, -124.382639, -124.388361, -124.388444, 
    -124.396167, -124.399806, -124.402611, -124.388056, -124.386889, 
    -124.375278, -124.375389, -124.368861, -124.362528, -124.356417, 
    -124.346972, -124.327083, -124.319889, -124.322722, -124.320056, 
    -124.313167, -124.306639, -124.302111, -124.296611, -124.285083, 
    -124.27875, -124.258056, -124.258056, -124.241167, -124.227861, 
    -124.216639, -124.217333, -124.207667, -124.189806, -124.175333, 
    -124.179667, -124.186861, -124.187944, -124.198639, -124.195861, 
    -124.200083, -124.198389, -124.190028, -124.20025, -124.208361, 
    -124.219111, -124.221861, -124.213556, -124.202167, -124.198389, 
    -124.192194, -124.198, -124.204889, -124.222139, -124.229167, -124.23475, 
    -124.239944, -124.246444, -124.251389, -124.265556, -124.272167, 
    -124.280611, -124.283944, -124.308222, -124.319139, -124.332917, 
    -124.339083, -124.301806, -124.2635, -124.230833, -124.206722, 
    -124.195667, -124.186694, -124.188778, -124.194667, -124.206028, 
    -124.192667, -124.166528, -124.141694, -124.135806, -124.130083, 
    -124.126361, -124.138, -124.123833, -124.123778, -124.128778, 
    -124.123806, -124.129611, -124.122111, -124.117111, -124.115472, 
    -124.111278, -124.115472, -124.108806, -124.115472, -124.110444, 
    -124.113833, -124.108806, -124.102889, -124.10875, -124.109583, 
    -124.094583, -124.084667, -124.072528, -124.060083, -124.056278, 
    -124.058389, -124.053417, -124.042556, -124.04, -124.030861, -124.026278, 
    -124.027472, -124.035861, -124.048361, -124.073389, -124.077556, 
    -124.082972, -124.081278, -124.085472, -124.077167, -124.067972, 
    -124.06875, -124.050861, -124.048389, -124.041278, -124.045472, 
    -124.040889, -124.025889, -124.018, -124.013444, -124.003778, 
    -124.009167, -124.023417, -124.023833, -124.0275, -124.046694, 
    -124.065028, -124.057944, -124.060861, -124.073389, -124.081278, 
    -124.079194, -124.072556, -124.06875, -124.057944, -124.05875, -124.0655, 
    -124.067972, -124.075417, -124.073778, -124.06875, -124.072917, 
    -124.073778, -124.06375, -124.063806, -124.068806, -124.065417, 
    -124.069611, -124.067583, -124.060472, -124.049639, -124.025056, 
    -124.028361, -124.017111, -124.012972, -124.018778, -124.016306, 
    -124.027139, -124.0255, -124.010028, -124.012611, -124.005194, 
    -124.004611, -124.016, -124.017778, -124.01425, -124.016, -124.009361, 
    -124.011667, -124.008556, -123.989917, -123.975944, -123.969528, 
    -123.972389, -123.971389, -123.974139, -123.981028, -123.97275, 
    -123.965083, -123.956667, -123.957583, -123.962694, -123.962389, 
    -123.971056, -123.97725, -124.00825, -124.008806, -123.999139, 
    -123.994028, -123.992944, -123.981139, -123.973833, -123.959667, 
    -123.952361, -123.961056, -123.962222, -123.958583, -123.952444, 
    -123.938333, -123.932528, -123.940056, -123.961694, -123.974139, 
    -123.970778, -123.975917, -123.963472, -123.956917, -123.956056, 
    -123.944667, -123.937861, -123.916306, -123.889917, -123.893167, 
    -123.881861, -123.878833, -123.869111, -123.865167, -123.869639, 
    -123.883944, -123.88325, -123.890306, -123.888472, -123.898417, 
    -123.898194, -123.908472, -123.896333, -123.90275, -123.905528, 
    -123.913583, -123.914722, -123.918139, -123.934139, -123.943778, 
    -123.958528, -123.942417, -123.941222, -123.93275, -123.926028, 
    -123.925278, -123.922083, -123.904528, -123.906, -123.901, -123.904167, 
    -123.893806, -123.893778, -123.916278, -123.920694, -123.930861, 
    -123.934528, -123.929972, -123.937333, -123.940111, -123.939056, 
    -123.945056, -123.96525, -123.969611, -123.979778, -123.984389, 
    -123.969889, -123.970278, -123.96425, -123.962417, -123.965194, 
    -123.969972, -123.966639, -123.968361, -123.971667, -123.978194, 
    -123.980028, -123.993472, -123.993556, -123.976389, -123.96875, 
    -123.940111, -123.92875, -123.91875, -123.927889, -123.933778, 
    -123.947944, -123.99625, -124.013139, -124.021722, -124.023361, 
    -124.019167, -124.011417, -123.994194, -123.990417, -123.995889, 
    -124.002139, -123.988389, -123.968361, -123.95175, -123.950028, 
    -123.909167, -123.901694, -123.878306, -123.865889, -123.862528, 
    -123.838389, -123.829194, -123.824167, -123.820444, -123.816639, 
    -123.808833, -123.813417, -123.825861, -123.844194, -123.860861, 
    -123.868333, -123.845889, -123.820861, -123.797556, -123.795833, 
    -123.779222, -123.770417, -123.768389, -123.758417, -123.76375, 
    -123.760444, -123.753333, -123.726694, -123.719667, -123.726722, 
    -123.724222, -123.717528, -123.7175, -123.689194, -123.6775, -123.628306, 
    -123.625056, -123.636278, -123.630806, -123.614222, -123.622583, 
    -123.605056, -123.595889, -123.589639, -123.587139, -123.577889, 
    -123.585528, -123.564167, -123.545861, -123.542139, -123.550444, 
    -123.542528, -123.493389, -123.482056, -123.470833, -123.441667, 
    -123.43375, -123.431306, -123.438333, -123.456694, -123.480028, 
    -123.498361, -123.518417, -123.530056, -123.5325, -123.561722, 
    -123.565056, -123.574222, -123.583361, -123.620889, -123.632556, 
    -123.6725, -123.681278, -123.678806, -123.681278, -123.687944, 
    -123.685472, -123.7025, -123.706722, -123.717111, -123.712917, 
    -123.718361, -123.725444, -123.729167, -123.749167, -123.765, 
    -123.776694, -123.786722, -123.804194, -123.819167, -123.836694, 
    -123.840806, -123.850833, -123.85125, -123.859222, -123.8675, 
    -123.870889, -123.875833, -123.909972, -123.923361, -123.929194, 
    -123.944167, -123.969667, -123.970056, -123.993389, -124.022861, 
    -124.030472, -124.039806, -124.048083, -124.051028, -124.034694, 
    -124.031611, -124.037194, -124.040444, -124.043778, -124.051444, 
    -124.056917, -124.082444, -124.088306, -124.084667, -124.072167, 
    -124.078028, -124.077722, -124.065806, -124.058528, -124.05675, 
    -124.066833, -124.059306, -124.046694, -124.028278, -124.030611, 
    -124.033694, -124.047083, -124.047167, -124.050944, -124.0375, 
    -124.02675, -124.023139, -124.024111, -124.028611, -124.029944, 
    -124.025139, -124.017333, -124.01475, -124.018694, -124.014861, 
    -124.008944, -123.999194, -123.995833, -123.980028, -123.980833, 
    -123.973389, -123.969194, -123.96125, -123.955028, -123.952556, 
    -123.949583, -123.952972, -123.952944, -123.940028, -123.93625, 
    -123.923806, -123.932083, -123.93125, -123.939639, -123.935083, 
    -123.923778, -123.926333, -123.921694, -123.895861, -123.8875, 
    -123.886306, -123.905833, -123.909639, -123.908778, -123.93, -123.937556, 
    -123.942972, -123.942972, -123.92625, -123.919556, -123.922556, 
    -123.9125, -123.897111, -123.898806, -123.892944, -123.898028, 
    -123.892944, -123.895861, -123.905917, -123.923, -123.920389, 
    -123.932083, -123.954583, -123.960528, -123.96125, -123.955028, 
    -123.944194, -123.930056, -123.916694, -123.915833, -123.932139, 
    -123.929194, -123.922889, -123.928361, -123.934222, -123.939583, 
    -123.937556, -123.92125, -123.920444, -123.9275, -123.921694, 
    -123.914194, -123.903389, -123.857583, -123.839194, -123.825083, 
    -123.819222, -123.81875, -123.831306, -123.825944, -123.830889, 
    -123.830444, -123.835, -123.840472, -123.8425, -123.846667, -123.848778, 
    -123.841639, -123.847528, -123.863389, -123.878389, -123.886694, -123.89, 
    -123.8875, -123.890861, -123.900889, -123.914278, -123.917972, 
    -123.91125, -123.925889, -123.947611, -123.975833, -123.974611, 
    -123.985472, -123.973833, -123.987972, -123.965806, -123.9675, 
    -123.972528, -123.984194, -124.000944, -124.017778, -124.028222, 
    -124.0355, -124.035861, -124.039806, -124.091972, -124.095194, 
    -124.095833, -124.104333, -124.124306, -124.138361, -124.125361, 
    -124.117944, -124.110861, -124.109806, -124.095139, -124.089111, 
    -124.095917, -124.101083, -124.0945, -124.084944, -124.084639, 
    -124.072417, -124.066056, -124.043944, -124.040361, -124.044528, 
    -124.054278, -124.063667, -124.053583, -124.050167, -124.042972, 
    -124.026917, -124.013389, -123.999583, -124.009944, -124.008639, 
    -124.003111, -124, -123.9825, -123.956667, -123.934222, -123.875833, 
    -123.850056, -123.822528, -123.80625, -123.811722, -123.834139, 
    -123.876694, -123.892528, -123.8975, -123.926722, -123.947528, 
    -123.950472, -123.945917, -123.916694, -123.915472, -123.925111, 
    -123.986667, -124.013278, -124.02125, -124.012194, -124.008278, 
    -124.019722, -124.019694, -124.028472, -124.046806, -124.052194, 
    -124.054472, -124.054139, -124.058139, -124.063333, -124.12075, 
    -124.145389, -124.151417, -124.145389, -124.135917, -124.13875, 
    -124.129083, -124.12775, -124.124528, -124.12675, -124.132472, 
    -124.159861, -124.161806, -124.150889, -124.157472, -124.173861, 
    -124.167278, -124.176917, -124.180528, -124.184611, -124.189722, 
    -124.206, -124.241472, -124.260111, -124.2725, -124.273333, -124.279528, 
    -124.300972, -124.285111, -124.310167, -124.321528, -124.326333, 
    -124.338083, -124.339389, -124.344361, -124.341278, -124.344667, 
    -124.341417, -124.343028, -124.348139, -124.343583, -124.347, 
    -124.357194, -124.350028, -124.358278, -124.389917, -124.413528, 
    -124.425333, -124.434806, -124.431861, -124.449806, -124.4555, 
    -124.480639, -124.481833, -124.474861, -124.493389, -124.497278, 
    -124.503472, -124.515861, -124.526, -124.542861, -124.5415, -124.554389, 
    -124.553, -124.561417, -124.562861, -124.573111, -124.581111, 
    -124.594806, -124.604333, -124.613139, -124.611222, -124.633278, 
    -124.63125, -124.641472, -124.635972, -124.643028, -124.649583, 
    -124.643333, -124.642, -124.653583, -124.66225, -124.668833, -124.66575, 
    -124.679, -124.673778, -124.672778, -124.682139, -124.678, -124.683, 
    -124.683, -124.698833, -124.697222, -124.688056, -124.693, -124.696333, 
    -124.712222, -124.708833, -124.718111, -124.723056, -124.7335, 
    -124.735583, -124.733444, -124.722667, -124.715167, -124.705194, 
    -124.699722, -124.691417, -124.707222, -124.699306, -124.683778, 
    -124.679583, -124.686278, -124.680472, -124.680833, -124.669222, 
    -124.664667, -124.66125, -124.664611, -124.657167, -124.658861, 
    -124.673861, -124.670028, -124.679194, -124.683389, -124.690889, 
    -124.697611, -124.70875, -124.707917, -124.713389, -124.727111, 
    -124.731278, -124.719222, -124.705056, -124.691722, -124.680056, 
    -124.675861, -124.667472, -124.65175, -124.63675, -124.637083, 
    -124.620028, -124.610056, -124.590083, -124.577556, -124.571722, 
    -124.564139, -124.539194, -124.52425, -124.512583, -124.490083, 
    -124.448333, -124.439167, -124.416694, -124.395083, -124.381778, 
    -124.358417, -124.339167, -124.300028, -124.302111, -124.297556, 
    -124.298361, -124.282472, -124.276667, -124.265056, -124.248389, 
    -124.219194, -124.180972, -124.14175, -124.128528, -124.11175, 
    -124.105972, -124.101389, -124.105944, -124.107583, -124.109278, 
    -124.072639, -124.049333, -124.023444, -124.020167, -124.000972, 
    -123.981806, -123.967639, -123.961778, -123.961, -123.945139, 
    -123.938444, -123.921861, -123.874278, -123.868472, -123.844222, 
    -123.829333, -123.819306, -123.810167, -123.778389, -123.757639, 
    -123.738444, -123.735139, -123.726778, -123.728417, -123.718417, 
    -123.707194, -123.709306, -123.704278, -123.70175, -123.671861, 
    -123.648444, -123.637194, -123.641, -123.626833, -123.589278, 
    -123.557611, -123.547639, -123.521778, -123.508417, -123.473444, 
    -123.445139, -123.404306, -123.401361, -123.40425, -123.428444, 
    -123.453417, -123.460556, -123.455889, -123.440194, -123.436, 
    -123.431833, -123.425944, -123.414278, -123.408472, -123.403528, 
    -123.37175, -123.345194, -123.33925, -123.323472, -123.310917, 
    -123.287583, -123.278444, -123.247611, -123.221833, -123.196778, 
    -123.181833, -123.154278, -123.103472, -123.105944, -123.134333, 
    -123.145083, -123.145472, -123.142611, -123.141833, -123.140139, 
    -123.156, -123.184694, -123.154306, -123.151, -123.149278, -123.131778, 
    -123.130083, -123.120917, -123.082667, -123.065111, -123.040528, 
    -123.045139, -123.047611, -123.053056, -123.049333, -123.046778, 
    -123.045472, -123.0405, -123.044694, -123.021861, -123.016833, -123.006, 
    -122.999278, -122.998889, -123.004694, -123.012194, -123.005556, 
    -123.007194, -123.0235, -123.021778, -123.041833, -123.040972, 
    -122.965972, -122.917611, -122.928056, -122.926361, -122.917583, 
    -122.874278, -122.858889, -122.862611, -122.887583, -122.886722, 
    -122.854194, -122.836806, -122.828028, -122.830972, -122.853472, 
    -122.860889, -122.880167, -122.893861, -122.881389, -122.886417, 
    -122.857583, -122.839278, -122.832667, -122.7885, -122.756806, 
    -122.763083, -122.751389, -122.765917, -122.780139, -122.798417, 
    -122.801417, -122.789278, -122.780139, -122.765556, -122.770556, 
    -122.764278, -122.755083, -122.750972, -122.735972, -122.727222, 
    -122.731806, -122.733, -122.728861, -122.731417, -122.71875, -122.719667, 
    -122.705028, -122.685028, -122.680444, -122.677111, -122.684611, 
    -122.681361, -122.684167, -122.686694, -122.697528, -122.699583, 
    -122.694222, -122.694194, -122.688361, -122.679194, -122.669167, 
    -122.658333, -122.652972, -122.65375, -122.645083, -122.638389, 
    -122.616722, -122.610472, -122.620889, -122.630083, -122.634639, 
    -122.648333, -122.668333, -122.692583, -122.692194, -122.681278, 
    -122.689639, -122.705028, -122.72175, -122.744194, -122.747972, 
    -122.7455, -122.749583, -122.7455, -122.75125, -122.749667, -122.757944, 
    -122.759583, -122.769167, -122.783778, -122.783861, -122.772111, 
    -122.778389, -122.8025, -122.812556, -122.832972, -122.827167, 
    -122.81375, -122.813778, -122.808778, -122.812111, -122.796306, 
    -122.788806, -122.791278, -122.787139, -122.796306, -122.793778, 
    -122.81425, -122.822139, -122.824639, -122.816306, -122.822139, 
    -122.840083, -122.852583, -122.854639, -122.846278, -122.850444, 
    -122.859194, -122.868778, -122.867944, -122.862972, -122.849611, 
    -122.852111, -122.858417, -122.864222, -122.873361, -122.872972, 
    -122.875861, -122.883806, -122.886306, -122.895472, -122.890444, 
    -122.908861, -122.902917, -122.903778, -122.920028, -122.929222, 
    -122.943361, -122.9575, -122.955889, -122.966722, -122.982611, 
    -122.986222, -122.981333, -122.988444, -123.007722, -123.01675, -123.033, 
    -123.040889, -123.0375, -123.050028, -123.056972, -123.101306, 
    -123.110444, -123.115222, -123.111833, -123.132722, -123.140778, 
    -123.148667, -123.157611, -123.155028, -123.158556, -123.142111, 
    -123.127222, -123.120722, -123.111861, -123.10625, -123.089639, 
    -123.073778, -123.07125, -123.048083, -123.045861, -123.052028, 
    -123.053278, -123.061861, -123.085833, -123.094333, -123.113333, 
    -123.121972, -123.083611, -123.073778, -123.055972, -123.070472, 
    -123.068583, -123.042056, -123.033556, -123.033389, -123.019278, 
    -122.996722, -122.984972, -122.975444, -122.976306, -122.971306, 
    -122.965083, -122.946722, -122.924167, -122.917972, -122.9205, 
    -122.916667, -122.90175, -122.878389, -122.870028, -122.85, -122.835861, 
    -122.827083, -122.838778, -122.838389, -122.805, -122.783417, -122.75175, 
    -122.747111, -122.749667, -122.739639, -122.731333, -122.714167, 
    -122.692139, -122.682611, -122.669222, -122.655028, -122.645, 
    -122.631722, -122.624167, -122.610861, -122.580889, -122.585528, 
    -122.578333, -122.567194, -122.567972, -122.575389, -122.573806, 
    -122.586306, -122.592972, -122.587083, -122.597556, -122.615028, 
    -122.614611, -122.620417, -122.617556, -122.605889, -122.596306, 
    -122.588389, -122.558389, -122.5375, -122.524611, -122.527083, 
    -122.512972, -122.513833, -122.507167, -122.506306, -122.500056, 
    -122.483306, -122.482111, -122.493361, -122.506333, -122.500917, 
    -122.482194, -122.477944, -122.471278, -122.470444, -122.473361, 
    -122.487528, -122.551722, -122.550472, -122.582972, -122.582194, -122.59, 
    -122.605028, -122.606333, -122.615861, -122.627556, -122.629611, 
    -122.62375, -122.644167, -122.652528, -122.654639, -122.660444, 
    -122.652139, -122.650889, -122.645028, -122.640083, -122.636306, 
    -122.639611, -122.631667, -122.634639, -122.631694, -122.620889, 
    -122.615417, -122.618778, -122.612972, -122.615472, -122.600917, 
    -122.591278, -122.597139, -122.592972, -122.602472, -122.610889, 
    -122.616722, -122.630889, -122.644972, -122.662111, -122.6625, 
    -122.677972, -122.674639, -122.684222, -122.6925, -122.692194, 
    -122.702111, -122.709611, -122.705833, -122.697556, -122.694222, 
    -122.687167, -122.686278, -122.692111, -122.686306, -122.688806, 
    -122.684639, -122.678833, -122.680472, -122.6775, -122.672556, 
    -122.667556, -122.662111, -122.665417, -122.6625, -122.655, -122.646722, 
    -122.633361, -122.622111, -122.625056, -122.653361, -122.670917, 
    -122.676722, -122.693778, -122.685861, -122.672583, -122.6625, 
    -122.64925, -122.637583, -122.627528, -122.6225, -122.606722, 
    -122.588389, -122.569278, -122.554222, -122.548861, -122.543778, 
    -122.551278, -122.538361, -122.532167, -122.542083, -122.539583, 
    -122.545417, -122.523417, -122.518389, -122.503389, -122.494583, 
    -122.517944, -122.522111, -122.530472, -122.534639, -122.533, 
    -122.549639, -122.553, -122.549639, -122.538806, -122.57175, -122.585, 
    -122.591333, -122.576278, -122.569583, -122.547944, -122.554611, 
    -122.570278, -122.5555, -122.532167, -122.532111, -122.549667, 
    -122.544167, -122.535028, -122.516722, -122.510028, -122.485, 
    -122.452556, -122.433333, -122.437167, -122.430917, -122.421694, 
    -122.426333, -122.419167, -122.421306, -122.418333, -122.405444, 
    -122.412944, -122.410861, -122.400889, -122.396278, -122.405833, 
    -122.410028, -122.423389, -122.434222, -122.445917, -122.444222, 
    -122.435861, -122.425111, -122.408417, -122.392528, -122.380028, 
    -122.374278, -122.335056, -122.32625, -122.323806, -122.327944, 
    -122.349611, -122.356722, -122.365083, -122.382972, -122.368806, 
    -122.3705, -122.361278, -122.365389, -122.3875, -122.39875, -122.394611, 
    -122.401278, -122.39625, -122.402083, -122.412056, -122.422111, 
    -122.384222, -122.371722, -122.36175, -122.360056, -122.358417, 
    -122.345889, -122.344222, -122.339667, -122.34675, -122.374222, 
    -122.381667, -122.385028, -122.400889, -122.411722, -122.423389, 
    -122.437944, -122.413361, -122.403778, -122.410444, -122.405444, 
    -122.406333, -122.384194, -122.377139, -122.374583, -122.384639, 
    -122.382167, -122.395472, -122.397167, -122.393, -122.394639, 
    -122.385833, -122.353389, -122.337917, -122.330444, -122.333778, 
    -122.327944, -122.322139, -122.311306, -122.313028, -122.30675, 
    -122.282556, -122.255889, -122.23675, -122.219583, -122.219583, 
    -122.225056, -122.227167, -122.218333, -122.215472, -122.226306, 
    -122.217167, -122.213, -122.215167, -122.20675, -122.194278, -122.182611, 
    -122.178417, -122.178028, -122.179667, -122.196833, -122.201028, 
    -122.208917, -122.207611, -122.193917, -122.209306, -122.211389, 
    -122.205972, -122.211806, -122.227694, -122.228472, -122.243472, 
    -122.268472, -122.292667, -122.293444, -122.281833, -122.285556, 
    -122.275972, -122.273889, -122.281, -122.291833, -122.296778, 
    -122.301806, -122.321778, -122.328417, -122.3455, -122.348833, 
    -122.364722, -122.363, -122.370556, -122.365528, -122.364722, 
    -122.372278, -122.355556, -122.358889, -122.357194, -122.362972, 
    -122.366333, -122.372667, -122.384639, -122.381778, -122.387667, 
    -122.39175, -122.395167, -122.410167, -122.425167, -122.429278, 
    -122.450167, -122.453889, -122.451333, -122.448472, -122.443, 
    -122.441361, -122.458444, -122.46425, -122.466028, -122.476778, 
    -122.475944, -122.466361, -122.476333, -122.478861, -122.473861, 
    -122.474694, -122.465556, -122.460528, -122.450083, -122.440944, 
    -122.427583, -122.421778, -122.411028, -122.383417, -122.366389, 
    -122.359667, -122.3585, -122.377639, -122.388472, -122.393861, 
    -122.400917, -122.415972, -122.425111, -122.445139, -122.468417, 
    -122.478417, -122.487611, -122.493417, -122.500944, -122.510972, 
    -122.52475, -122.532222, -122.538889, -122.534667, -122.541389, 
    -122.534694, -122.52925, -122.500972, -122.492639, -122.482639, 
    -122.473833, -122.469278, -122.45925, -122.430972, -122.417667, 
    -122.414278, -122.395944, -122.398889, -122.394722, -122.394694, 
    -122.38975, -122.388444, -122.389667, -122.381389, -122.383861, 
    -122.376389, -122.385583, -122.38225, -122.394278, -122.396361, 
    -122.388444, -122.399278, -122.402583, -122.421778, -122.420917, 
    -122.425139, -122.432611, -122.444278, -122.455194, -122.478944, 
    -122.475083, -122.468444, -122.446833, -122.466806, -122.478472, 
    -122.489306, -122.491806, -122.491778, -122.49675, -122.500972, 
    -122.503917, -122.502167, -122.507667, -122.506389, -122.4985, 
    -122.508056, -122.510194, -122.520944, -122.521778, -122.534306, 
    -122.535556, -122.555556, -122.555528, -122.572222, -122.570944, 
    -122.559694, -122.549722, -122.549333, -122.555889, -122.567667, 
    -122.571, -122.5785, -122.579722, -122.596778, -122.609306, -122.614306, 
    -122.624306, -122.629306, -122.636806, -122.651806, -122.656778, 
    -122.658889, -122.651417, -122.654222, -122.665056, -122.666833, 
    -122.677278, -122.67975, -122.668472, -122.662194, -122.663889, 
    -122.65475, -122.658944, -122.665528, -122.667222, -122.677639, 
    -122.680194, -122.686, -122.702639, -122.703028, -122.688417, 
    -122.671778, -122.614306, -122.603472, -122.598833, -122.598472, 
    -122.606806, -122.6105, -122.594722, -122.587222, -122.591333, 
    -122.584361, -122.574306, -122.572222, -122.573917, -122.579722, 
    -122.576361, -122.579333, -122.581361, -122.570139, -122.558528, 
    -122.538833, -122.5235, -122.517639, -122.515139, -122.516, -122.510972, 
    -122.50175, -122.500944, -122.4985, -122.488444, -122.483444, -122.491, 
    -122.478389, -122.473833, -122.476333, -122.470583, -122.470583, 
    -122.483111, -122.487222, -122.480639, -122.483889, -122.48725, 
    -122.498056, -122.501361, -122.505111, -122.524306, -122.540139, 
    -122.560111, -122.558083, -122.562194, -122.555917, -122.551806, 
    -122.540111, -122.496806, -122.488139, -122.496417, -122.492667, 
    -122.490111, -122.4835, -122.470111, -122.468444, -122.460083, 
    -122.468889, -122.465556, -122.468889, -122.468833, -122.457667, 
    -122.45175, -122.456361, -122.446, -122.444306, -122.438444, -122.432222, 
    -122.428, -122.440111, -122.454333, -122.469278, -122.491806, 
    -122.495972, -122.505083, -122.512222, -122.510972, -122.500944, 
    -122.491389, -122.4955, -122.501389, -122.497972, -122.506806, 
    -122.505556, -122.509222, -122.521417, -122.516778, -122.509722, 
    -122.508056, -122.493861, -122.495556, -122.48925, -122.491417, 
    -122.527583, -122.54175, -122.569306, -122.576778, -122.573917, 
    -122.57675, -122.580972, -122.585944, -122.600139, -122.609694, 
    -122.610083, -122.636417, -122.650889, -122.654278, -122.660556, 
    -122.66675, -122.674278, -122.676417, -122.662222, -122.657194, 
    -122.649722, -122.647556, -122.661806, -122.6785, -122.69675, 
    -122.702639, -122.707194, -122.704806, -122.714278, -122.712222, 
    -122.719722, -122.7485, -122.778444, -122.790111, -122.796417, 
    -122.782611, -122.770972, -122.755083, -122.748889, -122.750583, 
    -122.771778, -122.788444, -122.796, -122.821833, -122.825556, 
    -122.819306, -122.776833, -122.771361, -122.77425, -122.786028, 
    -122.790528, -122.775972, -122.750083, -122.736833, -122.733444, 
    -122.736389, -122.731361, -122.752694, -122.759301454927, -122.773361, 
    -122.824194, -122.864167, -122.875, -122.889611, -122.880944, 
    -122.876306, -122.881278, -122.878389, -122.859611, -122.863361, 
    -122.900889, -122.968361, -122.986694, -123, -123.020028, -123.044222, 
    -123.057917, -123.047556, -123.032107851209, -123.02225, -123.025972, 
    -123.049333, -123.086806, -123.09021981915, -123.100917, -123.130028, 
    -123.129167, -123.104194, -123.100917, -123.098833, -123.101306, 
    -123.114222, -123.119972, -123.152472, -123.154222, -123.161333, 
    -123.160806, -123.122056, -123.154611, -123.153389, -123.135833, 
    -123.130028, -123.148361, -123.16675, -123.17875, -123.187111, 
    -123.170833, -123.167083, -123.168361, -123.151667, -123.125917, 
    -123.121722, -123.108306, -123.097528, -123.088389, -123.075389, 
    -123.081222, -123.081667, -123.08925, -123.1175, -123.121722, 
    -123.127528, -123.144222, -123.166694, -123.196667, -123.196222, 
    -123.201333, -123.155833, -123.15375, -123.155833, -123.172556, 
    -123.208361, -123.211306, -123.208361, -125.815889, -128.475, -133.35425, 
    -134, -134, -134, -134, -134, -134, -130.298861, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, NaN, -114, 
    NaN, -125.672556, -125.672167, -125.672167, -125.677111, -125.673806, 
    -125.693778, -125.685, -125.688361, -125.705889, -125.743333, 
    -125.765056, -125.780028, -125.785056, -125.799194, -125.810861, 
    -125.815028, -125.82, -125.829194, -125.852556, -125.858361, -125.874167, 
    -125.881694, -125.887972, -125.874222, -125.872972, -125.890056, 
    -125.895861, -125.900917, -125.903778, -125.9005, -125.913806, 
    -125.913806, -125.9075, -125.8875, -125.884556, -125.887972, -125.882111, 
    -125.884556, -125.880861, -125.875083, -125.867556, -125.873778, 
    -125.864222, -125.855028, -125.847139, -125.860444, -125.859583, 
    -125.852083, -125.859194, -125.845444, -125.855472, -125.84675, 
    -125.840028, -125.832111, -125.835056, -125.818361, -125.822472, 
    -125.834611, -125.833361, -125.804222, -125.78, -125.780472, -125.774194, 
    -125.767528, -125.764194, -125.758333, -125.755889, -125.74425, 
    -125.740472, -125.747528, -125.738361, -125.730833, -125.736306, 
    -125.72925, -125.724167, -125.724611, -125.755472, -125.747583, 
    -125.718417, -125.721694, -125.71425, -125.706667, -125.704222, 
    -125.696722, -125.683417, -125.674194, -125.654222, -125.671306, 
    -125.662972, -125.666667, -125.673361, -125.678722, -125.675028, 
    -125.665056, -125.648417, -125.637972, -125.634667, -125.62375, 
    -125.630944, -125.633417, -125.636333, -125.632944, -125.637528, 
    -125.638833, -125.63, -125.65, -125.653778, -125.6575, -125.664278, 
    -125.671306, -125.667139, -125.671306, -125.664583, -125.680444, 
    -125.677111, -125.682528, -125.686278, -125.685861, -125.691694, 
    -125.698389, -125.710472, -125.70125, -125.713, -125.713778, -125.724139, 
    -125.732917, -125.731333, -125.744194, -125.741306, -125.75, -125.767083, 
    -125.757944, -125.760833, -125.7775, -125.7875, -125.790889, -125.782611, 
    -125.781694, -125.770083, -125.76625, -125.769694, -125.766306, 
    -125.754611, -125.757056, -125.752528, -125.74375, -125.749583, 
    -125.747111, -125.751361, -125.752139, -123.969667, -123.956722, 
    -123.948778, -123.940417, -123.926278, -123.927056, -123.917528, 
    -123.90425, -123.893806, -123.896278, -123.88875, -123.887889, 
    -123.897111, -123.895, -123.885806, -123.864222, -123.847583, 
    -123.835861, -123.803361, -123.787528, -123.771667, -123.769222, 
    -123.814639, -123.802972, -123.803806, -123.793361, -123.776278, 
    -123.767944, -123.770083, -123.757083, -123.759667, -123.754194, 
    -123.747111, -123.747056, -123.754167, -123.762583, -123.767556, 
    -123.783333, -123.790083, -123.791361, -123.7875, -123.7775, -123.767167, 
    -123.761313895368, -123.761333, -123.758083, -123.772639, -123.771806, 
    -123.778472, -123.787583, -123.793444, -123.804391766201, 
    -123.806866557692, -123.804694, -123.806778, -123.810313641544, 
    -123.8375, -123.847556, -123.852556, -123.858, -123.855833, -123.848361, 
    -123.846667, -123.844194, -123.822321036215, -123.821833, -123.808528, 
    -123.803417, -123.778444, -123.774306, -123.771806, -123.755944, 
    -123.738917, -123.7185, -123.709306, -123.706361, -123.708833, 
    -123.705972, -123.702194, -123.698, -123.698, -123.69175, -123.690917, 
    -123.686389, -123.688056, -123.682611, -123.680139, -123.673861, 
    -123.672583, -123.678, -123.67425, -123.665972, -123.660944, -123.648444, 
    -123.636806, -123.620972, -123.616778, -123.594333, -123.588, 
    -123.584667, -123.587694, -123.600139, -123.60975, -123.600917, 
    -123.597139, -123.590111, -123.563944, -123.56475, -123.558, -123.565139, 
    -123.580583, -123.570528, -123.577639, -123.582583, -123.586778, 
    -123.597667, -123.596361, -123.604278, -123.620111, -123.631778, 
    -123.635528, -123.646389, -123.640083, -123.636361, -123.645556, 
    -123.582583, -123.557556, -123.554278, -123.534694, -123.533028, 
    -123.539278, -123.5485, -123.555083, -123.556361, -123.553111, 
    -123.530528, -123.518861, -123.523833, -123.52225, -123.514667, 
    -123.520972, -123.548472, -123.557222, -123.555556, -123.543833, 
    -123.542167, -123.548083, -123.542611, -123.535556, -123.5385, 
    -123.507639, -123.487639, -123.475917, -123.47175, -123.463, -123.471306, 
    -123.466417, -123.48225, -123.476389, -123.481333, -123.481333, 
    -123.466333, -123.470139, -123.47925, -123.479667, -123.474306, 
    -123.446444, -123.451861, -123.472611, -123.473444, -123.4785, 
    -123.482639, -123.489722, -123.483417, -123.475528, -123.475167, 
    -123.486306, -123.481806, -123.438417, -123.420139, -123.403472, 
    -123.405528, -123.40175, -123.398028, -123.397667, -123.411806, 
    -123.415056, -123.422194, -123.416, -123.414667, -123.4205, -123.409278, 
    -123.410111, -123.406778, -123.399278, -123.400917, -123.392222, 
    -123.396389, -123.393083, -123.409722, -123.388833, -123.388444, 
    -123.377639, -123.372611, -123.370528, -123.367194, -123.361389, 
    -123.364694, -123.330194, -123.317611, -123.316028, -123.305972, 
    -123.299722, -123.301361, -123.275111, -123.265556, -123.279278, 
    -123.289306, -123.298083, -123.290583, -123.291444, -123.300944, 
    -123.306361, -123.298028, -123.294306, -123.304306, -123.313417, 
    -123.320917, -123.327639, -123.333444, -123.33925, -123.350167, 
    -123.353472, -123.375944, -123.385111, -123.391361, -123.387667, 
    -123.375139, -123.370972, -123.371806, -123.396778, -123.394694, 
    -123.407611, -123.415972, -123.419306, -123.421722, -123.432556, 
    -123.433472, -123.436861, -123.440583, -123.437583, -123.4205, 
    -123.435167, -123.436389, -123.432167, -123.434306, -123.455917, 
    -123.449778, -123.450556, -123.445528, -123.447222, -123.454722, 
    -123.487222, -123.485972, -123.47925, -123.477167, -123.482639, 
    -123.502639, -123.502611, -123.513444, -123.519278, -123.543056, 
    -123.539306, -123.526361, -123.535111, -123.558833, -123.538889, 
    -123.540083, -123.55925, -123.565972, -123.57925, -123.583472, 
    -123.591778, -123.600917, -123.603083, -123.600139, -123.596778, 
    -123.593056, -123.590111, -123.593417, -123.602694, -123.60425, 
    -123.627639, -123.633056, -123.628806, -123.634722, -123.637611, 
    -123.654278, -123.654306, -123.667667, -123.685167, -123.701722, 
    -123.708444, -123.709278, -123.713472, -123.716333, -123.705111, 
    -123.703833, -123.715944, -123.717194, -123.700944, -123.68175, 
    -123.680139, -123.672556, -123.663417, -123.655917, -123.651778, 
    -123.635972, -123.638861, -123.634722, -123.647556, -123.652583, 
    -123.660472, -123.655083, -123.655139, -123.665111, -123.6785, 
    -123.683861, -123.690111, -123.6985, -123.712611, -123.723444, 
    -123.730556, -123.723528, -123.716778, -123.710472, -123.730167, 
    -123.751833, -123.765139, -123.777583, -123.785944, -123.796806, 
    -123.823472, -123.836778, -123.864306, -123.900194, -123.921778, 
    -123.93925, -123.949306, -123.980167, -123.986361, -123.991778, 
    -124.013444, -124.037556, -124.072528, -124.095889, -124.109222, 
    -124.117556, -124.158389, -124.175028, -124.207583, -124.25175, 
    -124.292556, -124.293778, -124.3125, -124.365889, -124.397583, 
    -124.400028, -124.408389, -124.419167, -124.432611, -124.443361, 
    -124.448389, -124.459611, -124.451722, -124.426722, -124.401278, 
    -124.402083, -124.4125, -124.451722, -124.469194, -124.475028, 
    -124.495889, -124.552583, -124.553361, -124.556667, -124.589167, 
    -124.610056, -124.619167, -124.648417, -124.655917, -124.679194, 
    -124.690056, -124.715861, -124.739139, -124.755083, -124.765861, 
    -124.771667, -124.778361, -124.785028, -124.800028, -124.815833, 
    -124.825, -124.830833, -124.850917, -124.855833, -124.852917, 
    -124.861667, -124.871667, -124.887583, -124.91175, -124.95, -124.975917, 
    -124.986694, -125.002528, -125.02, -125.065889, -125.101722, -125.106639, 
    -125.117972, -125.119639, -125.130417, -125.133028, -125.129222, 
    -125.128778, -125.135444, -125.134583, -125.117972, -125.118333, 
    -125.129194, -125.143778, -125.147111, -125.156694, -125.15625, 
    -125.160028, -125.162139, -125.167139, -125.167583, -125.177528, 
    -125.187556, -125.190028, -125.2, -125.204222, -125.210861, -125.217111, 
    -125.218722, -125.212944, -125.215472, -125.209972, -125.193389, 
    -125.1925, -125.184222, -125.182139, -125.187167, -125.18, -125.171694, 
    -125.170028, -125.16675, -125.163417, -125.157556, -125.144167, 
    -125.140444, -125.142917, -125.139222, -125.139611, -125.134639, 
    -125.137083, -125.13125, -125.120028, -125.114167, -125.111306, 
    -125.107111, -125.108722, -125.100056, -125.091722, -125.076667, 
    -125.077556, -125.070861, -125.053361, -125.050028, -125.050861, 
    -125.040056, -125.033306, -125.032944, -125.026694, -125.005417, 
    -125.004167, -125.013833, -125.005389, -125.009194, -125.010056, 
    -125.016639, -125.018333, -125.024278, -125.025806, -125.029167, 
    -125.034583, -125.037111, -125.026278, -125.035444, -125.030472, 
    -125.031694, -125.023417, -125.021639, -125.00425, -125.005861, 
    -124.986611, -124.988722, -124.980333, -124.990389, -124.983278, 
    -124.983278, -124.969194, -124.950778, -124.948306, -124.907472, 
    -124.898333, -124.894556, -124.884139, -124.864222, -124.864222, 
    -124.855472, -124.84125, -124.835444, -124.838, -124.832917, -124.813778, 
    -124.817111, -124.810472, -124.812944, -124.787111, -124.792972, 
    -124.791278, -124.80675, -124.814639, -124.810472, -124.82625, 
    -124.822139, -124.829639, -124.825083, -124.807139, -124.813861, 
    -124.825083, -124.823, -124.832972, -124.830111, -124.851694, 
    -124.852556, -124.863361, -124.882167, -124.878389, -124.8605, 
    -124.863778, -124.870889, -124.891163735156, -124.897472, -124.914139, 
    -124.938278, -124.956583, -124.971667, -124.974917, -124.975806, 
    -124.984917, -124.987833, -124.978722, -124.981639, -124.993253834092, 
    -125.032167, -125.022944, -125.02675, -125.033306, -125.045833, 
    -125.04625, -125.012926, -125.013778, -125.000833, -124.993639, 
    -125.002556, -125.015056, -125.024222, -125.030917, -125.034583, 
    -125.033778, -125.020472, -125.028361, -125.033389, -125.039194, 
    -125.036722, -125.040083, -125.04175, -125.047111, -125.049167, 
    -125.065056, -125.083361, -125.082139, -125.087139, -125.087528, 
    -125.09675, -125.104194, -125.114222, -125.121667, -125.128778, 
    -125.127056, -125.133806, -125.137417836421, -125.142756270286, 
    -125.142528, -125.150417, -125.150186936053, -125.140444, -125.146722, 
    -125.1560803059, -125.155472, -125.163417, -125.16675, -125.171694, 
    -125.186694, -125.187556, -125.178306, -125.177979864954, -125.148806, 
    -125.148806, -125.136333, -125.142111, -125.138306, -125.136278, 
    -125.150806, -125.1625, -125.167528, -125.197472, -125.213778, 
    -125.173333, -125.165056, -125.151222, -125.143778, -125.150889, 
    -125.153444, -125.161667, -125.168778, -125.154639, -125.154556, 
    -125.164972, -125.176722, -125.177583, -125.180833, -125.185861, 
    -125.193045925887, -125.195389, -125.18375, -125.193806, -125.189556, 
    -125.194667, -125.192972, -125.199194, -125.200861, -125.2055, 
    -125.200028, -125.206306, -125.212611, -125.227917, -125.21625, 
    -125.210389, -125.214167, -125.223306, -125.245028, -125.251278, 
    -125.250861, -125.275056, -125.278833, -125.272111, -125.273417, 
    -125.279611, -125.280056, -125.286639, -125.288722, -125.2825, 
    -125.277583, -125.283389, -125.285056, -125.303361, -125.312556, 
    -125.3175, -125.324222, -125.323333, -125.3025, -125.291306, -125.295417, 
    -125.298, -125.304503309505, -125.322139, -125.309139, -125.293444, 
    -125.290056, -125.28, -125.280056, -125.275028, -125.274194, -125.251694, 
    -125.206667, -125.199167, -125.218417, -125.225, -125.262583, 
    -125.293389, -125.301722, -125.303389, -125.308333, -125.313333, 
    -125.329194, -125.335056, -125.348361, -125.353333, -125.360917, 
    -125.354639, -125.3605, -125.367270458015, -125.3675, -125.393306, 
    -125.392111, -125.396639, -125.417528, -125.426667, -125.434167, 
    -125.444167, -125.445833, -125.460056, -125.46875, -125.480056, 
    -125.483417, -125.483361, -125.505, -125.500528, -125.502556, 
    -125.506778, -125.51175, -125.517528, -125.521333, -125.517917, 
    -125.524194, -125.528444, -125.547556, -125.559222, -125.576722, 
    -125.580028, -125.586306, -125.585444, -125.591278, -125.570056, 
    -125.567111, -125.575083, -125.568361, -125.565889, -125.561639, 
    -125.555889, -125.550028, -125.527917, -125.535472, -125.528, 
    -125.530917, -125.546694, -125.548722, -125.541222, -125.545444, 
    -125.544222, -125.551722, -125.555833, -125.576667, -125.579194, 
    -125.586639, -125.590861, -125.593361, -125.596361, -125.593417, 
    -125.607194, -125.603778, -125.610444, -125.609667, -125.615, 
    -125.619583, -125.61925, -125.614611, -125.613778, -125.635056, 
    -125.632912545383, -125.657963732562, -125.658778, -125.657556, 
    -125.665056, -125.66675, -125.672556, -125.674167, -125.672556, NaN, 
    -114.324167, -114.3275, -114.336944, -114.339722, -114.343333, 
    -114.352778, -114.355278, -114.3475, -114.349167, -114.353889, 
    -114.360556, -114.369167, -114.390833, -114.400556, -114.4075, -114.41, 
    -114.411944, -114.398611, -114.4, -114.3925, -114.38, -114.374444, 
    -114.367778, -114.364167, -114.369167, -114.409167, -114.420833, 
    -114.433333, -114.441389, -114.439444, -114.428889, -114.427222, 
    -114.432222, -114.418889, -114.415, -114.413056, -114.42, -114.440833, 
    -114.450556, -114.449444, -114.460278, -114.481389, -114.518611, 
    -114.565, -114.605556, -114.635, -114.659444, -114.686389, -114.699722, 
    -114.708056, -114.721667, -114.716111, -114.719167, -114.745556, 
    -114.766667, -114.774444, -114.805833, -114.832222, -114.856111, -114.86, 
    -114.857222, -114.828889, -114.805, -114.800556, -114.813056, -114.81, 
    -114.796111, -114.765, -114.732222, -114.727778, -114.741389, 
    -114.734722, -114.715278, -114.696111, -114.710556, -114.700833, 
    -114.665833, -114.655278, -114.637222, -114.6325, -114.623889, 
    -114.572778, -114.561944, -114.55, -114.542222, -114.516944, -114.503611, 
    -114.491389, -114.459167, -114.455556, -114.456389, -114.450833, 
    -114.443056, -114.4325, -114.413056, -114.393056, -114.390556, 
    -114.403611, -114.401944, -114.395833, -114.374167, -114.375, 
    -114.358333, -114.351389, -114.3475, -114.334444, -114.322222, 
    -114.319444, -114.33, -114.281944, -114.252778, -114.235, -114.196944, 
    -114.155, -114.110278, -114.107222, -114.08, -114.084444, -114.071944, 
    -114.053056, -114.039722, -114.016944, -114.001111, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, -114, 
    -114, -114, -114, -114, -114, -114, -114, -114.002778, -114.007222, 
    -114.017778, -114.019722, -114.026944, -114.058056, -114.072222, 
    -114.103889, -114.1225, -114.142778, -114.144722, -114.154167, 
    -114.180833, -114.210556, -114.225556, -114.251944, -114.255556, 
    -114.2575, -114.253611, -114.245, -114.246944, -114.282778, -114.286389, 
    -114.298889, -114.308056, -114.330556, -114.352222, -114.370278, 
    -114.381111, -114.3875, -114.3875, -114.370278, -114.373056, -114.365833, 
    -114.343056, -114.316944, -114.309722, -114.314167, -114.3275, 
    -114.329167, -114.335, -114.333889, -114.323611, -114.332222, 
    -114.324167, NaN, -122.371722, -122.370111, -122.353, -122.347972, 
    -122.357972, -122.374667, -122.378389, -122.39625, -122.395472, 
    -122.387583, -122.402472, -122.416694, -122.430861, -122.444667, 
    -122.446333, -122.441306, -122.443806, -122.454972, -122.475, 
    -122.484222, -122.498389, -122.513361, -122.523417, -122.546694, 
    -122.552972, -122.5455, -122.542056, -122.560944, -122.585083, -122.601, 
    -122.608028, -122.598861, -122.5955, -122.598, -122.614778, -122.599722, 
    -122.610611, -122.61925, -122.631, -122.661028, -122.670917, -122.673472, 
    -122.675139, -122.680083, -122.692667, -122.712639, -122.737639, 
    -122.747583, -122.761806, -122.767222, -122.770583, -122.753861, 
    -122.733917, -122.724694, -122.693056, -122.669694, -122.6655, 
    -122.665139, -122.63425, -122.63225, -122.637194, -122.628472, 
    -122.611833, -122.598444, -122.594333, -122.587639, -122.58475, 
    -122.586417, -122.579639, -122.595194, -122.564278, -122.530944, 
    -122.525111, -122.514306, -122.505556, -122.505556, -122.527611, 
    -122.558444, -122.559306, -122.563889, -122.561389, -122.584361, 
    -122.602639, -122.624278, -122.627222, -122.622194, -122.625972, 
    -122.632639, -122.643083, -122.646861, -122.633056, -122.636806, 
    -122.645944, -122.663917, -122.652194, -122.653056, -122.660111, 
    -122.674333, -122.713472, -122.7285, -122.734306, -122.732222, 
    -122.726333, -122.722611, -122.715944, -122.693444, -122.680972, 
    -122.673472, -122.660167, -122.647556, -122.645972, -122.635139, 
    -122.627611, -122.605556, -122.603, -122.597667, -122.587222, 
    -122.580583, -122.567194, -122.566361, -122.558917, -122.572167, 
    -122.556444, -122.54725, -122.549722, -122.540111, -122.537194, 
    -122.540972, -122.528444, -122.520972, -122.512222, -122.518028, 
    -122.513889, -122.527194, -122.52425, -122.506806, -122.491778, 
    -122.445139, -122.430972, -122.406778, -122.400111, -122.376833, 
    -122.371722, NaN, -123.000972, -123.004222, -123.023417, -123.030944, 
    -123.040139, -123.052583, -123.066361, -123.06975, -123.063861, 
    -123.065111, -123.072639, -123.077639, -123.075972, -123.084222, 
    -123.094278, -123.105167, -123.1085, -123.110111, -123.119333, 
    -123.133417, -123.143, -123.146806, -123.153861, -123.153861, 
    -123.164722, -123.163111, -123.169694, -123.178889, -123.172611, 
    -123.163417, -123.158, -123.154306, -123.163417, -123.165139, 
    -123.173944, -123.172167, -123.165111, -123.161806, -123.153444, 
    -123.150972, -123.151306, -123.158861, -123.147639, -123.138889, 
    -123.144306, -123.150917, -123.160167, -123.164278, -123.173028, 
    -123.172194, -123.166361, -123.167667, -123.163444, -123.156806, 
    -123.153056, -123.158889, -123.152194, -123.152667, -123.141, 
    -123.140139, -123.148056, -123.143389, -123.120917, -123.119278, 
    -123.102556, -123.098056, -123.10425, -123.082611, -123.076861, 
    -123.05925, -123.04925, -123.035167, -123.014306, -123.007167, 
    -123.007167, -123.017694, -123.019306, -123.007583, -122.998444, 
    -122.996417, -122.988472, -122.9835, -122.979278, -122.9705, -122.973444, 
    -122.983417, -122.996806, -123.005083, -123.015167, -123.016833, 
    -123.021333, -123.021333, -123.016361, -123.022194, -123.022194, 
    -123.008028, -123.011361, -123.007583, -122.989306, -122.970972, 
    -122.96675, -122.971833, -122.960611, -122.964278, -123.000972, NaN, 
    -122.947167, -122.947167, -122.934778, -122.926722, -122.919694, 
    -122.923028, -122.91925, -122.931833, -122.936861, -122.932611, 
    -122.929361, -122.921778, -122.915583, -122.914694, -122.918917, 
    -122.923861, -122.92225, -122.908472, -122.902583, -122.894333, 
    -122.892222, -122.885111, -122.88425, -122.874278, -122.8735, 
    -122.866417, -122.866389, -122.875583, -122.877222, -122.874306, 
    -122.861833, -122.853083, -122.860583, -122.867167, -122.875528, 
    -122.851472, -122.857194, -122.856417, -122.862222, -122.85675, 
    -122.845139, -122.843889, -122.854722, -122.848444, -122.840972, 
    -122.830111, -122.824694, -122.832278, -122.829639, -122.833444, 
    -122.83475, -122.819306, -122.813861, -122.81975, -122.815194, -122.806, 
    -122.801417, -122.809722, -122.81475, -122.805139, -122.805056, 
    -122.817611, -122.829278, -122.82925, -122.834361, -122.843417, 
    -122.840944, -122.861833, -122.862667, -122.850611, -122.85675, 
    -122.85675, -122.871806, -122.878472, -122.895972, -122.895972, 
    -122.880556, -122.8805, -122.890139, -122.890139, -122.875944, 
    -122.876389, -122.870972, -122.865528, -122.878417, -122.894306, 
    -122.895167, -122.897639, -122.901778, -122.909333, -122.913444, 
    -122.903056, -122.910111, -122.918833, -122.913417, -122.919306, 
    -122.927583, -122.928444, -122.931833, -122.936778, -122.942667, 
    -122.947167, NaN, -123.598861, -123.598917, -123.593028, -123.595889, 
    -123.575944, -123.546778, -123.528444, -123.504306, -123.498056, 
    -123.503389, -123.495139, -123.494333, -123.426806, -123.421, 
    -123.452639, -123.463472, -123.47425, -123.4805, -123.47425, -123.468417, 
    -123.428444, -123.425556, -123.4285, -123.44675, -123.444278, 
    -123.469333, -123.488472, -123.4855, -123.490167, -123.500583, 
    -123.494333, -123.482583, -123.487222, -123.484278, -123.474306, 
    -123.469278, -123.455111, -123.432667, -123.427583, -123.421778, 
    -123.407639, -123.394222, -123.390139, -123.380167, -123.375583, 
    -123.367167, -123.374278, -123.379778, -123.381389, -123.388444, 
    -123.395083, -123.399278, -123.405139, -123.414306, -123.430972, 
    -123.444278, -123.460917, -123.4485, -123.435583, -123.426361, 
    -123.476806, -123.500972, -123.525111, -123.550111, -123.563944, 
    -123.562583, -123.54925, -123.5455, -123.553889, -123.550139, 
    -123.540111, -123.525139, -123.518861, -123.559333, -123.570083, 
    -123.573, -123.570139, -123.563444, -123.563028, -123.550944, 
    -123.532167, -123.573417, -123.581417, -123.578833, -123.593056, 
    -123.589667, -123.593028, -123.588083, -123.5955, -123.598861, NaN, 
    -123.000528, -123.000528, -123.005972, -123.008889, -123.024222, 
    -123.031389, -123.032167, -123.021389, -123.010972, -122.991806, 
    -122.982667, -122.962639, -122.95975, -122.962639, -122.950167, 
    -122.943056, -122.950972, -122.925944, -122.910167, -122.895972, 
    -122.885111, -122.878444, -122.868472, -122.854333, -122.828444, 
    -122.826861, -122.804361, -122.801806, -122.74225, -122.755111, 
    -122.756389, -122.76675, -122.780139, -122.781778, -122.788917, 
    -122.784278, -122.799722, -122.799639, -122.810528, -122.800167, 
    -122.817667, -122.825944, -122.829278, -122.832583, -122.833444, 
    -122.838472, -122.842583, -122.845972, -122.869333, -122.875944, 
    -122.88225, -122.887222, -122.901806, -122.902583, -122.909306, 
    -122.925556, -122.918056, -122.912194, -122.912222, -122.907611, 
    -122.895167, -122.883028, -122.878, -122.863917, -122.866, -122.881778, 
    -122.88675, -122.889278, -122.903472, -122.906806, -122.907611, 
    -122.915972, -122.936778, -122.938417, -122.950167, -122.958056, 
    -122.953028, -122.960139, -122.971833, -122.984306, -122.993889, 
    -122.987611, -122.989694, -122.980556, -122.979333, -122.992583, 
    -122.99475, -123.000528, NaN, -116.531111, -116.530833, -116.523889, 
    -116.507778, -116.505278, -116.515278, -116.5475, -116.550278, 
    -116.546389, -116.561944, -116.559722, -116.531111, -116.485, 
    -116.445556, -116.430278, -116.429722, -116.434444, -116.449722, 
    -116.451111, -116.438333, -116.415556, -116.415278, -116.410556, 
    -116.383056, -116.288056, -116.275, -116.263889, -116.2575, -116.2125, 
    -116.190278, -116.190833, -116.209167, -116.225, -116.25, -116.254444, 
    -116.255833, -116.275556, -116.279167, -116.277222, -116.301667, 
    -116.350833, -116.358611, -116.391667, -116.405556, -116.420556, 
    -116.430833, -116.441111, -116.466667, -116.489444, -116.507778, 
    -116.523611, -116.550278, -116.570278, -116.572222, -116.557222, 
    -116.523333, -116.514167, -116.503056, -116.4875, -116.464444, 
    -116.458056, -116.448889, -116.432222, -116.426944, -116.421389, 
    -116.401944, -116.391667, -116.381389, -116.359444, -116.354722, 
    -116.370556, -116.378889, -116.395278, -116.4175, -116.435833, 
    -116.445833, -116.470556, -116.516667, -116.531111, NaN, -119.593444, 
    -119.596944, -119.658972, -119.692611, -119.700556, -119.702694, 
    -119.708139, -119.717139, -119.723694, -119.744833, -119.755944, 
    -119.760167, -119.772944, -119.791222, -119.795917, -119.809, -119.8185, 
    -119.841528, -119.852083, -119.866472, -119.877028, -119.888444, 
    -119.880222, -119.8775, -119.885583, -119.898667, -119.915917, 
    -119.925972, -119.931, -119.921222, -119.924139, -119.921694, 
    -119.919333, -119.911111, -119.892889, -119.882444, -119.865472, 
    -119.857639, -119.825444, -119.818556, -119.814611, -119.811056, 
    -119.800694, -119.798444, -119.76725, -119.766222, -119.759806, 
    -119.754389, -119.748, -119.737472, -119.726833, -119.712278, -119.70325, 
    -119.691528, -119.686111, -119.676083, -119.669028, -119.654389, 
    -119.651667, -119.638222, -119.618028, -119.6065, -119.610722, 
    -119.610056, -119.588361, -119.576, -119.563917, -119.556222, -119.5315, 
    -119.521611, -119.528139, -119.543417, -119.546861, -119.557611, 
    -119.578056, -119.593444, NaN, -122.208889, -122.211389, -122.218056, 
    -122.224444, -122.226667, -122.236111, -122.257222, -122.261389, 
    -122.2875, -122.298611, -122.311667, -122.325556, -122.339167, 
    -122.350278, -122.359167, -122.353333, -122.332778, -122.33, -122.370833, 
    -122.400833, -122.385278, -122.3775, -122.389444, -122.407222, 
    -122.414444, -122.415833, -122.425556, -122.442222, -122.445, 
    -122.440556, -122.418056, -122.4075, -122.401111, -122.391111, 
    -122.381389, -122.371111, -122.286944, -122.264167, -122.243611, 
    -122.231667, -122.225833, -122.2175, -122.199167, -122.1775, -122.14, 
    -122.110278, -122.093333, -122.093056, -122.101111, -122.136667, 
    -122.152222, -122.165556, -122.191111, -122.195556, -122.193611, 
    -122.1675, -122.164444, -122.166944, -122.175278, -122.201944, 
    -122.228056, -122.240833, -122.266389, -122.274167, -122.276389, 
    -122.270556, -122.244167, -122.243333, -122.216111, -122.208889, NaN, 
    -114.157222, -114.160556, -114.164722, -114.156944, -114.107222, 
    -114.088333, -114.060833, -114.046111, -114.041111, -114.037222, 
    -114.063889, -114.068056, -114.064722, -114.059167, -114.054722, 
    -114.048056, -114.040556, -114.037222, -114.029444, -114.0175, 
    -114.008889, -114, -114, -114.019722, -114.015833, -114.021111, 
    -114.0475, -114.058611, -114.068611, -114.080833, -114.097778, -114.105, 
    -114.112778, -114.1175, -114.123889, -114.128333, -114.146389, -114.2, 
    -114.207778, -114.208889, -114.195556, -114.158611, -114.157778, 
    -114.140278, -114.143333, -114.153333, -114.1725, -114.178889, 
    -114.199167, -114.244167, -114.256111, -114.265, -114.274444, 
    -114.316667, -114.318611, -114.2975, -114.285, -114.24, -114.214167, 
    -114.1675, -114.151944, -114.143056, -114.131944, -114.122778, 
    -114.119444, -114.108333, -114.106111, -114.116389, -114.150278, 
    -114.157222, NaN, -118.307556, -118.309222, -118.306444, -118.315528, 
    -118.316583, -118.322, -118.328583, -118.340139, -118.348, -118.363278, 
    -118.365667, -118.351583, -118.355833, -118.367194, -118.367639, 
    -118.353389, -118.331667, -118.320694, -118.315861, -118.303111, 
    -118.294194, -118.286806, -118.277722, -118.265861, -118.258028, 
    -118.257389, -118.265722, -118.270833, -118.276361, -118.284222, 
    -118.284111, -118.278556, -118.270639, -118.251528, -118.225611, 
    -118.219111, -118.227306, -118.225583, -118.22775, -118.219, -118.226778, 
    -118.225583, -118.238333, -118.245, -118.24975, -118.248472, -118.262194, 
    -118.267917, -118.273528, -118.28025, -118.299667, -118.297333, 
    -118.299028, -118.2875, -118.283972, -118.288917, -118.289083, 
    -118.295778, -118.296417, -118.303556, -118.297472, -118.295944, 
    -118.300778, -118.295972, -118.293167, -118.2935, -118.316472, 
    -118.30775, -118.307556, NaN, -121.934722, -121.938889, -121.945278, 
    -121.951667, -121.956389, -121.944444, -121.945833, -121.950833, 
    -121.966667, -121.977222, -121.9725, -121.975556, -121.994722, 
    -121.998611, -121.9975, -122.003889, -122.016944, -122.042222, 
    -122.048056, -122.057778, -122.080278, -122.0825, -122.049167, 
    -122.038056, -122.025556, -122.010833, -121.997222, -121.984167, 
    -121.974167, -121.968611, -121.961111, -121.954444, -121.942778, 
    -121.932778, -121.901667, -121.905833, -121.910833, -121.944722, 
    -121.944722, -121.939722, -121.927778, -121.909444, -121.893611, 
    -121.880556, -121.8525, -121.835278, -121.819722, -121.811389, 
    -121.804722, -121.820833, -121.8275, -121.818333, -121.826389, 
    -121.816111, -121.813333, -121.825, -121.898889, -121.915556, 
    -121.948333, -121.961389, -121.983889, -121.983333, -121.976389, 
    -121.946111, -121.934167, -121.925833, -121.934722, NaN, -118.607139, 
    -118.607083, -118.585, -118.569194, -118.550889, -118.538333, 
    -118.530028, -118.523361, -118.522528, -118.503333, -118.498333, 
    -118.478389, -118.473361, -118.463361, -118.445056, -118.424194, 
    -118.396722, -118.389139, -118.38, -118.370889, -118.367111, -118.370444, 
    -118.367944, -118.35875, -118.353361, -118.331278, -118.324583, 
    -118.326333, -118.3175, -118.310417, -118.303778, -118.304611, 
    -118.317528, -118.330861, -118.350028, -118.355, -118.375833, 
    -118.413389, -118.420833, -118.442528, -118.466667, -118.482917, 
    -118.491278, -118.484583, -118.487139, -118.48125, -118.481667, 
    -118.47625, -118.482917, -118.489611, -118.506639, -118.507917, 
    -118.504167, -118.512917, -118.513361, -118.525, -118.536694, 
    -118.537556, -118.564167, -118.565861, -118.575417, -118.57375, 
    -118.585861, -118.595861, -118.602556, -118.607139, NaN, -115.365806, 
    -115.365528, -115.356917, -115.356917, -115.352389, -115.350194, 
    -115.3275, -115.315528, -115.292639, -115.2625, -115.251722, -115.250944, 
    -115.247472, -115.259056, -115.267444, -115.270778, -115.28, -115.267611, 
    -115.268444, -115.271056, -115.265139, -115.264222, -115.253222, 
    -115.2315, -115.218306, -115.21325, -115.213333, -115.191639, 
    -115.187556, -115.178389, -115.179194, -115.170722, -115.171861, 
    -115.160917, -115.150778, -115.153361, -115.150833, -115.153222, 
    -115.167639, -115.173417, -115.169139, -115.172639, -115.168167, 
    -115.171056, -115.182694, -115.183306, -115.177306, -115.179333, 
    -115.185, -115.191, -115.203167, -115.231278, -115.237417, -115.243306, 
    -115.255222, -115.252278, -115.258306, -115.265889, -115.276528, 
    -115.293389, -115.302528, -115.321083, -115.338583, -115.350694, 
    -115.365806, NaN, -120, -119.99875, -119.987278, -119.978972, 
    -119.980556, -119.969361, -119.999389, -120.018611, -120.023139, 
    -120.048583, -120.048722, -120.07, -120.081472, -120.099528, -120.108611, 
    -120.109278, -120.117806, -120.134722, -120.137917, -120.152972, 
    -120.159944, -120.162139, -120.16725, -120.173, -120.180722, -120.189806, 
    -120.199556, -120.209778, -120.221639, -120.224222, -120.238361, 
    -120.242556, -120.248778, -120.252167, -120.242833, -120.239528, 
    -120.228861, -120.209528, -120.195944, -120.186528, -120.177611, 
    -120.166278, -120.152722, -120.149417, -120.139917, -120.11975, 
    -120.116222, -120.092861, -120.075861, -120.055972, -120.043833, 
    -120.043028, -120.049611, -120.046472, -120.039667, -120.015667, 
    -120.012361, -120, NaN, -122.594667, -122.594611, -122.575861, 
    -122.571306, -122.57, -122.564167, -122.559611, -122.565417, -122.566306, 
    -122.564639, -122.555833, -122.548361, -122.541694, -122.530389, 
    -122.531722, -122.535028, -122.543444, -122.545917, -122.543333, 
    -122.528361, -122.524194, -122.519194, -122.510028, -122.503778, 
    -122.509639, -122.497972, -122.518778, -122.490028, -122.493028, 
    -122.489611, -122.495111, -122.500861, -122.515139, -122.519972, 
    -122.525111, -122.538361, -122.538806, -122.518389, -122.500917, 
    -122.496278, -122.497917, -122.515444, -122.483417, -122.480833, 
    -122.508333, -122.523417, -122.537111, -122.544222, -122.54925, 
    -122.555889, -122.564194, -122.570861, -122.577944, -122.575472, 
    -122.579639, -122.594667, NaN, -120.123889, -120.121111, -120.065833, 
    -120.018056, -119.998889, -119.979722, -120.01, -120.037778, -120.051944, 
    -120.11, -120.154722, -120.172222, -120.179167, -120.168889, -120.169722, 
    -120.185278, -120.2075, -120.250556, -120.278333, -120.336389, 
    -120.382778, -120.433056, -120.457778, -120.474444, -120.510278, 
    -120.5225, -120.562222, -120.591111, -120.627222, -120.644444, 
    -120.656389, -120.663611, -120.665833, -120.6575, -120.633611, 
    -120.628611, -120.616111, -120.575833, -120.565278, -120.546389, 
    -120.513056, -120.499444, -120.482778, -120.462778, -120.448333, 
    -120.416944, -120.330556, -120.259167, -120.233611, -120.219167, 
    -120.204722, -120.199722, -120.202222, -120.177222, -120.123889, NaN, 
    -115.775833, -115.786944, -115.829444, -115.881667, -115.891667, 
    -115.894167, -115.899722, -115.910833, -115.925278, -115.961667, 
    -115.989722, -116.016944, -116.041389, -116.088333, -116.121667, 
    -116.158611, -116.2025, -116.2325, -116.241389, -116.261944, -116.278056, 
    -116.299722, -116.285833, -116.283333, -116.315833, -116.312222, 
    -116.298889, -116.283611, -116.273056, -116.248889, -116.240833, 
    -116.240833, -116.270278, -116.273611, -116.268611, -116.259444, -116.21, 
    -116.128333, -116.081667, -116.043611, -116.029444, -116.014167, 
    -115.984167, -115.952222, -115.933333, -115.913333, -115.83, -115.757778, 
    -115.738056, -115.7225, -115.713611, -115.720278, -115.729167, 
    -115.775833, NaN, -123.590111, -123.590389, -123.590389, -123.577556, 
    -123.559758451579, -123.543528, -123.506, -123.48675, -123.466806, 
    -123.439278, -123.412667, -123.408472, -123.401778, -123.379306, 
    -123.347667, -123.337222, -123.336778, -123.341778, -123.333444, 
    -123.326806, -123.328056, -123.323472, -123.313028, -123.318056, 
    -123.311333, -123.315194, -123.330056, -123.336833, -123.349306, 
    -123.352639, -123.357583, -123.386806, -123.393, -123.389667, 
    -123.400583, -123.390528, -123.393417, -123.400111, -123.406778, 
    -123.404694, -123.407639, -123.412194, -123.410167, -123.42675, 
    -123.490139, -123.50175, -123.50175, -123.523417, -123.542667, 
    -123.573472, -123.576333, -123.58475, -123.590111, NaN, -116.775278, 
    -116.779167, -116.802778, -116.813611, -116.791944, -116.780278, -116.78, 
    -116.783611, -116.804444, -116.846389, -116.848056, -116.841389, 
    -116.815833, -116.808056, -116.805278, -116.818056, -116.836111, 
    -116.919444, -116.926389, -116.918611, -116.896944, -116.886944, 
    -116.875833, -116.853333, -116.838333, -116.8125, -116.773333, -116.75, 
    -116.747222, -116.758889, -116.779444, -116.796944, -116.805833, 
    -116.809444, -116.818611, -116.83, -116.841389, -116.841944, -116.835556, 
    -116.800278, -116.773056, -116.770278, -116.779167, -116.766667, 
    -116.766111, -116.761667, -116.746111, -116.675833, -116.658333, 
    -116.654722, -116.723333, -116.775278, NaN, -122.527972, -122.527972, 
    -122.523806, -122.515444, -122.516306, -122.527972, -122.527972, 
    -122.514667, -122.512111, -122.512194, -122.495917, -122.482139, 
    -122.476306, -122.466722, -122.45125, -122.458833, -122.459611, 
    -122.448389, -122.441722, -122.432917, -122.442194, -122.438806, 
    -122.429611, -122.438028, -122.437083, -122.425028, -122.395861, 
    -122.372972, -122.400889, -122.422556, -122.431694, -122.443806, 
    -122.455028, -122.460917, -122.474639, -122.473833, -122.464194, 
    -122.455056, -122.432139, -122.439667, -122.440889, -122.463333, 
    -122.465861, -122.451694, -122.445444, -122.450889, -122.474167, 
    -122.484583, -122.493389, -122.51925, -122.527972, NaN, -118.547528, 
    -118.547, -118.544167, -118.521417, -118.493639, -118.459833, 
    -118.447806, -118.424306, -118.36625, -118.349389, -118.357417, 
    -118.363194, -118.393639, -118.402472, -118.405111, -118.415833, 
    -118.42525, -118.43075, -118.435222, -118.440083, -118.445667, 
    -118.451639, -118.477222, -118.490778, -118.49325, -118.501278, 
    -118.504389, -118.509972, -118.5095, -118.522194, -118.521167, 
    -118.533389, -118.540833, -118.54325, -118.548194, -118.545972, 
    -118.554194, -118.574917, -118.588806, -118.596722, -118.606278, 
    -118.607972, -118.595056, -118.586694, -118.574194, -118.565444, 
    -118.559611, -118.553361, -118.547972, -118.547528, NaN, -122.2025, 
    -122.2, -122.249722, -122.235278, -122.239167, -122.249167, -122.264444, 
    -122.270556, -122.271667, -122.265, -122.24, -122.234444, -122.236667, 
    -122.256389, -122.290556, -122.306944, -122.316389, -122.321667, 
    -122.317778, -122.308889, -122.300278, -122.288056, -122.270833, 
    -122.265, -122.260556, -122.263889, -122.253611, -122.237222, 
    -122.234722, -122.238333, -122.232778, -122.221111, -122.210556, 
    -122.197778, -122.185278, -122.192778, -122.183889, -122.178056, 
    -122.1925, -122.195, -122.219722, -122.223889, -122.2175, -122.196111, 
    -122.192778, -122.191667, -122.2025, NaN, -123.000528, -123, -123.017694, 
    -123.016722, -123.013056, -123.015083, -123.010111, -123.007639, 
    -123.006861, -122.982611, -122.970111, -122.971361, -122.967639, 
    -122.96675, -122.938444, -122.94475, -122.936, -122.930528, -122.933917, 
    -122.931389, -122.924333, -122.90925, -122.903833, -122.918444, 
    -122.925972, -122.92425, -122.936778, -122.940528, -122.93925, 
    -122.950944, -122.942194, -122.94675, -122.95175, -122.963472, 
    -122.968417, -122.971, -122.981028, -122.990528, -122.990528, 
    -122.985972, -122.97925, -122.973833, -122.982194, -122.982611, 
    -122.988472, -122.986306, -123.000528, NaN, -121.479722, -121.483611, 
    -121.488611, -121.525833, -121.539444, -121.544722, -121.548611, 
    -121.5575, -121.556111, -121.551667, -121.528611, -121.512778, 
    -121.504167, -121.494167, -121.480556, -121.476667, -121.479444, 
    -121.476111, -121.445556, -121.445278, -121.441944, -121.434722, 
    -121.420833, -121.413611, -121.370278, -121.354444, -121.347778, 
    -121.341111, -121.345556, -121.364722, -121.389722, -121.394167, 
    -121.394722, -121.387222, -121.357778, -121.361389, -121.3825, 
    -121.395278, -121.409167, -121.422778, -121.425278, -121.418056, 
    -121.4225, -121.449722, -121.459167, -121.479722, NaN, -115.964444, 
    -115.970278, -115.991944, -116.030833, -116.047222, -116.058611, 
    -116.062222, -116.044167, -116.037222, -116.029722, -116.022222, 
    -115.959444, -115.938333, -115.9225, -115.891389, -115.871667, 
    -115.862222, -115.855278, -115.836944, -115.822778, -115.808889, 
    -115.789722, -115.756111, -115.706111, -115.700833, -115.700278, 
    -115.695556, -115.683889, -115.68, -115.666389, -115.641667, -115.614722, 
    -115.61, -115.595, -115.593611, -115.606111, -115.636944, -115.648056, 
    -115.6625, -115.690833, -115.743889, -115.768611, -115.912222, 
    -115.934167, -115.964444, NaN, -119.923056, -119.924444, -119.923333, 
    -119.928056, -119.951667, -119.970833, -119.984444, -119.994444, 
    -120.008056, -120.027222, -120.047778, -120.075556, -120.088056, 
    -120.113889, -120.130833, -120.135, -120.150278, -120.151111, 
    -120.147222, -120.136111, -120.118333, -120.108889, -120.1075, 
    -120.086667, -120.090556, -120.0675, -120.049722, -120.030833, 
    -120.004444, -119.978889, -119.965278, -119.950278, -119.941389, 
    -119.940556, -119.932778, -119.936111, -119.930278, -119.942222, 
    -119.919167, -119.917778, -119.923056, NaN, -122.813333, -122.823056, 
    -122.845278, -122.876389, -122.88, -122.879722, -122.897778, -122.899722, 
    -122.894722, -122.885278, -122.821389, -122.775833, -122.759722, 
    -122.740833, -122.732778, -122.718333, -122.72, -122.716389, -122.691111, 
    -122.676111, -122.651389, -122.645278, -122.628333, -122.622222, 
    -122.616944, -122.615, -122.635833, -122.648889, -122.679444, -122.6975, 
    -122.661389, -122.649444, -122.644722, -122.649167, -122.706111, 
    -122.731389, -122.756944, -122.769722, -122.785278, -122.796667, 
    -122.813333, NaN, -119.042222, -119.0425, -119.043056, -119.048056, 
    -119.069722, -119.100556, -119.115833, -119.145833, -119.161944, 
    -119.179444, -119.188611, -119.191389, -119.186944, -119.181667, 
    -119.142778, -119.133611, -119.128889, -119.139444, -119.124444, 
    -119.1125, -119.114444, -119.111389, -119.100556, -119.067222, 
    -119.063611, -119.066111, -119.085, -119.124722, -119.165556, 
    -119.169167, -119.161389, -119.137778, -119.104722, -119.088611, 
    -119.083889, -119.078889, -119.071944, -119.066389, -119.045278, 
    -119.042222, NaN, -120.364167, -120.365278, -120.37375, -120.383222, 
    -120.40875, -120.414944, -120.417667, -120.428278, -120.4395, 
    -120.449694, -120.452639, -120.448139, -120.449111, -120.438444, 
    -120.430333, -120.417917, -120.418333, -120.414778, -120.411556, 
    -120.402444, -120.389917, -120.372556, -120.367028, -120.369944, 
    -120.367639, -120.361444, -120.3565, -120.354278, -120.359222, 
    -120.355167, -120.340528, -120.331583, -120.317611, -120.306417, 
    -120.294, -120.294917, -120.314667, -120.349194, -120.356917, 
    -120.364167, NaN, -119.327222, -119.331667, -119.335833, -119.341389, 
    -119.353889, -119.356111, -119.341944, -119.347778, -119.355, 
    -119.363889, -119.398889, -119.411667, -119.420556, -119.425833, 
    -119.435278, -119.43, -119.420556, -119.420278, -119.429722, -119.428333, 
    -119.402222, -119.355278, -119.335556, -119.314167, -119.305, 
    -119.298056, -119.278611, -119.270556, -119.246111, -119.183056, 
    -119.158889, -119.147222, -119.147778, -119.155556, -119.201389, 
    -119.240833, -119.275278, -119.292222, -119.308889, -119.327222, NaN, 
    -121.064167, -121.063056, -121.080556, -121.093889, -121.1125, 
    -121.117778, -121.110833, -121.081944, -121.068611, -121.044722, 
    -121.017222, -121.003333, -121.005, -121.023611, -121.025278, 
    -121.023056, -121, -121.000556, -121.0225, -121.034444, -121.036389, 
    -121.056111, -121.058611, -121.056512774235, -121.068333, 
    -121.083374538379, -121.083611, -121.065833, -121.062222, -121.056389, 
    -121.023056, -121.021944, -121.0475, -121.054167, -121.047222, 
    -121.029722, -121.028056, -121.035833, -121.064167, NaN, -122.750583, 
    -122.750583, -122.737639, -122.725944, -122.726333, -122.718028, 
    -122.720528, -122.713083, -122.715556, -122.706361, -122.701, 
    -122.693056, -122.703861, -122.705528, -122.699306, -122.694278, 
    -122.693444, -122.693056, -122.702167, -122.705583, -122.718028, 
    -122.730556, -122.705972, -122.690111, -122.693056, -122.686389, 
    -122.684778, -122.681833, -122.668833, -122.671389, -122.683444, 
    -122.691806, -122.696833, -122.725083, -122.733222, -122.743861, 
    -122.740528, -122.750583, NaN, -123.328806, -123.328806, -123.327639, 
    -123.320528, -123.319694, -123.328944, -123.32425, -123.308417, 
    -123.301722, -123.291833, -123.285167, -123.277194, -123.27675, 
    -123.271861, -123.255944, -123.249667, -123.239694, -123.257639, 
    -123.274278, -123.274278, -123.258056, -123.268083, -123.256, 
    -123.241806, -123.240139, -123.231333, -123.232611, -123.256806, 
    -123.308444, -123.315111, -123.313028, -123.321389, -123.309722, 
    -123.318889, -123.31225, -123.315111, -123.305528, -123.328806, NaN, 
    -124.329444, -124.331111, -124.3475, -124.376667, -124.418889, 
    -124.448333, -124.450556, -124.433333, -124.413333, -124.396667, -124.38, 
    -124.3575, -124.349722, -124.348889, -124.339167, -124.288056, 
    -124.248333, -124.217778, -124.198333, -124.165278, -124.146944, 
    -124.093611, -124.070556, -124.052222, -124.057778, -124.105, -124.13, 
    -124.136389, -124.131944, -124.140278, -124.199722, -124.214444, 
    -124.238889, -124.256389, -124.273611, -124.284167, -124.329444, NaN, 
    -118.549444, -118.556667, -118.571111, -118.588056, -118.590833, 
    -118.566944, -118.535278, -118.511111, -118.472222, -118.453056, 
    -118.435278, -118.429167, -118.428889, -118.432778, -118.450833, 
    -118.475, -118.495278, -118.500833, -118.495833, -118.489444, 
    -118.463889, -118.441389, -118.436944, -118.435833, -118.43, -118.419444, 
    -118.422778, -118.42, -118.406944, -118.401389, -118.409444, -118.385833, 
    -118.3875, -118.401389, -118.445278, -118.469444, -118.549444, NaN, 
    -120.386111, -120.391667, -120.424722, -120.441944, -120.480833, 
    -120.501667, -120.499722, -120.484444, -120.478611, -120.490833, 
    -120.481944, -120.483333, -120.502778, -120.494167, -120.471944, 
    -120.4725, -120.459722, -120.4625, -120.471667, -120.476389, -120.477222, 
    -120.471944, -120.402222, -120.372222, -120.368611, -120.370833, 
    -120.358333, -120.356389, -120.346111, -120.326667, -120.321389, 
    -120.320278, -120.312778, -120.315556, -120.336389, -120.359167, 
    -120.386111, NaN, -119.497778, -119.500278, -119.507222, -119.5175, 
    -119.585, -119.598056, -119.648611, -119.658611, -119.664722, 
    -119.691389, -119.695, -119.681389, -119.671944, -119.629444, -119.6125, 
    -119.605556, -119.597778, -119.574167, -119.563056, -119.522222, 
    -119.468611, -119.454722, -119.4425, -119.434444, -119.424722, 
    -119.401111, -119.411944, -119.450278, -119.463889, -119.481667, 
    -119.485278, -119.484167, -119.478889, -119.475833, -119.486944, 
    -119.497778, NaN, -120.213056, -120.219722, -120.226667, -120.243889, 
    -120.328333, -120.367778, -120.414167, -120.443889, -120.441111, 
    -120.4075, -120.349444, -120.326667, -120.285278, -120.260556, 
    -120.245278, -120.239722, -120.232778, -120.230278, -120.2325, 
    -120.241944, -120.273889, -120.295278, -120.306667, -120.308611, 
    -120.303889, -120.287222, -120.280833, -120.199167, -120.163889, 
    -120.155833, -120.151944, -120.157222, -120.18, -120.187778, -120.213056, 
    NaN, -114.700083, -114.701361, -114.711528, -114.716056, -114.714139, 
    -114.753611, -114.772722, -114.792611, -114.800306, -114.801083, 
    -114.795833, -114.795861, -114.764917, -114.747778, -114.728556, 
    -114.709667, -114.71125, -114.705972, -114.655806, -114.641722, 
    -114.640722, -114.643389, -114.640611, -114.643194, -114.657, -114.662, 
    -114.676222, -114.683056, -114.687861, -114.681806, -114.688222, 
    -114.692639, -114.690083, -114.688639, -114.700083, NaN, -118.088611, 
    -118.086667, -118.093333, -118.111944, -118.118611, -118.117778, 
    -118.151389, -118.168889, -118.205556, -118.215, -118.221667, 
    -118.226944, -118.191667, -118.187778, -118.163056, -118.149444, 
    -118.142778, -118.163611, -118.170833, -118.187778, -118.193056, 
    -118.203889, -118.202222, -118.198611, -118.155556, -118.149444, 
    -118.123889, -118.124722, -118.115, -118.094444, -118.083333, 
    -118.083889, -118.069444, -118.088611, NaN, -120.664444, -120.663333, 
    -120.669167, -120.678889, -120.705556, -120.716389, -120.720278, 
    -120.727222, -120.739167, -120.759722, -120.765278, -120.766944, 
    -120.755, -120.764444, -120.804444, -120.8025, -120.792778, -120.7775, 
    -120.767222, -120.727222, -120.721111, -120.721944, -120.703333, 
    -120.696667, -120.698611, -120.692222, -120.685, -120.667778, 
    -120.659722, -120.654722, -120.651389, -120.6525, -120.657778, 
    -120.664444, NaN, -114.354722, -114.356389, -114.375833, -114.373889, 
    -114.391667, -114.398056, -114.396389, -114.387778, -114.365833, 
    -114.335278, -114.324444, -114.304167, -114.295833, -114.285833, 
    -114.171667, -114.135, -114.113056, -114.065, -114.062778, -114.073889, 
    -114.096944, -114.123611, -114.139167, -114.1675, -114.200833, 
    -114.218056, -114.276111, -114.290833, -114.312222, -114.3325, -114.34, 
    -114.35, -114.355556, -114.354722, NaN, -124.000472, -124, -123.992556, 
    -123.992167, -123.986667, -123.979972, -123.971222, -123.976694, 
    -123.985056, -123.987917, -123.978778, -123.978389, -123.975417, 
    -123.974611, -123.970889, -123.966278, -123.970028, -123.962556, 
    -123.942889, -123.942111, -123.947917, -123.945472, -123.935472, 
    -123.940833, -123.965889, -123.971361, -123.965472, -123.968806, 
    -123.991694, -123.995028, -124.003, -124.004472, -124.000472, NaN, 
    -123.347167, -123.346833, -123.324306, -123.314333, -123.302639, 
    -123.299639, -123.307222, -123.292667, -123.28675, -123.277611, 
    -123.258472, -123.245528, -123.246806, -123.261722, -123.27225, 
    -123.244722, -123.24975, -123.246361, -123.254778, -123.231806, 
    -123.228028, -123.238444, -123.242583, -123.250139, -123.276778, 
    -123.281778, -123.3285, -123.3285, -123.321333, -123.334694, -123.323028, 
    -123.347167, NaN, -121.055833, -121.057222, -121.060833, -121.069722, 
    -121.082222, -121.099167, -121.131389, -121.151111, -121.168056, 
    -121.209444, -121.214167, -121.208611, -121.207222, -121.211111, 
    -121.191667, -121.165278, -121.149444, -121.14, -121.134444, -121.113333, 
    -121.105556, -121.129167, -121.131389, -121.126389, -121.101111, 
    -121.087778, -121.068056, -121.061667, -121.055, -121.050833, 
    -121.051111, -121.055833, NaN, -114.905833, -114.899314, -114.890833, 
    -114.874722, -114.845556, -114.827222, -114.824722, -114.82, -114.793889, 
    -114.718889, -114.692778, -114.674722, -114.671389, -114.6725, 
    -114.658333, -114.656667, -114.659722, -114.676111, -114.697222, 
    -114.721667, -114.731111, -114.741667, -114.769722, -114.774444, 
    -114.810556, -114.821667, -114.834722, -114.854722, -114.864444, 
    -114.878056, -114.885278, -114.905833, NaN, -122.245, -122.249444, 
    -122.260278, -122.264444, -122.271667, -122.275278, -122.278611, 
    -122.285278, -122.281389, -122.293056, -122.258333, -122.246389, 
    -122.236944, -122.220833, -122.209444, -122.187778, -122.192222, 
    -122.186667, -122.175833, -122.169722, -122.1575, -122.151389, 
    -122.143056, -122.120556, -122.1125, -122.105278, -122.109444, 
    -122.163889, -122.184167, -122.212778, -122.231667, -122.245, NaN, 
    -118.731111, -118.738333, -118.753611, -118.755833, -118.762778, 
    -118.785, -118.806944, -118.853611, -118.886667, -118.953056, 
    -118.958056, -118.96, -118.948056, -118.938611, -118.854167, -118.833889, 
    -118.815278, -118.800833, -118.783056, -118.769444, -118.761944, 
    -118.749444, -118.740833, -118.729444, -118.706667, -118.668333, 
    -118.660833, -118.660833, -118.682778, -118.689167, -118.731111, NaN, 
    -119.486361, -119.485528, -119.4605, -119.429944, -119.437472, 
    -119.439222, -119.451722, -119.459667, -119.476806, -119.484611, 
    -119.499583, -119.515028, -119.520722, -119.534083, -119.546917, 
    -119.567028, -119.566583, -119.575611, -119.574694, -119.580167, 
    -119.573278, -119.561611, -119.556861, -119.551889, -119.540111, 
    -119.535861, -119.528306, -119.499278, -119.487472, -119.486361, NaN, 
    -118.259722, -118.262222, -118.267222, -118.282222, -118.293889, 
    -118.311111, -118.32, -118.335, -118.339167, -118.338333, -118.329167, 
    -118.31, -118.302222, -118.307778, -118.304167, -118.282778, -118.290833, 
    -118.3175, -118.326667, -118.311389, -118.303889, -118.280556, 
    -118.274167, -118.234722, -118.220556, -118.2175, -118.233889, 
    -118.251389, -118.259722, NaN, -123.215556, -123.215472, -123.211778, 
    -123.2035, -123.200083, -123.197222, -123.20175, -123.178389, 
    -123.203861, -123.203444, -123.195139, -123.186778, -123.127556, 
    -123.110972, -123.100139, -123.044722, -123.047694, -123.061, 
    -123.112639, -123.093444, -123.089722, -123.094306, -123.131806, 
    -123.132556, -123.142611, -123.159278, -123.2035, -123.202972, 
    -123.215556, NaN, -114.638333, -114.638333, -114.643889, -114.641389, 
    -114.646944, -114.665278, -114.655833, -114.655, -114.676389, 
    -114.678889, -114.678889, -114.666667, -114.669444, -114.658889, 
    -114.615833, -114.594444, -114.590556, -114.583056, -114.579722, 
    -114.594722, -114.597778, -114.607778, -114.646389, -114.653889, 
    -114.6525, -114.635, -114.632778, -114.638333, NaN, -125.122111, 
    -125.121667, -125.109583, -125.108806, -125.113722, -125.109278, 
    -125.103778, -125.109583, -125.097889, -125.099222, -125.086694, 
    -125.090389, -125.082583, -125.071667, -125.068389, -125.051667, 
    -125.047167, -125.057944, -125.058833, -125.068306, -125.081667, 
    -125.086694, -125.101694, -125.105861, -125.114222, -125.122111, NaN, 
    -122.74225, -122.742194, -122.730556, -122.731417, -122.720889, 
    -122.712611, -122.706778, -122.705111, -122.695556, -122.693, -122.7005, 
    -122.668861, -122.672611, -122.676806, -122.698083, -122.697639, 
    -122.691806, -122.684306, -122.685111, -122.723528, -122.725611, 
    -122.722194, -122.740556, -122.74225, NaN, -121.084444, -121.085833, 
    -121.095556, -121.110278, -121.119444, -121.125556, -121.128056, 
    -121.125278, -121.131667, -121.163611, -121.171667, -121.181389, 
    -121.189444, -121.196389, -121.205833, -121.204444, -121.189722, -121.16, 
    -121.112222, -121.085, -121.073889, -121.069722, -121.0725, -121.084444, 
    NaN, -121.116389, -121.125556, -121.134722, -121.149167, -121.174167, 
    -121.174444, -121.161111, -121.146944, -121.138611, -121.1325, 
    -121.135833, -121.128889, -121.118333, -121.111944, -121.113889, 
    -121.111111, -121.093611, -121.075556, -121.067778, -121.064167, 
    -121.070833, -121.080556, -121.109167, -121.116389, NaN, -122.724722, 
    -122.724694, -122.7185, -122.705111, -122.695917, -122.690917, 
    -122.683028, -122.670917, -122.665194, -122.662583, -122.659333, 
    -122.646861, -122.635111, -122.628444, -122.625056, -122.618861, 
    -122.609278, -122.622667, -122.636806, -122.676028, -122.690583, 
    -122.705111, -122.720139, -122.724722, NaN, -118.7225, -118.729722, 
    -118.746389, -118.752222, -118.738889, -118.738056, -118.756667, 
    -118.756944, -118.748056, -118.753889, -118.745833, -118.733056, 
    -118.697778, -118.684722, -118.670833, -118.656111, -118.646944, 
    -118.646389, -118.660278, -118.659722, -118.663333, -118.706389, 
    -118.7225, NaN, -122.922167, -122.92225, -122.916361, -122.917556, 
    -122.92225, -122.920139, -122.906833, -122.878861, -122.885972, 
    -122.910167, -122.913111, -122.902667, -122.898417, -122.891, 
    -122.885972, -122.894278, -122.902667, -122.908861, -122.898417, 
    -122.915194, -122.915972, -122.911361, -122.922167, NaN, -123.347222, 
    -123.347278, -123.321, -123.305972, -123.292611, -123.271778, 
    -123.268861, -123.270944, -123.285944, -123.295111, -123.298861, 
    -123.310528, -123.315194, -123.338, -123.342194, -123.340167, -123.33475, 
    -123.337222, -123.331778, -123.328028, -123.328806, -123.332278, 
    -123.347222, NaN, -125.278778, -125.278361, -125.26675, -125.270028, 
    -125.262583, -125.250861, -125.239222, -125.235861, -125.23675, 
    -125.2275, -125.227111, -125.241694, -125.240917, -125.246722, 
    -125.250917, -125.255889, -125.261667, -125.250389, -125.258361, 
    -125.271722, -125.272111, -125.278778, NaN, -122.841417, -122.841361, 
    -122.838472, -122.833056, -122.830972, -122.818444, -122.789306, 
    -122.790194, -122.79725, -122.796389, -122.791, -122.7885, -122.783861, 
    -122.798472, -122.8185, -122.818444, -122.821778, -122.827194, 
    -122.817194, -122.818889, -122.83175, -122.841417, NaN, -120.148333, 
    -120.146389, -120.138611, -120.139167, -120.148056, -120.232778, 
    -120.240278, -120.244167, -120.248611, -120.270278, -120.278333, 
    -120.275278, -120.268889, -120.2525, -120.246944, -120.245278, 
    -120.238889, -120.2225, -120.179167, -120.175833, -120.163333, 
    -120.148333, NaN, -123.239694, -123.239694, -123.237556, -123.211778, 
    -123.205583, -123.205972, -123.210528, -123.207667, -123.185167, 
    -123.179278, -123.175139, -123.164694, -123.170556, -123.16725, 
    -123.173472, -123.176833, -123.205917, -123.182611, -123.182222, 
    -123.187667, -123.21675, -123.239694, NaN, -123.204722, -123.204722, 
    -123.198083, -123.189333, -123.180889, -123.174667, -123.183, 
    -123.178889, -123.180056, -123.187194, -123.185111, -123.179278, 
    -123.171333, -123.181306, -123.178111, -123.183528, -123.186389, 
    -123.186778, -123.191417, -123.196778, -123.204722, NaN, -121.734167, 
    -121.740556, -121.751667, -121.758333, -121.764167, -121.774167, -121.8, 
    -121.803056, -121.800556, -121.786389, -121.741944, -121.721389, 
    -121.694167, -121.679167, -121.671111, -121.671111, -121.662222, 
    -121.668889, -121.678056, -121.723889, -121.734167, NaN, -121.084444, 
    -121.086111, -121.078889, -121.085, -121.100556, -121.101667, 
    -121.110278, -121.162778, -121.16, -121.130833, -121.122778, -121.094444, 
    -121.082778, -121.055278, -121.053056, -121.057222, -121.0975, 
    -121.106389, -121.108889, -121.086111, -121.084444, NaN, -119.133056, 
    -119.139722, -119.166944, -119.194167, -119.206389, -119.207222, 
    -119.194722, -119.158056, -119.142222, -119.119167, -119.099722, 
    -119.082778, -119.0675, -119.054167, -119.035, -119.0425, -119.054722, 
    -119.075, -119.124444, -119.133056, NaN, -123.677111, -123.677111, 
    -123.661722, -123.666306, -123.661722, -123.643389, -123.644222, 
    -123.6505, -123.645028, -123.633333, -123.635833, -123.628778, 
    -123.634639, -123.634583, -123.649222, -123.660083, -123.660861, 
    -123.667528, -123.677111, NaN, -123.409639, -123.409333, -123.397167, 
    -123.405528, -123.403472, -123.363444, -123.355167, -123.352167, 
    -123.355167, -123.365528, -123.359667, -123.360889, -123.377222, 
    -123.365111, -123.365167, -123.383444, -123.405528, -123.395556, 
    -123.409639, NaN, -123.671389, -123.671389, -123.669333, -123.662639, 
    -123.661806, -123.644278, -123.640556, -123.642611, -123.636333, 
    -123.638, -123.629694, -123.631778, -123.639306, -123.639306, 
    -123.652583, -123.658028, -123.663028, -123.658944, -123.671389, NaN, 
    -118.944722, -118.952222, -118.996667, -119.021667, -119.052778, 
    -119.037222, -119.01, -118.992778, -118.983056, -118.949722, -118.937778, 
    -118.930556, -118.926111, -118.917222, -118.8775, -118.875833, 
    -118.896111, -118.906389, -118.944722, NaN, -116.085556, -116.089444, 
    -116.101389, -116.106667, -116.092778, -116.093056, -116.095, 
    -116.111111, -116.12, -116.125, -116.122778, -116.086944, -116.061944, 
    -116.046944, -116.043611, -116.050278, -116.054722, -116.080556, 
    -116.085556, NaN, -122.655556, -122.655528, -122.653833, -122.64725, 
    -122.653861, -122.653, -122.645167, -122.630111, -122.611778, 
    -122.581806, -122.573917, -122.590167, -122.59175, -122.603556, 
    -122.628444, -122.640944, -122.653472, -122.655556, NaN, -116.041389, 
    -116.042778, -116.045278, -116.053889, -116.066111, -116.080278, 
    -116.089167, -116.112778, -116.104167, -116.097778, -116.079167, 
    -116.065833, -116.058056, -116.054722, -116.046111, -116.042778, 
    -116.045, -116.041389, NaN, -120.750833, -120.753333, -120.7575, 
    -120.763056, -120.769722, -120.7975, -120.790278, -120.789167, 
    -120.778611, -120.761389, -120.728889, -120.712778, -120.696111, 
    -120.698333, -120.7175, -120.742222, -120.750833, NaN, -122.833083, 
    -122.833083, -122.826861, -122.816806, -122.816806, -122.811861, 
    -122.793444, -122.770556, -122.780083, -122.795944, -122.800167, 
    -122.804361, -122.811806, -122.824778, -122.818056, -122.828111, 
    -122.833083, NaN, -118.734167, -118.736389, -118.741667, -118.7525, 
    -118.742222, -118.744444, -118.760833, -118.772222, -118.770833, 
    -118.757778, -118.738333, -118.722778, -118.712778, -118.720833, -118.72, 
    -118.734167, NaN, -123.072167, -123.072167, -123.051722, -123.042583, 
    -123.027583, -123.025056, -123.012667, -123.009722, -123.008944, 
    -123.004694, -123.012194, -123.005556, -123.017611, -123.044306, 
    -123.040056, -123.072167, NaN, -122.653, -122.653, -122.645167, 
    -122.6335, -122.626056, -122.620139, -122.618, -122.629722, -122.623417, 
    -122.612222, -122.607222, -122.608833, -122.615944, -122.625083, 
    -122.635917, -122.653, NaN, -125.294611, -125.294694, -125.293361, 
    -125.289194, -125.281722, -125.274194, -125.264583, -125.276667, 
    -125.277528, -125.282556, -125.292583, -125.290833, -125.277083, 
    -125.291667, -125.290417, -125.294611, NaN, -122.849167, -122.849167, 
    -122.842778, -122.845556, -122.868056, -122.896111, -122.902222, 
    -122.912222, -122.911389, -122.869722, -122.859444, -122.829444, 
    -122.831944, -122.851389, -122.858889, -122.849167, NaN, -123.703056, 
    -123.702944, -123.702944, -123.702472, -123.695861, -123.6875, 
    -123.689639, -123.685861, -123.659095260324, -123.653, -123.674722, 
    -123.669333, -123.675944, -123.680139, -123.691806, -123.703056, NaN, 
    -122.080556, -122.089167, -122.125, -122.148056, -122.159167, -122.155, 
    -122.145833, -122.133056, -122.098333, -122.0775, -122.066944, 
    -122.053056, -122.05, -122.064722, -122.080556, NaN, -123.258056, 
    -123.258056, -123.250139, -123.235056, -123.204278, -123.173806, 
    -123.187639, -123.183056, -123.186722, -123.208472, -123.216806, 
    -123.231028, -123.234222, -123.2485, -123.258056, NaN, -118.613889, 
    -118.611667, -118.606111, -118.603889, -118.619167, -118.64, -118.651111, 
    -118.658611, -118.655, -118.649722, -118.642222, -118.641667, 
    -118.637222, -118.63, -118.613889, NaN, -119.3845, -119.384167, 
    -119.380806, -119.389417, -119.402389, -119.410194, -119.420222, 
    -119.425694, -119.427361, -119.446028, -119.424139, -119.409028, 
    -119.392917, -119.3845, NaN, -122.6675, -122.668333, -122.681944, 
    -122.698056, -122.708889, -122.726111, -122.723611, -122.699167, 
    -122.690278, -122.685, -122.681944, -122.683333, -122.665278, -122.6675, 
    NaN, -125.163806, -125.163806, -125.158333, -125.143389, -125.142917, 
    -125.133417, -125.123361, -125.120028, -125.115472, -125.1325, 
    -125.140917, -125.15175, -125.163806, NaN, -123.721278, -123.721278, 
    -123.704222, -123.697528, -123.692111, -123.693389, -123.687556, 
    -123.68625, -123.695917, -123.684139, -123.674583, -123.697528, 
    -123.721278, NaN, -125.363833, -125.36375, -125.358333, -125.35675, 
    -125.350833, -125.35, -125.337917, -125.340028, -125.348389, -125.348361, 
    -125.355889, -125.356639, -125.363833, NaN, -119.597778, -119.596944, 
    -119.595556, -119.61, -119.636389, -119.69, -119.695833, -119.686667, 
    -119.665833, -119.644167, -119.630833, -119.612778, -119.597778, NaN, 
    -123.736278, -123.736306, -123.732528, -123.718806, -123.724556, 
    -123.723361, -123.726722, -123.726694, -123.730861, -123.734583, 
    -123.726306, -123.730889, -123.736278, NaN, -118.600278, -118.597778, 
    -118.595556, -118.600833, -118.628056, -118.622222, -118.625556, 
    -118.618056, -118.596944, -118.593056, -118.591667, -118.600278, NaN, 
    -123.333861, -123.333889, -123.327194, -123.330972, -123.310111, 
    -123.305583, -123.291361, -123.296389, -123.302194, -123.29925, 
    -123.319278, -123.333861, NaN, -115.599, -115.599194, -115.598, 
    -115.582917, -115.577333, -115.571306, -115.568361, -115.572528, 
    -115.569139, -115.570917, -115.586306, -115.599, NaN, -122.447139, 
    -122.447139, -122.442111, -122.440028, -122.435861, -122.433389, 
    -122.428361, -122.422083, -122.419611, -122.430833, -122.435861, 
    -122.447139, NaN, -116.9225, -116.924167, -116.930833, -116.937222, 
    -116.930278, -116.935833, -116.932222, -116.922778, -116.902778, 
    -116.909722, -116.915833, -116.9225, NaN, -114.139222, -114.138611, 
    -114.130056, -114.116306, -114.117472, -114.124222, -114.130639, 
    -114.138, -114.141917, -114.145083, -114.146917, -114.139222, NaN, 
    -123.379639, -123.378444, -123.358444, -123.348472, -123.335528, 
    -123.336833, -123.350917, -123.358028, -123.356028, -123.353083, 
    -123.357583, -123.379639, NaN, -120.129722, -120.134444, -120.166667, 
    -120.176389, -120.155278, -120.12, -120.113611, -120.091944, -120.095556, 
    -120.101944, -120.108889, -120.129722, NaN, -122.641667, -122.6375, 
    -122.633333, -122.636111, -122.6625, -122.682222, -122.696389, 
    -122.712222, -122.708333, -122.668889, -122.652778, -122.641667, NaN, 
    -114.604917, -114.607, -114.630667, -114.65475, -114.666333, -114.6715, 
    -114.660611, -114.606611, -114.596472, -114.594889, -114.599222, 
    -114.604917, NaN, -123.939667, -123.942222, -123.949167, -123.950472, 
    -123.956806, -123.956028, -123.951556, -123.942056, -123.936, 
    -123.940722, -123.939667, NaN, -116.9225, -116.924444, -116.933889, 
    -116.933889, -116.929167, -116.909167, -116.893056, -116.894167, 
    -116.898889, -116.913611, -116.9225, NaN, -114.064556, -114.064944, 
    -114.068444, -114.071028, -114.079972, -114.071, -114.055972, 
    -114.059167, -114.057944, -114.060583, -114.064556, NaN, -123.330833, 
    -123.326944, -123.322778, -123.344167, -123.354722, -123.401667, 
    -123.411389, -123.411667, -123.4, -123.3475, -123.330833, NaN, 
    -125.336333, -125.336306, -125.331278, -125.331722, -125.326667, 
    -125.317583, -125.312111, -125.328361, -125.329194, -125.335056, 
    -125.336333, NaN, -123.234667, -123.234694, -123.221833, -123.188861, 
    -123.204333, -123.210556, -123.205583, -123.210917, -123.222611, 
    -123.224333, -123.234667, NaN, -114.385778, -114.3845, -114.381639, 
    -114.370583, -114.381083, -114.392083, -114.396167, -114.40225, 
    -114.399194, -114.390917, -114.385778, NaN, -114.421444, -114.421389, 
    -114.417917, -114.419, -114.432722, -114.446, -114.4475, -114.440889, 
    -114.441972, -114.426333, -114.421444, NaN, -122.195278, -122.193611, 
    -122.191944, -122.198611, -122.207222, -122.217222, -122.22, -122.234722, 
    -122.219722, -122.202778, -122.195278, NaN, -122.610278, -122.616389, 
    -122.643889, -122.652778, -122.651944, -122.618333, -122.602778, 
    -122.594722, -122.586389, -122.586944, -122.610278, NaN, -125.350444, 
    -125.350417, -125.340472, -125.344194, -125.3275, -125.323722, 
    -125.33175, -125.333361, -125.343333, -125.350444, NaN, -116.128806, 
    -116.128778, -116.120889, -116.115, -116.110472, -116.104583, 
    -116.113333, -116.117556, -116.126639, -116.128806, NaN, -123.388056, 
    -123.387972, -123.376833, -123.375972, -123.374306, -123.365139, 
    -123.360528, -123.372194, -123.371722, -123.388056, NaN, -114.55575, 
    -114.556111, -114.54175, -114.535722, -114.537472, -114.544444, 
    -114.548222, -114.551306, -114.555944, -114.55575, NaN, -125.22625, 
    -125.226306, -125.214194, -125.205028, -125.2025, -125.197083, 
    -125.212611, -125.215, -125.223389, -125.22625, NaN, -124.164444, 
    -124.165278, -124.168889, -124.195833, -124.197778, -124.190833, 
    -124.184444, -124.176944, -124.163889, -124.164444, NaN, -118.218889, 
    -118.221389, -118.231111, -118.241944, -118.245, -118.244444, -118.2325, 
    -118.217778, -118.211111, -118.218889, NaN, -122.379694, -122.379694, 
    -122.375861, -122.366306, -122.362917, -122.3705, -122.362917, 
    -122.363389, -122.372972, -122.379694, NaN, -124.010278, -124.006944, 
    -124.003139, -124.006472, -124.027278, -124.031694, -124.033611, 
    -124.025972, -124.023111, -124.010278, NaN, -123.103861, -123.103861, 
    -123.075944, -123.076722, -123.0635, -123.061778, -123.051417, 
    -123.060111, -123.071778, -123.103861, NaN, -123.628806, -123.628722, 
    -123.625056, -123.617556, -123.609972, -123.598389, -123.590472, 
    -123.589639, -123.595917, -123.628806, NaN, -123.5255, -123.5255, 
    -123.508333, -123.503778, -123.504194, -123.4905, -123.491694, 
    -123.510028, -123.514222, -123.5255, NaN, -125.320444, -125.320444, 
    -125.308389, -125.307083, -125.312083, -125.302583, -125.291278, 
    -125.314167, -125.320444, NaN, -114.131278, -114.131389, -114.129778, 
    -114.117639, -114.118194, -114.125444, -114.116056, -114.126139, 
    -114.131278, NaN, -122.899444, -122.900556, -122.908333, -122.916111, 
    -122.908889, -122.898333, -122.891389, -122.891944, -122.899444, NaN, 
    -125.265472, -125.265444, -125.260833, -125.24375, -125.253389, 
    -125.255861, -125.260889, -125.261278, -125.265472, NaN, -123.165528, 
    -123.165528, -123.15925, -123.150111, -123.149306, -123.141833, 
    -123.136361, -123.145083, -123.165528, NaN, -119.030778, -119.030556, 
    -119.032972, -119.041861, -119.048444, -119.039361, -119.031528, 
    -119.028639, -119.030778, NaN, -122.335528, -122.335528, -122.330972, 
    -122.324306, -122.311806, -122.303889, -122.310917, -122.327639, 
    -122.335528, NaN, -123.556278, -123.556278, -123.545861, -123.539194, 
    -123.530028, -123.52875, -123.538306, -123.5475, -123.556278, NaN, 
    -123.622139, -123.622194, -123.596694, -123.572472, -123.567194, 
    -123.568361, -123.584139, -123.604194, -123.622139, NaN, -123.500444, 
    -123.500444, -123.479167, -123.453806, -123.470056, -123.480861, 
    -123.487944, -123.495889, -123.500444, NaN, -122.505472, -122.505472, 
    -122.495889, -122.480028, -122.478778, -122.4855, -122.484194, 
    -122.495917, -122.505472, NaN, -122.701361, -122.701361, -122.675972, 
    -122.663889, -122.659722, -122.669306, -122.679278, -122.700083, 
    -122.701361, NaN, -125.335444, -125.335444, -125.332194, -125.337556, 
    -125.348389, -125.351306, -125.34986117776, -125.335373044127, 
    -125.335444, NaN, -123.630111, -123.631972, -123.631972, -123.626667, 
    -123.618122656598, -123.614694, -123.619278, -123.623417, -123.630111, 
    NaN, -125.208833, -125.208833, -125.203333, -125.201722, -125.185, 
    -125.190028, -125.2055, -125.204139, -125.208833, NaN, -123.055528, 
    -123.055528, -123.050111, -123.046722, -123.043444, -123.038028, 
    -123.050111, -123.055528, NaN, -123.627917, -123.627917, -123.615861, 
    -123.606278, -123.618389, -123.624667, -123.6225, -123.627917, NaN, 
    -123.167222, -123.165111, -123.120972, -123.115944, -123.107583, 
    -123.108028, -123.132583, -123.167222, NaN, -122.5955, -122.595139, 
    -122.588, -122.587639, -122.579722, -122.582611, -122.584278, -122.5955, 
    NaN, -124.136833, -124.13925, -124.148417, -124.149111, -124.139444, 
    -124.125361, -124.130083, -124.136833, NaN, -125.327167, -125.327083, 
    -125.322528, -125.316722, -125.318361, -125.311278, -125.314972, 
    -125.327167, NaN, -123.479639, -123.479639, -123.456667, -123.440889, 
    -123.435472, -123.439167, -123.473361, -123.479639, NaN, -125.353806, 
    -125.353778, -125.345889, -125.334167, -125.330028, -125.339167, 
    -125.339167, -125.353806, NaN, -123.388833, -123.388861, -123.38475, 
    -123.38675, -123.364694, -123.3735, -123.385111, -123.388833, NaN, 
    -123.574694, -123.574694, -123.552639, -123.535944, -123.535944, 
    -123.557611, -123.558444, -123.574694, NaN, -122.824778, -122.824778, 
    -122.819667, -122.816806, -122.806389, -122.811861, -122.822611, 
    -122.824778, NaN, -123.251361, -123.251361, -123.245972, -123.229333, 
    -123.225528, -123.233417, -123.243417, -123.251361, NaN, -122.001944, 
    -122.008889, -122.018056, -121.998333, -121.992222, -121.986111, 
    -121.983333, -122.001944, NaN, -115.566417, -115.566417, -115.566722, 
    -115.559917, -115.553139, -115.554861, -115.562056, -115.566417, NaN, 
    -123.435556, -123.435556, -123.420139, -123.411806, -123.397194, 
    -123.396861, -123.41675, -123.435556, NaN, -122.945556, -122.943444, 
    -122.934306, -122.924333, -122.910556, -122.92425, -122.935167, 
    -122.945556, NaN, -123, -123.001306, -123.004778, -123.003917, 
    -123.009722, -123.005, -123.001389, -123, NaN, -123.201389, -123.201389, 
    -123.184722, -123.188861, -123.187556, -123.196833, -123.196833, 
    -123.201389, NaN, -123.000972, -123, -122.994333, -122.989333, 
    -122.995111, -123.006861, -123.008889, -123.000972, NaN, -125.369556, 
    -125.36925, -125.35425, -125.351306, -125.360056, -125.362528, 
    -125.369556, NaN, -121.832778, -121.836944, -121.851944, -121.855, 
    -121.829722, -121.826111, -121.832778, NaN, -115.799194, -115.799167, 
    -115.796778, -115.792583, -115.795139, -115.798639, -115.799194, NaN, 
    -121.811389, -121.82, -121.818889, -121.8075, -121.793056, -121.796389, 
    -121.811389, NaN, -125.181278, -125.18125, -125.1775, -125.17, 
    -125.162944, -125.168361, -125.181278, NaN, -122.768889, -122.768028, 
    -122.766778, -122.763889, -122.758028, -122.761806, -122.768889, NaN, 
    -123.426361, -123.4255, -123.423472, -123.412639, -123.407194, 
    -123.420139, -123.426361, NaN, -124.032083, -124.031, -124.018694, 
    -124.013611, -124.029222, -124.034, -124.032083, NaN, -124.024889, 
    -124.02575, -124.029056, -124.030222, -124.02125, -124.021861, 
    -124.024889, NaN, -123.027278, -123.027278, -123.023444, -123.019222, 
    -123.020944, -123.025194, -123.027278, NaN, -122.713861, -122.713861, 
    -122.701806, -122.69475, -122.698472, -122.704278, -122.713861, NaN, 
    -116.801611, -116.800222, -116.801639, -116.804778, -116.811556, 
    -116.808861, -116.801611, NaN, -123.301333, -123.300556, -123.299278, 
    -123.288417, -123.281333, -123.282611, -123.301333, NaN, -122.553833, 
    -122.553917, -122.552583, -122.548472, -122.543861, -122.548472, 
    -122.553833, NaN, -122.781389, -122.781417, -122.774278, -122.769694, 
    -122.780167, -122.778083, -122.781389, NaN, -115.543833, -115.544083, 
    -115.544139, -115.537472, -115.529861, -115.5375, -115.543833, NaN, 
    -124.003528, -124.004222, -124.009417, -124.006083, -123.998806, 
    -123.999167, -124.003528, NaN, -122.714667, -122.714667, -122.707667, 
    -122.687167, -122.691722, -122.706778, -122.714667, NaN, -118.283889, 
    -118.282583, -118.279833, -118.281722, -118.290806, -118.289028, 
    -118.283889, NaN, -122.838, -122.837222, -122.835917, -122.827667, 
    -122.824694, -122.832611, -122.838, NaN, -125.351306, -125.351306, 
    -125.345806, -125.332972, -125.342528, -125.351306, NaN, -123.713861, 
    -123.713861, -123.711722, -123.70175, -123.692111, -123.713861, NaN, 
    -123.963861, -123.963778, -123.961306, -123.955889, -123.960472, 
    -123.963861, NaN, -122.539722, -122.539722, -122.529306, -122.524722, 
    -122.527583, -122.539722, NaN, -122.578889, -122.578861, -122.574306, 
    -122.559694, -122.560944, -122.578889, NaN, -125.387917, -125.387917, 
    -125.381722, -125.377917, -125.383333, -125.387917, NaN, -123.66875, 
    -123.66875, -123.645861, -123.641306, -123.652528, -123.66875, NaN, 
    -122.616389, -122.616389, -122.600944, -122.600472, -122.609278, 
    -122.616389, NaN, -123.993806, -123.993778, -123.980889, -123.971667, 
    -123.969583, -123.993806, NaN, -123.28725, -123.287194, -123.272639, 
    -123.27225, -123.278444, -123.28725, NaN, -122.973917, -122.972694, 
    -122.967583, -122.941417, -122.951, -122.973917, NaN, -114.475, 
    -114.474167, -114.474, -114.476806, -114.480944, -114.475, NaN, 
    -119.830583, -119.829389, -119.824472, -119.829111, -119.832083, 
    -119.830583, NaN, -116.792639, -116.792028, -116.787472, -116.786833, 
    -116.799222, -116.792639, NaN, -125.519639, -125.519583, -125.517528, 
    -125.510889, -125.514139, -125.519639, NaN, -117.250972, -117.248556, 
    -117.241639, -117.239222, -117.245111, -117.250972, NaN, -125.277056, 
    -125.277139, -125.265056, -125.265833, -125.271667, -125.277056, NaN, 
    -123.674639, -123.674556, -123.664222, -123.652139, -123.655028, 
    -123.674639, NaN, -118.293583, -118.292278, -118.297528, -118.3, 
    -118.298139, -118.293583, NaN, -123.633833, -123.633861, -123.630083, 
    -123.623833, -123.625083, -123.633833, NaN, -123.252167, -123.252222, 
    -123.244333, -123.241389, -123.250083, -123.252167, NaN, -122.493056, 
    -122.493028, -122.487611, -122.480556, -122.490083, -122.493056, NaN, 
    -119.364139, -119.359611, -119.357417, -119.363306, -119.380889, 
    -119.364139, NaN, -123.545444, -123.545028, -123.524194, -123.517917, 
    -123.541694, -123.545444, NaN, -123.879611, -123.879556, -123.863361, 
    -123.854583, -123.866639, -123.879611, NaN, -123.548889, -123.548944, 
    -123.547694, -123.538444, -123.537639, -123.548889, NaN, -123.328861, 
    -123.328889, -123.321778, -123.3155, -123.318444, -123.328861, NaN, 
    -123.259722, -123.259722, -123.253417, -123.253444, -123.255944, 
    -123.259722, NaN, -125.352083, -125.351306, -125.346667, -125.339556, 
    -125.349222, -125.352083, NaN, -125.331278, -125.330028, -125.321694, 
    -125.321694, -125.328333, -125.331278, NaN, -125.096278, -125.096278, 
    -125.094222, -125.088, -125.089167, -125.096278, NaN, -123.612972, 
    -123.612972, -123.579222, -123.580139, -123.594333, -123.612972, NaN, 
    -115.384, -115.384194, -115.374444, -115.372528, -115.381028, -115.384, 
    NaN, -122.850556, -122.849361, -122.837611, -122.828028, -122.837611, 
    -122.850556, NaN, -122.50975, -122.508861, -122.505944, -122.493889, 
    -122.498444, -122.50975, NaN, -114.087583, -114.088194, -114.091056, 
    -114.089278, -114.085861, -114.087583, NaN, -114.069917, -114.06925, 
    -114.071083, -114.075917, -114.071083, -114.069917, NaN, -120.329528, 
    -120.328556, -120.331361, -120.338, -120.333722, -120.329528, NaN, 
    -123.697222, -123.69725, -123.687167, -123.691806, -123.693444, 
    -123.697222, NaN, -125.383722, -125.383806, -125.377528, -125.373806, 
    -125.375917, -125.383722, NaN, -124.027833, -124.029778, -124.036833, 
    -124.044417, -124.041778, -124.027833, NaN, -122.364611, -122.363389, 
    -122.356722, -122.352083, -122.358417, -122.364611, NaN, -123.323861, 
    -123.323861, -123.320944, -123.314722, -123.318472, -123.323861, NaN, 
    -123.6105, -123.610528, -123.602611, -123.600556, -123.605167, -123.6105, 
    NaN, -123.089694, -123.089694, -123.086778, -123.079722, -123.080972, 
    -123.089694, NaN, -114.074222, -114.073611, -114.071306, -114.069194, 
    -114.071444, -114.074222, NaN, -124.653917, -124.653167, -124.647056, 
    -124.643917, -124.651889, -124.653917, NaN, -122.842167, -122.842167, 
    -122.840083, -122.83675, -122.838472, -122.842167, NaN, -122.390528, 
    -122.390528, -122.386806, -122.384722, -122.389278, -122.390528, NaN, 
    -123.00175, -123, -123, -123.009667, -123.008444, -123.00175, NaN, 
    -114.498111, -114.498278, -114.49925, -114.495917, -114.494278, 
    -114.498111, NaN, -125.416278, -125.414583, -125.413417, -125.405472, 
    -125.410028, -125.416278, NaN, -123.41475, -123.41475, -123.407611, 
    -123.401361, -123.410167, -123.41475, NaN, -123.752139, -123.752167, 
    -123.745028, -123.744194, -123.749194, -123.752139, NaN, -125.3705, 
    -125.370417, -125.365, -125.359667, -125.363389, -125.3705, NaN, 
    -117.26375, -117.262333, -117.256722, -117.258333, -117.261583, 
    -117.26375, NaN, -122.560528, -122.559778, -122.559306, -122.55475, 
    -122.556833, -122.560528, NaN, -124.738778, -124.738833, -124.735861, 
    -124.731278, -124.735056, -124.738778, NaN, -124.092722, -124.096861, 
    -124.09575, -124.089806, -124.088389, -124.092722, NaN, -125.253722, 
    -125.253778, -125.245417, -125.247528, -125.253722, NaN, -125.291278, 
    -125.29, -125.283778, -125.285083, -125.291278, NaN, -122.851389, 
    -122.851389, -122.845139, -122.846806, -122.851389, NaN, -114.146056, 
    -114.146056, -114.138333, -114.138668045857, NaN, NaN, -123.673861, 
    -123.673861, -123.658028, -123.667667, -123.673861, NaN, -125.364611, 
    -125.364556, -125.354556, -125.356722, -125.364611, NaN, -123.624611, 
    -123.624667, -123.613778, -123.618333, -123.624611, NaN, -123.522972, 
    -123.523028, -123.511278, -123.517528, -123.522972, NaN, -125.320444, 
    -125.320444, -125.312972, -125.3175, -125.320444, NaN, -123.96875, 
    -123.96875, -123.96425, -123.962139, -123.96875, NaN, -124.60125, 
    -124.601306, -124.595889, -124.594194, -124.60125, NaN, -124.758056, 
    -124.758083, -124.752611, -124.747222, -124.758056, NaN, -123.39725, 
    -123.397167, -123.391361, -123.390917, -123.39725, NaN, -123.093056, 
    -123.093111, -123.084667, -123.088389, -123.093056, NaN, -120.458639, 
    -120.459389, -120.461389, -120.454778, -120.458639, NaN, -122.738833, 
    -122.738056, -122.733417, -122.73475, -122.738833, NaN, -122.779694, 
    -122.779694, -122.775194, -122.775583, -122.779694, NaN, -114.069194, 
    -114.070611, -114.07275, -114.066028, -114.069194, NaN, -125.584639, 
    -125.584611, -125.578333, -125.572139, -125.584639, NaN, -123.594806, 
    -123.59325, -123.590944, -123.5955, -123.594806, NaN, -122.895111, 
    -122.895556, -122.882639, -122.881861, -122.895111, NaN, -125.089639, 
    -125.089556, -125.078722, -125.085056, -125.089639, NaN, -123.018806, 
    -123.018028, -123.014361, -123.015528, -123.018806, NaN, -123.242194, 
    -123.242194, -123.236833, -123.229667, -123.242194, NaN, -120.43625, 
    -120.434389, -120.434778, -120.441556, -120.43625, NaN, -114.072667, 
    -114.073278, -114.076917, -114.069528, -114.072667, NaN, -123.17225, 
    -123.17225, -123.16175, -123.161417, -123.17225, NaN, -124.996972, 
    -124.997028, -124.990778, -124.987056, -124.996972, NaN, -124.509417, 
    -124.507861, -124.505972, -124.5115, -124.509417, NaN, -123.019778, 
    -123.019778, -123.010528, -123.017694, -123.019778, NaN, -123.308, 
    -123.308, -123.304278, -123.303, -123.308, NaN, -122.930556, -122.930556, 
    -122.926806, -122.923083, -122.930556, NaN, -122.582194, -122.582194, 
    -122.576417, -122.579278, -122.582194, NaN, -123.401389, -123.401417, 
    -123.395972, -123.3955, -123.401389, NaN, -123.243944, -123.241778, 
    -123.233444, -123.234278, -123.243944, NaN, -123.189667, -123.189667, 
    -123.17975, -123.182639, -123.189667, NaN, -124.07525, -124.074083, 
    -124.069056, -124.073611, -124.07525, NaN, -125.372972, -125.372972, 
    -125.366306, -125.368361, -125.372972, NaN, -114.982056, -114.984, 
    -114.985028, -114.980833, -114.982056, NaN, -125.321333, -125.321222, 
    -125.310861, -125.311667, -125.321333, NaN, -123.684722, -123.683444, 
    -123.6755, -123.677583, -123.684722, NaN, -123.010417, -123.011833, 
    -123.015639, -123.014139, -123.010417, NaN, -122.932167, -122.932167, 
    -122.918, -122.928389, -122.932167, NaN, -123.244722, -123.244722, 
    -123.239306, -123.23475, -123.244722, NaN, -123.628917, -123.628056, 
    -123.625056, -123.624278, -123.628917, NaN, -125.320389, -125.320472, 
    -125.314583, -125.315889, -125.320389, NaN, -115.504389, -115.503917, 
    -115.500917, -115.502694, -115.504389, NaN, -123.499583, -123.499583, 
    -123.495028, -123.495028, -123.499583, NaN, -115.356556, -115.3565, 
    -115.353444, -115.355028, -115.356556, NaN, -125.647111, -125.647139, 
    -125.645028, -125.642111, -125.647111, NaN, -125.390528, -125.389583, 
    -125.385417, -125.3875, -125.390528, NaN, -125.120417, -125.120028, 
    -125.10625, -125.116694, -125.120417, NaN, -123.452167, -123.452167, 
    -123.441306, -123.445139, -123.452167, NaN, -114.280917, -114.279778, 
    -114.274167, -114.27875, -114.280917, NaN, -114.4125, -114.412278, 
    -114.417333, -114.414278, -114.4125, NaN, -123.327167, -123.327194, 
    -123.320972, -123.3155, -123.327167, NaN, -123.34225, -123.34225, 
    -123.334278, -123.330972, -123.34225, NaN, -123.629778, -123.629222, 
    -123.621833, -123.618472, -123.629778, NaN, -125.174583, -125.174639, 
    -125.165833, -125.166667, -125.174583, NaN, -125.297944, -125.297944, 
    -125.294222, -125.288028, -125.297944, NaN, -115.355972, -115.355806, 
    -115.351556, -115.353528, -115.355972, NaN, -117.300306, -117.297278, 
    -117.293222, -117.300333, -117.300306, NaN, -115.36175, -115.361639, 
    -115.358444, -115.357694, -115.36175, NaN, -123.993806, -123.993861, 
    -123.987556, -123.983806, -123.993806, NaN, -123.733806, -123.733806, 
    -123.72375, -123.730028, -123.733806, NaN, -123.033556, -123.033972, 
    -123.031944, -123.030917, -123.033556, NaN, -123.457083, -123.457083, 
    -123.438722, -123.436694, -123.457083, NaN, -115.365917, -115.365583, 
    -115.356806, -115.363222, -115.365917, NaN, -114.877472, -114.875917, 
    -114.874917, -114.878306, -114.877472, NaN, -125.527972, -125.527972, 
    -125.525, -125.523722, -125.527972, NaN, -125.377139, -125.377056, 
    -125.374167, -125.3705, -125.377139, NaN, -122.4705, -122.470028, 
    -122.465472, -122.468417, -122.4705, NaN, -122.426278, -122.426278, 
    -122.420472, -122.423361, -122.426278, NaN, -123.388861, -123.388861, 
    -123.3855, -123.386806, -123.388861, NaN, -123.269694, -123.269722, 
    -123.263861, -123.265139, -123.269694, NaN, -125.328806, -125.328806, 
    -125.323306, -125.323333, -125.328806, NaN, -125.205444, -125.205417, 
    -125.200889, -125.199583, -125.205444, NaN, -125.313778, -125.313861, 
    -125.310028, -125.309167, -125.313778, NaN, -124.548472, -124.548944, 
    -124.546, -124.542667, -124.548472, NaN, -122.899667, -122.899667, 
    -122.898444, -122.894778, -122.899667, NaN, -114.164806, -114.16575, 
    -114.16375, -114.161917, -114.164806, NaN, -123.281333, -123.280556, 
    -123.27675, -123.275583, -123.281333, NaN, -123.982333, -123.982583, 
    -123.98475, -123.986861, -123.982333, NaN, -125.334639, -125.334667, 
    -125.330889, -125.330417, -125.334639, NaN, -122.976389, -122.976389, 
    -122.972667, -122.968889, -122.976389, NaN, -123.155528, -123.155528, 
    -123.15175, -123.150528, -123.155528, NaN, -125.326333, -125.326333, 
    -125.320917, -125.319556, -125.326333, NaN, -125.269611, -125.269583, 
    -125.263778, -125.265056, -125.269611, NaN, -125.211306, -125.211306, 
    -125.206667, -125.206667, -125.211306, NaN, -125.377083, -125.377083, 
    -125.374194, -125.372056, -125.377083, NaN, -125.329583, -125.329639, 
    -125.325, -125.322917, -125.329583, NaN, -125.117083, -125.117167, 
    -125.112083, -125.115861, -125.117083, NaN, -123.392167, -123.391389, 
    -123.38925, -123.388056, -123.392167, NaN, -122.541361, -122.541361, 
    -122.537583, -122.537139, -122.541361, NaN, -119.049361, -119.048222, 
    -119.045639, -119.047694, -119.049361, NaN, -123.013861, -123.013444, 
    -123.008889, -123.010972, -123.013861, NaN, -115.768361, -115.767583, 
    -115.77075, -115.770972, -115.768361, NaN, -123.60975, -123.608889, 
    -123.605167, -123.604667, -123.60975, NaN, -117.26425, -117.26175, 
    -117.260778, -117.263944, -117.26425, NaN, -124.63125, -124.629889, 
    -124.630389, -124.63125, NaN, -115.811806, -115.810861, -115.810694, 
    -115.811806, NaN, -115.7875, -115.786917, -115.786889, -115.7875, NaN, 
    -118.37075, -118.369861, -118.369167, -118.37075, NaN, -115.781111, 
    -115.780444, -115.780139, -115.781111, NaN, -115.788306, -115.787444, 
    -115.786278, -115.788306, NaN, -115.775972, -115.775778, -115.774278, 
    -115.775972, NaN, -115.69075, -115.689694, -115.689111, -115.69075, NaN, 
    -123.986667, -123.986556, -123.990889, -123.986667, NaN, -114.068333, 
    -114.068639, -114.068639, -114.068333, NaN, -124.727472, -124.726917, 
    -124.73275, -124.727472, NaN, -122.828861, -122.828861, -122.821306, 
    -122.828861, NaN, -115.778389, -115.779111, -115.776389, -115.778389, 
    NaN, -115.783611, -115.783083, -115.782333, -115.783611, NaN, 
    -115.784972, -115.784333, -115.784361, -115.784972, NaN, -115.802917, 
    -115.802861, -115.803278, -115.802917, NaN, -125.097917, -125.097944, 
    -125.092917, -125.097917, NaN, -125.472972, -125.472944, -125.467972, 
    -125.472972, NaN, -123.276361, -123.276361, -123.269722, -123.276361, 
    NaN, -123.292222, -123.292222, -123.283083, -123.292222, NaN, 
    -123.458889, -123.458889, -123.453861, -123.458889, NaN, -122.482222, 
    -122.482194, -122.474722, -122.482222, NaN, -124.422083, -124.421306, 
    -124.421389, -124.422083, NaN, -125.137139, -125.134222, -125.128806, 
    -125.137139, NaN, -125.101306, -125.101306, -125.097139, -125.101306, 
    NaN, -124.593583, -124.592333, -124.594444, -124.593583, NaN, 
    -123.647972, -123.647944, -123.642111, -123.647972, NaN, -125.337917, 
    -125.336694, -125.332194, -125.337917, NaN, -125.288833, -125.288806, 
    -125.281306, -125.288833, NaN, -125.357111, -125.357194, -125.352167, 
    -125.357111, NaN, -123.987361, -123.987389, -123.991167, -123.987361, 
    NaN, -123.94925, -123.949472, -123.954444, -123.94925, NaN, -125.292944, 
    -125.292972, -125.28625, -125.292944, NaN, -125.015472, -125.015444, 
    -125.011278, -125.015472, NaN, -123.531222, -123.531111, -123.529778, 
    -123.531222, NaN, -123.642222, -123.64225, -123.638472, -123.642222, NaN, 
    -123.65475, -123.65475, -123.650972, -123.65475, NaN, -123.67975, 
    -123.679278, -123.6785, -123.67975, NaN, -123.6355, -123.6355, 
    -123.632194, -123.6355, NaN, -123.332194, -123.332194, -123.329333, 
    -123.332194, NaN, -123.134722, -123.134722, -123.128917, -123.134722, 
    NaN, -122.341278, -122.34125, -122.335444, -122.341278, NaN, -123.330583, 
    -123.330139, -123.327639, -123.330583, NaN, -123.439667, -123.439722, 
    -123.433861, -123.439667, NaN, -123.376444, -123.376361, -123.3705, 
    -123.376444, NaN, -123.277278, -123.277278, -123.273889, -123.277278, 
    NaN, -118.29125, -118.292028, -118.2915, -118.29125, NaN, -122.92475, 
    -122.924333, -122.917583, -122.92475, NaN, -122.572222, -122.572222, 
    -122.568, -122.572222, NaN, -123.472278, -123.472167, -123.468889, 
    -123.472278, NaN, -123.273056, -123.271778, -123.267167, -123.273056, 
    NaN, -123.134722, -123.134722, -123.130556, -123.134722, NaN, 
    -123.273111, -123.272583, -123.269306, -123.273111, NaN, -123.710556, 
    -123.70975, -123.705528, -123.710556, NaN, -125.327083, -125.326722, 
    -125.323722, -125.327083, NaN, -123.817111, -123.816278, -123.813361, 
    -123.817111, NaN, -123.902056, -123.901278, -123.898722, -123.902056, 
    NaN, -125.245417, -125.245444, -125.243333, -125.245417, NaN, 
    -125.299639, -125.299556, -125.295417, -125.299639, NaN, -115.808028, 
    -115.807222, -115.806806, -115.808028, NaN, -115.810194, -115.809528, 
    -115.8095, -115.810194, NaN, -123.105639, -123.107972, -123.106667, 
    -123.105639, NaN, -123.481333, -123.48125, -123.475417, -123.481333, NaN, 
    -123.628806, -123.628806, -123.621333, -123.628806, NaN, -115.764194, 
    -115.7655, -115.764222, -115.764194, NaN, -123.302194, -123.302194, 
    -123.294639, -123.302194, NaN, -125.362167, -125.362139, -125.353778, 
    -125.362167, NaN, -123.102556, -123.103694, -123.101861, -123.102556, 
    NaN, -123.763778, -123.763833, -123.757972, -123.763778, NaN, 
    -123.566222, -123.566278, -123.559611, -123.566222, NaN, -123.637972, 
    -123.636667, -123.630861, -123.637972, NaN, -123.983417, -123.981722, 
    -123.987222, -123.983417, NaN, -124.686556, -124.687972, -124.685694, 
    -124.686556, NaN, -118.301611, -118.300528, -118.299194, -118.301611, 
    NaN, -115.765417, -115.765111, -115.767167, -115.765417, NaN, 
    -124.696389, -124.697833, -124.693694, -124.696389, NaN, -125.297083, 
    -125.297167, -125.292139, -125.297083, NaN, -123.213083, -123.213083, 
    -123.206389, -123.213083, NaN, -122.829722, -122.829722, -122.822222, 
    -122.829722, NaN, -114.070111, -114.07075, -114.071361, -114.070111, NaN, 
    -125.354639, -125.354583, -125.349611, -125.354639, NaN, -114.442472, 
    -114.442722, -114.441111, -114.442472, NaN, -123.126139, -123.127056, 
    -123.127722, -123.126139, NaN, -123.438556, -123.437472, -123.437861, 
    -123.438556, NaN, -123.050583, -123.049778, -123.050139, -123.050583, 
    NaN, -118.617111, -118.617056, -118.612944, -118.617111, NaN, 
    -115.772639, -115.773639, -115.771833, -115.772639, NaN, -123.858806, 
    -123.858806, -123.853333, -123.858806, NaN, -114.627444, -114.626611, 
    -114.628444, -114.627444, NaN, -114.356889, -114.355167, -114.354639, 
    -114.356889, NaN, -123.217972, -123.217639, -123.210944, -123.217972, 
    NaN, -123.1, -123.098278, -123.095889, -123.1, NaN, -122.473833, 
    -122.473778, -122.471278, -122.473833, NaN, -115.815083, -115.814278, 
    -115.814917, -115.815083, NaN, -115.761167, -115.760861, -115.764444, 
    -115.761167, NaN, -115.436833, -115.435778, -115.434194, -115.436833, 
    NaN, -123.141333, -123.140139, -123.137194, -123.141333, NaN, 
    -125.042083, -125.041278, -125.037056, -125.042083, NaN, -122.482222, 
    -122.481806, -122.477167, -122.482222, NaN, -118.593778, -118.593806, 
    -118.590389, -118.593778, NaN, -122.893083, -122.893083, -122.889694, 
    -122.893083, NaN, -123.396417, -123.396333, -123.391389, -123.396417, 
    NaN, -123.300556, -123.300472, -123.297194, -123.300556, NaN, 
    -123.463889, -123.462611, -123.460528, -123.463889, NaN, -123.041389, 
    -123.041389, -123.032222, -123.041389, NaN, -123.278861, -123.278861, 
    -123.2755, -123.278861, NaN, -123.684694, -123.68425, -123.681778, 
    -123.684694, NaN, -124.763056, -124.763056, -124.758944, -124.763056, 
    NaN, -124.758083, -124.758056, -124.754694, -124.758083, NaN, 
    -125.172083, -125.172111, -125.168778, -125.172083, NaN, -125.307917, 
    -125.308, -125.304583, -125.307917, NaN, -125.321306, -125.321333, 
    -125.317139, -125.321306, NaN, -125.154667, -125.154556, -125.1505, 
    -125.154667, NaN, -125.242889, -125.242944, -125.240861, -125.242889, 
    NaN, -125.123778, -125.123806, -125.120833, -125.123778, NaN, 
    -125.235444, -125.235056, -125.231278, -125.235444, NaN, -125.386278, 
    -125.386306, -125.382944, -125.386278, NaN, -125.366222, -125.36625, 
    -125.362139, -125.366222, NaN, -123.717111, -123.717139, -123.713778, 
    -123.717111, NaN, -115.817167, -115.817361, -115.815056, -115.817167, 
    NaN, -115.808778, -115.807861, -115.807361, -115.808778, NaN, 
    -115.774444, -115.774389, -115.776667, -115.774444, NaN, -124.015056, 
    -124.015139, -124.012194, -124.015056, NaN, -123.981111, -123.982278, 
    -123.983583, -123.981111, NaN, -115.554222, -115.553889, -115.551556, 
    -115.554222, NaN, -123.688028, -123.687639, -123.682667, -123.688028, 
    NaN, -115.538194, -115.537917, -115.535806, -115.538194, NaN, 
    -115.568444, -115.568361, -115.567278, -115.568444, NaN, -115.559083, 
    -115.558889, -115.556806, -115.559083, NaN, -115.5615, -115.561444, 
    -115.559111, -115.5615, NaN, -115.570861, -115.570722, -115.568583, 
    -115.570861, NaN, -115.350944, -115.350778, -115.348611, -115.350944, 
    NaN, -115.577417, -115.577306, -115.575056, -115.577417, NaN, 
    -115.575028, -115.574778, -115.5725, -115.575028, NaN, -115.548333, 
    -115.547944, -115.545611, -115.548333, NaN, -115.791861, -115.791528, 
    -115.789167, -115.791861, NaN, -123.486361, -123.486361, -123.474694, 
    -123.486361, NaN, -115.281611, -115.281556, -115.279417, -115.281611, 
    NaN, -115.601472, -115.601472, -115.599389, -115.601472, NaN, 
    -115.565056, -115.564917, -115.562472, -115.565056, NaN, -115.341722, 
    -115.341667, -115.33975, -115.341722, NaN, -122.372917, -122.372972, 
    -122.3705, -122.372917, NaN, -123.907083, -123.905056, -123.902972, 
    -123.907083, NaN, -123.895472, -123.8955, -123.892083, -123.895472, NaN, 
    -125.114611, -125.114167, -125.112056, -125.114611, NaN, -125.347917, 
    -125.347528, -125.345889, -125.347917, NaN, -123.488056, -123.487972, 
    -123.483806, -123.488056, NaN, -123.379694, -123.379694, -123.376361, 
    -123.379694, NaN, -122.824778, -122.824778, -122.821361, -122.824778, 
    NaN, -123.615528, -123.615083, -123.610972, -123.615528, NaN, 
    -122.914667, -122.914667, -122.911417, -122.914667, NaN, -122.8705, 
    -122.870139, -122.868472, -122.8705, NaN, -115.543167, -115.543028, 
    -115.54075, -115.543167, NaN, -115.570611, -115.570611, -115.567639, 
    -115.570611, NaN, -123.329667, -123.329667, -123.326389, -123.329667, 
    NaN, -123.651389, -123.650972, -123.649278, -123.651389, NaN, -123.6605, 
    -123.660083, -123.655944, -123.6605, NaN, -125.163806, -125.163333, 
    -125.160472, -125.163806, NaN, -115.261472, -115.261722, -115.25925, 
    -115.261472, NaN, -115.355333, -115.355333, -115.351083, -115.355333, 
    NaN, -115.361028, -115.360639, -115.358444, -115.361028, NaN, 
    -115.329417, -115.329222, -115.325972, -115.329417, NaN, -115.256778, 
    -115.256639, -115.253417, -115.256778, NaN, -115.350694, -115.350639, 
    -115.34775, -115.350694, NaN, -115.358556, -115.358472, -115.355833, 
    -115.358556, NaN, -115.377444, -115.37725, -115.372611, -115.377444, NaN ;

 lat_coast = NaN, NaN, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28.008611, 31.564194, 31.565, 
    31.568528, 31.584444, 31.589889, 31.587611, 31.594694, 31.599056, 
    31.599806, 31.604972, 31.595472, 31.594389, 31.588583, 31.586333, 
    31.600667, 31.610278, 31.611639, 31.618694, 31.619139, 31.614361, 
    31.61275, 31.623444, 31.604111, 31.609556, 31.613667, 31.617639, 
    31.612639, 31.604889, 31.613167, 31.618444, 31.618306, 31.621667, 
    31.624778, 31.620917, 31.620194, 31.614278, 31.618861, 31.624028, 
    31.621528, 31.624444, 31.636694, 31.626056, 31.608944, 31.604806, 
    31.611389, 31.615361, 31.628361, 31.630972, 31.617389, 31.616472, 
    31.630861, 31.641944, 31.648028, 31.644389, 31.660167, 31.638861, 
    31.618556, 31.605361, 31.585944, 31.583278, 31.582806, 31.596583, 
    31.591389, 31.587861, 31.588917, 31.575611, 31.573611, 31.571556, 
    31.568556, 31.568417, 31.564139, 31.560722, 31.58025, 31.56325, 
    31.544833, 31.539833, 31.5233866447477, 31.52225, 31.525, 31.531972, 
    31.536556, 31.539306, 31.542861, 31.538917, 31.540083, 31.536611, 
    31.533806, 31.520694, 31.522, 31.517944, 31.513028, 31.5115, 31.514861, 
    31.509583, 31.508889, 31.506639, 31.508222, 31.51825, 31.525806, 
    31.523167, 31.516917, 31.503833, 31.493333, 31.489806, 31.488083, 
    31.491667, 31.490472, 31.493861, 31.507139, 31.527361, 31.544167, 
    31.560917, 31.576417, 31.581556, 31.593, 31.598111, 31.607944, 31.628139, 
    31.634889, 31.645611, 31.648306, 31.652056, 31.659861, 31.670333, 
    31.676778, 31.680639, 31.691611, 31.696583, 31.703528, 31.720139, 
    31.735889, 31.748972, 31.778139, 31.753139, 31.763472, 31.760667, 
    31.763306, 31.772722, 31.813278, 31.820861, 31.834139, 31.824305, 
    31.821472, 31.822278, 31.839833, 31.854667, 31.864111, 31.874306, 
    31.871611, 31.884306, 31.873472, 31.868556, 31.864194, 31.868528, 31.881, 
    31.870889, 31.864194, 31.863361, 31.86925, 31.869083, 31.860556, 
    31.852389, 31.83425, 31.829139, 31.831361, 31.809333, 31.807444, 
    31.810083, 31.807333, 31.831639, 31.806528, 31.809222, 31.806583, 
    31.807778, 31.7895, 31.734972, 31.682167, 31.664139, 31.639139, 31.6225, 
    31.61225, 31.610278, 31.601139, 31.598333, 31.587611, 31.580917, 
    31.564333, 31.551583, 31.530556, 31.488528, 31.459944, 31.434583, 
    31.425361, 31.418111, 31.408167, 31.40575, 31.394889, 31.369028, 
    31.310417, 31.301194, 31.298944, 31.287389, 31.285, 31.293389, 31.302639, 
    31.292361, 31.288917, 31.289889, 31.30225, 31.290972, 31.289167, 
    31.289068, 31.284417, 31.280889, 31.274833, 31.280111, 31.266028, 
    31.261889, 31.268111, 31.271694, 31.273333, 31.278056, 31.273306, 
    31.268083, 31.264778, 31.2775, 31.265722, 31.266639, 31.265, 31.261917, 
    31.258306, 31.260694, 31.256583, 31.267861, 31.259222, 31.26325, 
    31.258278, 31.258, 31.253861, 31.256833, 31.255194, 31.249194, 31.253306, 
    31.247778, 31.244639, 31.24475, 31.239583, 31.241167, 31.234611, 
    31.236778, 31.243111, 31.235833, 31.233389, 31.230944, 31.256694, 
    31.265833, 31.254889, 31.239583, 31.2365, 31.232472, 31.236, 31.237611, 
    31.249667, 31.25175, 31.236583, 31.207611, 31.208556, 31.217972, 
    31.211556, 31.218083, 31.210528, 31.205833, 31.204944, 31.157722, 
    31.118722, 31.093472, 31.088944, 31.083222, 31.074, 31.069, 31.055944, 
    31.055583, 31.049111, 31.043778, 31.040556, 31.022056, 31.008333, 
    31.001111, 30.990194, 30.978333, 30.9375, 30.912694, 30.878944, 30.87575, 
    30.876472, 30.868167, 30.847611, 30.819889, 30.790583, 30.815056, 
    30.812417, 30.785444, 30.758083, 30.757167, 30.754306, 30.744083, 
    30.739056, 30.714139, 30.681639, 30.629333, 30.587278, 30.577611, 
    30.566639, 30.557028, 30.545583, 30.538806, 30.530722, 30.500806, 
    30.491444, 30.470139, 30.457, 30.441861, 30.419111, 30.373972, 30.364611, 
    30.346528, 30.343944, 30.348139, 30.339389, 30.337694, 30.31525, 
    30.297056, 30.289083, 30.284306, 30.27925, 30.265333, 30.257417, 
    30.241444, 30.226667, 30.218139, 30.198194, 30.184806, 30.174472, 
    30.166778, 30.141694, 30.128833, 30.121083, 30.111972, 30.088222, 30.078, 
    30.069472, 30.052361, 30.032278, 30.026778, 30.011306, 30.002583, 
    29.983222, 29.969556, 29.95675, 29.95425, 29.949861, 29.912583, 
    29.908861, 29.909861, 29.889889, 29.869472, 29.849861, 29.829361, 
    29.826444, 29.824028, 29.825889, 29.820139, 29.814694, 29.809417, 
    29.802667, 29.800028, 29.809778, 29.808444, 29.801083, 29.791556, 
    29.775944, 29.771556, 29.77075, 29.760056, 29.747556, 29.743222, 
    29.741556, 29.745861, 29.742417, 29.742361, 29.758333, 29.756389, 
    29.759278, 29.755806, 29.758278, 29.766361, 29.765667, 29.771472, 
    29.773306, 29.769139, 29.764111, 29.768361, 29.766806, 29.760639, 
    29.763306, 29.750028, 29.744194, 29.727333, 29.707194, 29.700472, 
    29.690778, 29.694139, 29.692472, 29.674111, 29.662833, 29.652306, 
    29.640611, 29.630528, 29.597306, 29.594556, 29.580611, 29.581472, 
    29.581472, 29.566806, 29.554972, 29.5395, 29.526639, 29.522389, 
    29.514778, 29.505, 29.486528, 29.475722, 29.465, 29.459139, 29.453306, 
    29.438278, 29.432333, 29.427389, 29.420917, 28.003472, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28.021611, 28.088361, 28.091028, 
    28.0885, 28.053472, 28.044917, 28.040111, 28.023194, 28.011778, 
    28.000639, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28.004722, 28.005361, 28.019389, 28.015139, 
    28.016861, 28.022028, 28.026806, 28.030972, 28.037361, 28.03625, 
    28.032167, 28.032778, 28.02125, 28.026472, 28.022417, 28.014, 28.009556, 
    28.006694, 28.006, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28.027611, 
    28.044278, 28.041639, 28.055, 28.047806, 28.052778, 28.083611, 28.115, 
    28.124472, 28.157306, 28.189028, 28.195083, 28.193333, 28.186194, 
    28.17175, 28.145028, 28.11475, 28.109056, 28.110111, 28.105194, 
    28.113278, 28.111111, 28.114139, 28.119889, 28.121833, 28.118556, 
    28.121306, 28.126139, 28.129444, 28.13375, 28.136194, 28.149889, 
    28.156611, 28.160417, 28.162639, 28.186194, 28.218139, 28.196444, 
    28.194111, 28.203222, 28.21825, 28.236, 28.238806, 28.259472, 28.258278, 
    28.262917, 28.258444, 28.256667, 28.253806, 28.249583, 28.249, 28.252722, 
    28.249972, 28.24975, 28.246639, 28.240139, 28.241139, 28.252028, 
    28.257694, 28.34225, 28.391083, 28.427611, 28.465139, 28.474194, 
    28.487583, 28.499278, 28.510917, 28.519917, 28.524222, 28.547417, 
    28.55975, 28.563111, 28.559667, 28.56875, 28.594528, 28.623, 28.636444, 
    28.655667, 28.66575, 28.663889, 28.653861, 28.66325, 28.660667, 
    28.688139, 28.705639, 28.706556, 28.703222, 28.70575, 28.721944, 
    28.726556, 28.730222, 28.738194, 28.738167, 28.742778, 28.755917, 
    28.757944, 28.766306, 28.769861, 28.773083, 28.779833, 28.795222, 
    28.811639, 28.8125, 28.806417, 28.817056, 28.829722, 28.834472, 
    28.858917, 28.874556, 28.883389, 28.875222, 28.887833, 28.90625, 
    28.907306, 28.921528, 28.931722, 28.934389, 28.930056, 28.930944, 
    28.927389, 28.923056, 28.918667, 28.927694, 28.935611, 28.944056, 
    28.959833, 28.973806, 28.973028, 28.969972, 28.967556, 28.964889, 
    28.968444, 28.975778, 28.990222, 28.993444, 28.998694, 29.009528, 
    29.017472, 29.019333, 29.024083, 29.060167, 29.062889, 29.080667, 
    29.092194, 29.096806, 29.096556, 29.108306, 29.110833, 29.109167, 
    29.102056, 29.100667, 29.110833, 29.109167, 29.119833, 29.132528, 
    29.136861, 29.134944, 29.138722, 29.157083, 29.173361, 29.181083, 
    29.183417, 29.180972, 29.195611, 29.194111, 29.19675, 29.210028, 
    29.210917, 29.236056, 29.240167, 29.236778, 29.244083, 29.258611, 
    29.268111, 29.273167, 29.283111, 29.284694, 29.295833, 29.30375, 
    29.310778, 29.315111, 29.359278, 29.373222, 29.380889, 29.380778, 
    29.38575, 29.396694, 29.405944, 29.415833, 29.417556, 29.420806, 
    29.418222, 29.422472, 29.420972, 29.429222, 29.431778, 29.427444, 
    29.446444, 29.475056, 29.476833, 29.483944, 29.485611, 29.499472, 
    29.512444, 29.524972, 29.53975, 29.541667, 29.554972, 29.55925, 
    29.557389, 29.561917, 29.571556, 29.576806, 29.591639, 29.622444, 
    29.625778, 29.625778, 29.616611, 29.615056, 29.621139, 29.633222, 
    29.642389, 29.656556, 29.662889, 29.678389, 29.690556, 29.696806, 
    29.694139, 29.742417, 29.750194, 29.754833, 29.80925, 29.830722, 
    29.898389, 29.926667, 29.947306, 29.958333, 29.957333, 29.947556, 
    29.948667, 30.000889, 30.090111, 30.111583, 30.115806, 30.132417, 
    30.151972, 30.199861, 30.243194, 30.2805, 30.299417, 30.309222, 
    30.315583, 30.339917, 30.352889, 30.369861, 30.393306, 30.4015, 
    30.404944, 30.402472, 30.392472, 30.394806, 30.411472, 30.408472, 
    30.411472, 30.409889, 30.413167, 30.42175, 30.430611, 30.447417, 
    30.460778, 30.459806, 30.462833, 30.485583, 30.483278, 30.490056, 
    30.496972, 30.498861, 30.506139, 30.501833, 30.497528, 30.492111, 
    30.479083, 30.477167, 30.471444, 30.469556, 30.463444, 30.454944, 
    30.44975, 30.442889, 30.438111, 30.434, 30.427111, 30.427417, 30.441611, 
    30.450806, 30.453722, 30.450417, 30.455389, 30.454167, 30.4425, 
    30.432472, 30.425806, 30.4085, 30.391778, 30.379111, 30.377528, 
    30.380417, 30.381528, 30.373889, 30.365944, 30.357222, 30.359306, 
    30.364972, 30.373306, 30.375861, 30.389139, 30.424167, 30.432917, 
    30.435806, 30.456639, 30.463306, 30.4725, 30.493306, 30.499111, 
    30.572472, 30.663306, 30.699972, 30.7175, 30.772444, 30.8025, 30.819583, 
    30.821194, 30.81875, 30.822889, 30.85875, 30.862056, 30.859556, 
    30.861278, 30.875389, 30.886667, 30.913306, 30.917944, 30.932917, 
    30.932056, 30.965361, 30.968722, 30.961222, 30.954583, 30.956222, 
    30.964167, 30.976639, 31.093528, 31.15275, 31.189556, 31.206944, 
    31.213139, 31.224861, 31.2405, 31.252, 31.256889, 31.266417, 31.282083, 
    31.284056, 31.2905, 31.291694, 31.302889, 31.309806, 31.321361, 
    31.322556, 31.329083, 31.329806, 31.334139, 31.345167, 31.3515, 
    31.360056, 31.361583, 31.368611, 31.376722, 31.405667, 31.409056, 
    31.414306, 31.434639, 31.444167, 31.451389, 31.463333, 31.464111, 
    31.459278, 31.461028, 31.495083, 31.514056, 31.515889, 31.513167, 
    31.517111, 31.527139, 31.533833, 31.534583, 31.54875, 31.553361, 
    31.549028, 31.55275, 31.559, 31.571389, 31.570722, 31.579056, 31.579083, 
    31.582667, 31.590528, 31.599833, 31.614639, 31.645417, 31.663972, 
    31.693194, 31.697722, 31.702583, 31.705444, 31.714556, 31.709833, 
    31.712306, 31.715, 31.723417, 31.720528, 31.730972, 31.732694, 31.739806, 
    31.742278, 31.744222, 31.748972, 31.749, 31.732611, 31.728389, 31.718333, 
    31.718306, 31.724806, 31.738417, 31.769361, 31.772278, 31.765139, 
    31.752917, 31.749556, 31.725417, 31.71675, 31.7065, 31.699167, 31.698056, 
    31.709167, 31.713722, 31.722194, 31.750056, 31.763222, 31.765722, 
    31.77075, 31.779889, 31.816472, 31.842944, 31.852722, 31.855972, 
    31.859222, 31.857944, 31.845861, 31.858278, 31.862639, 31.859833, 
    31.895083, 31.894778, 31.900639, 31.902361, 31.910917, 31.9595, 
    31.974944, 31.975694, 31.979944, 31.977417, 31.992139, 32.002694, 
    32.017944, 32.032944, 32.077861, 32.085361, 32.129722, 32.163528, 
    32.167306, 32.202944, 32.226444, 32.240306, 32.248222, 32.257333, 
    32.264194, 32.268167, 32.268667, 32.283389, 32.328917, 32.346611, 
    32.374167, 32.394028, 32.439694, 32.448722, 32.468889, 32.486861, 
    32.535833, 32.568306, 32.603028, 32.620889, 32.660778, 32.681944, 
    32.689083, 32.689139, 32.683083, 32.68725, 32.696361, 32.70825, 
    32.715833, 32.716611, 32.714667, 32.708361, 32.698889, 32.678833, 
    32.677389, 32.682556, 32.680667, 32.671611, 32.653417, 32.634583, 
    32.631389, 32.624556, 32.621028, 32.612944, 32.603722, 32.601556, 
    32.615139, 32.629417, 32.63975, 32.667722, 32.669944, 32.673556, 
    32.687278, 32.686944, 32.689861, 32.70975, 32.724972, 32.727667, 
    32.728194, 32.722333, 32.725028, 32.721583, 32.720917, 32.718278, 
    32.704778, 32.696222, 32.689083, 32.686056, 32.682444, 32.666639, 
    32.664833, 32.667472, 32.672972, 32.699056, 32.726333, 32.744944, 
    32.759056, 32.765917, 32.783278, 32.800722, 32.822444, 32.831833, 
    32.844333, 32.848639, 32.853528, 32.850778, 32.856417, 32.880083, 
    32.902083, 32.914194, 32.925611, 32.953889, 33.008833, 33.035889, 33.125, 
    33.127667, 33.165528, 33.209, 33.212083, 33.25425, 33.332139, 33.364139, 
    33.378389, 33.38425, 33.399528, 33.411667, 33.444861, 33.460778, 
    33.460028, 33.462611, 33.459278, 33.459056, 33.481972, 33.485333, 
    33.496417, 33.509583, 33.514167, 33.54175, 33.546611, 33.551556, 
    33.553028, 33.560528, 33.565667, 33.574889, 33.582306, 33.593, 33.605722, 
    33.619417, 33.645194, 33.677889, 33.70875, 33.729556, 33.734167, 
    33.732056, 33.736222, 33.738722, 33.734611, 33.734556, 33.737917, 
    33.739583, 33.742917, 33.75125, 33.762056, 33.763722, 33.759556, 
    33.759556, 33.762083, 33.759556, 33.765417, 33.758778, 33.753361, 
    33.749944, 33.738778, 33.737889, 33.740361, 33.742472, 33.750389, 
    33.744583, 33.744972, 33.752083, 33.749167, 33.740389, 33.744556, 
    33.750861, 33.755778, 33.759167, 33.760389, 33.757056, 33.762083, 
    33.752056, 33.755417, 33.75, 33.744583, 33.742917, 33.745389, 33.742889, 
    33.739583, 33.741222, 33.744139, 33.751222, 33.746694, 33.73125, 
    33.731667, 33.737889, 33.7325, 33.723333, 33.722083, 33.735806, 
    33.752889, 33.765417, 33.769611, 33.769556, 33.76625, 33.771667, 
    33.769583, 33.772944, 33.765417, 33.767083, 33.762889, 33.766222, 33.76, 
    33.754556, 33.759583, 33.754583, 33.755806, 33.767917, 33.766667, 
    33.757889, 33.754972, 33.756222, 33.7525, 33.749139, 33.7375, 33.721667, 
    33.720806, 33.715, 33.713694, 33.724583, 33.718278, 33.714111, 33.709972, 
    33.705444, 33.705417, 33.710417, 33.714556, 33.71875, 33.727889, 
    33.734611, 33.738694, 33.737083, 33.742917, 33.742917, 33.737028, 
    33.742056, 33.742056, 33.754139, 33.775806, 33.783694, 33.792472, 
    33.801278, 33.806667, 33.840833, 33.8475, 33.884167, 33.961667, 
    33.967889, 33.976667, 33.977472, 33.982056, 33.98375, 33.982472, 
    33.979972, 33.978306, 33.977472, 33.973333, 33.972472, 33.972056, 
    33.969139, 33.964556, 33.985806, 33.991639, 33.994972, 34, 34.006389, 
    34.006722, 34.011806, 34.02875, 34.033833, 34.037361, 34.039917, 
    34.036667, 34.039, 34.035472, 34.038083, 34.030639, 34.031444, 34.028833, 
    34.033222, 34.025694, 34.020583, 34.008611, 34.005667, 34.000167, 
    34.033083, 34.038167, 34.040583, 34.044694, 34.042194, 34.046444, 
    34.058778, 34.065861, 34.065056, 34.081556, 34.084056, 34.097556, 
    34.098333, 34.093222, 34.099167, 34.141583, 34.144194, 34.149694, 
    34.167472, 34.223222, 34.245861, 34.247333, 34.240222, 34.2445, 34.251, 
    34.251194, 34.261611, 34.273222, 34.272583, 34.277639, 34.282556, 
    34.290083, 34.302389, 34.319306, 34.317556, 34.354111, 34.354361, 
    34.371722, 34.375167, 34.371972, 34.381778, 34.386056, 34.393361, 
    34.395167, 34.414222, 34.411639, 34.418417, 34.420056, 34.415028, 
    34.415111, 34.411556, 34.407306, 34.402694, 34.400806, 34.395194, 
    34.394139, 34.394111, 34.401694, 34.416722, 34.414333, 34.403278, 
    34.408472, 34.406639, 34.416639, 34.431611, 34.434778, 34.43575, 
    34.44825, 34.449083, 34.460111, 34.461806, 34.457389, 34.462444, 
    34.46075, 34.463083, 34.459028, 34.459917, 34.469944, 34.473417, 
    34.46825, 34.470917, 34.4665, 34.46975, 34.465694, 34.461528, 34.458389, 
    34.454222, 34.452639, 34.449194, 34.451028, 34.441722, 34.448333, 
    34.448111, 34.474306, 34.480694, 34.487944, 34.49225, 34.49425, 
    34.512333, 34.523278, 34.539083, 34.54, 34.550611, 34.556611, 34.556944, 
    34.552278, 34.553444, 34.560556, 34.559389, 34.563694, 34.571528, 
    34.576556, 34.578944, 34.586083, 34.592444, 34.603722, 34.61125, 
    34.649778, 34.689472, 34.692417, 34.693194, 34.70725, 34.712917, 
    34.731611, 34.7385, 34.745111, 34.749528, 34.757833, 34.807639, 
    34.840694, 34.861556, 34.880722, 34.887917, 34.899972, 34.899861, 
    34.902583, 34.926222, 34.930361, 34.939333, 34.985833, 35.051306, 
    35.104028, 35.135139, 35.143833, 35.151361, 35.153028, 35.158111, 
    35.174556, 35.174167, 35.178889, 35.178111, 35.171556, 35.159306, 
    35.162444, 35.168028, 35.177889, 35.187139, 35.209, 35.213139, 35.216389, 
    35.219, 35.23125, 35.234417, 35.247778, 35.249806, 35.257083, 35.262278, 
    35.275028, 35.275472, 35.28125, 35.294639, 35.316528, 35.347972, 35.37, 
    35.368778, 35.344611, 35.326333, 35.314611, 35.319472, 35.323944, 
    35.332389, 35.332972, 35.338917, 35.342389, 35.340417, 35.342444, 
    35.371222, 35.372333, 35.367167, 35.368028, 35.372139, 35.373972, 
    35.381444, 35.397083, 35.43125, 35.447972, 35.44625, 35.451306, 
    35.458833, 35.460028, 35.483361, 35.489944, 35.50325, 35.509472, 
    35.551667, 35.560528, 35.575639, 35.582861, 35.592861, 35.600028, 
    35.605583, 35.636583, 35.642861, 35.640972, 35.635861, 35.634306, 
    35.650972, 35.652056, 35.654333, 35.663833, 35.666222, 35.667083, 
    35.664333, 35.692556, 35.714389, 35.720861, 35.727222, 35.737667, 
    35.745167, 35.749667, 35.755306, 35.759861, 35.769778, 35.783389, 
    35.805028, 35.810278, 35.815806, 35.821806, 35.855778, 35.858722, 
    35.870389, 35.88775, 35.896806, 35.918972, 35.923417, 35.9265, 35.930222, 
    35.933611, 35.950111, 35.97, 36, 36.014194, 36.0185, 36.018389, 
    36.021667, 36.041611, 36.048528, 36.052861, 36.06325, 36.070972, 
    36.086583, 36.101806, 36.119306, 36.126139, 36.161972, 36.174472, 36.195, 
    36.210028, 36.210139, 36.227, 36.227583, 36.233361, 36.231722, 36.234167, 
    36.238528, 36.247667, 36.259361, 36.276611, 36.279389, 36.28875, 
    36.301722, 36.304278, 36.308694, 36.308556, 36.313222, 36.337444, 
    36.356528, 36.3645, 36.373694, 36.381917, 36.392444, 36.397861, 
    36.402444, 36.417194, 36.425806, 36.448389, 36.460222, 36.469611, 
    36.488167, 36.491583, 36.498361, 36.504861, 36.5205, 36.525139, 
    36.521861, 36.525028, 36.526444, 36.535833, 36.539444, 36.552, 36.560972, 
    36.5605, 36.56425, 36.565028, 36.559222, 36.5685, 36.580472, 36.585, 
    36.584944, 36.608194, 36.611639, 36.611861, 36.626806, 36.629472, 
    36.636444, 36.639, 36.636611, 36.625111, 36.623167, 36.602556, 36.604194, 
    36.612417, 36.647917, 36.68075, 36.712611, 36.751806, 36.7525, 36.757056, 
    36.807444, 36.851361, 36.853639, 36.931556, 36.963361, 36.977528, 
    36.977222, 36.970694, 36.954194, 36.964222, 36.960194, 36.950028, 
    36.951639, 36.947417, 36.949306, 36.947444, 36.949167, 36.9525, 
    36.954806, 36.964917, 36.9665, 36.974667, 36.975833, 36.987361, 
    36.987389, 36.992389, 36.99925, 37.008722, 37.013722, 37.02375, 
    37.024556, 37.042472, 37.06, 37.095417, 37.107056, 37.117083, 37.116278, 
    37.110389, 37.116667, 37.119972, 37.136639, 37.144583, 37.150833, 
    37.161639, 37.171639, 37.182083, 37.18125, 37.191611, 37.196639, 37.22, 
    37.2275, 37.233306, 37.25, 37.248722, 37.2625, 37.265, 37.270833, 
    37.321611, 37.3575, 37.361639, 37.375, 37.391667, 37.407472, 37.434972, 
    37.456611, 37.486667, 37.502028, 37.502111, 37.499944, 37.494556, 
    37.494583, 37.502472, 37.505833, 37.521667, 37.534167, 37.551639, 
    37.564194, 37.571639, 37.588278, 37.594139, 37.597028, 37.595389, 
    37.601611, 37.605861, 37.610806, 37.619972, 37.630778, 37.649139, 
    37.694944, 37.725, 37.781611, 37.787889, 37.789583, 37.809556, 37.80625, 
    37.810389, 37.808722, 37.812083, 37.807889, 37.791667, 37.778333, 
    37.774111, 37.772472, 37.764139, 37.759972, 37.754167, 37.752444, 
    37.74875, 37.748333, 37.747944, 37.741611, 37.739972, 37.733722, 
    37.73375, 37.728306, 37.724167, 37.719167, 37.716222, 37.719611, 
    37.723722, 37.722056, 37.718306, 37.711611, 37.709139, 37.7075, 37.68, 
    37.677444, 37.671611, 37.67125, 37.665833, 37.665417, 37.661611, 
    37.659972, 37.655778, 37.650806, 37.647917, 37.642472, 37.635833, 
    37.632917, 37.629583, 37.6275, 37.621639, 37.614139, 37.608306, 
    37.612111, 37.606639, 37.592889, 37.590361, 37.592056, 37.587917, 
    37.592083, 37.590389, 37.581611, 37.575389, 37.575389, 37.571194, 
    37.57625, 37.570389, 37.572889, 37.57125, 37.5625, 37.552083, 37.55375, 
    37.551667, 37.545806, 37.530444, 37.545444, 37.5425, 37.534556, 
    37.542083, 37.536694, 37.53, 37.516639, 37.50375, 37.513333, 37.5175, 
    37.5225, 37.524583, 37.518778, 37.521194, 37.510806, 37.504944, 
    37.497917, 37.498694, 37.502083, 37.507889, 37.507944, 37.504167, 
    37.469972, 37.46375, 37.463722, 37.4575, 37.45875, 37.451222, 37.452056, 
    37.447917, 37.450417, 37.450417, 37.445417, 37.45125, 37.449611, 
    37.453333, 37.459583, 37.461222, 37.455417, 37.46125, 37.464167, 
    37.46875, 37.468722, 37.464583, 37.49, 37.492889, 37.492083, 37.49625, 
    37.497028, 37.50125, 37.505389, 37.498694, 37.499139, 37.505806, 
    37.521667, 37.545833, 37.555806, 37.564139, 37.563333, 37.585806, 
    37.606639, 37.615, 37.6175, 37.625833, 37.629972, 37.639139, 37.645, 
    37.648361, 37.67, 37.695833, 37.697083, 37.692056, 37.697917, 37.697444, 
    37.7, 37.704111, 37.702917, 37.706667, 37.712083, 37.710417, 37.699583, 
    37.717917, 37.722083, 37.721611, 37.743333, 37.749556, 37.74875, 
    37.750417, 37.762056, 37.767861, 37.767028, 37.769556, 37.766667, 
    37.763722, 37.764556, 37.770389, 37.769556, 37.773333, 37.780417, 
    37.780417, 37.77625, 37.776222, 37.77875, 37.781639, 37.7975, 37.802056, 
    37.801222, 37.804139, 37.807083, 37.80375, 37.805806, 37.810389, 
    37.812083, 37.819972, 37.819583, 37.824167, 37.831639, 37.836222, 
    37.836639, 37.838778, 37.840806, 37.864139, 37.865417, 37.859556, 37.865, 
    37.865389, 37.868306, 37.867861, 37.871667, 37.874556, 37.871222, 
    37.871639, 37.888306, 37.89, 37.892056, 37.894972, 37.897056, 37.895361, 
    37.901667, 37.903306, 37.909583, 37.907889, 37.9125, 37.914583, 
    37.908694, 37.907889, 37.919111, 37.923722, 37.923306, 37.92, 37.905389, 
    37.90375, 37.910389, 37.905389, 37.919972, 37.929583, 37.932889, 
    37.943306, 37.946667, 37.951639, 37.966278, 37.962917, 37.957083, 
    37.952889, 37.955, 37.958722, 37.9575, 37.969556, 37.970417, 37.977083, 
    37.975417, 37.978306, 37.993333, 37.997472, 38.014833, 38.004083, 
    38.004167, 38.014083, 38.014111, 38.020417, 38.02475, 38.025806, 
    38.038917, 38.04025, 38.050361, 38.053972, 38.060833, 38.065472, 
    38.073083, 38.098917, 38.115778, 38.127306, 38.128278, 38.138889, 
    38.146361, 38.154917, 38.143861, 38.13725, 38.114028, 38.116111, 
    38.120583, 38.116472, 38.110944, 38.119855, 38.129139, 38.113333, 
    38.10575, 38.093222, 38.0915, 38.081417, 38.06675, 38.035056, 38.02475, 
    38.017417, 38.0165, 38.009139, 38.00575, 37.988333, 37.980361, 37.984583, 
    37.982889, 37.972889, 37.972917, 37.974972, 37.975444, 37.969972, 
    37.966667, 37.949194, 37.947083, 37.942056, 37.937056, 37.943722, 
    37.941639, 37.937944, 37.929167, 37.921222, 37.92125, 37.916694, 
    37.909167, 37.908333, 37.904556, 37.895389, 37.894583, 37.881667, 
    37.87125, 37.8725, 37.862056, 37.871639, 37.884583, 37.89375, 37.895, 
    37.890806, 37.877861, 37.883694, 37.88875, 37.887056, 37.89375, 
    37.892056, 37.885806, 37.882889, 37.882917, 37.876194, 37.870833, 
    37.86625, 37.859194, 37.849111, 37.839111, 37.833278, 37.833778, 
    37.825389, 37.826222, 37.820389, 37.824583, 37.825361, 37.819167, 
    37.815444, 37.824111, 37.828361, 37.832028, 37.835389, 37.841639, 
    37.843722, 37.85375, 37.853722, 37.859583, 37.859556, 37.875417, 
    37.877083, 37.881222, 37.900389, 37.905417, 37.907083, 37.893722, 
    37.902889, 37.926222, 37.93375, 37.936222, 37.94375, 37.942889, 
    37.947083, 37.947083, 37.967472, 37.981222, 37.986222, 38.004972, 
    38.019028, 38.028278, 38.029111, 38.034028, 38.034944, 38.031583, 
    38.030833, 38.02575, 38.013278, 37.999139, 37.99375, 37.989556, 
    37.994556, 37.992694, 37.994417, 38.001778, 38.004139, 38.011, 38.065806, 
    38.129, 38.151667, 38.176278, 38.182389, 38.185667, 38.199389, 38.213972, 
    38.221667, 38.237222, 38.240611, 38.238139, 38.230806, 38.236583, 
    38.251528, 38.269056, 38.2715, 38.292111, 38.310083, 38.311694, 
    38.306583, 38.2995, 38.298222, 38.301778, 38.315278, 38.322778, 
    38.323222, 38.339444, 38.363472, 38.3895, 38.395611, 38.410472, 
    38.430667, 38.452972, 38.455889, 38.461472, 38.464778, 38.467917, 
    38.474917, 38.494028, 38.5025, 38.510028, 38.512472, 38.510972, 
    38.532444, 38.53175, 38.539806, 38.547694, 38.555778, 38.559889, 
    38.566472, 38.565944, 38.573194, 38.58325, 38.590278, 38.597306, 
    38.597444, 38.604278, 38.609083, 38.610306, 38.614139, 38.616972, 
    38.630722, 38.635417, 38.63825, 38.641111, 38.64625, 38.648889, 
    38.649194, 38.655306, 38.659278, 38.674556, 38.679611, 38.683083, 
    38.689722, 38.704167, 38.706139, 38.718111, 38.726889, 38.737944, 
    38.741778, 38.751611, 38.756417, 38.759917, 38.766972, 38.777917, 
    38.784861, 38.790417, 38.80075, 38.800806, 38.809167, 38.807778, 
    38.811139, 38.812306, 38.819944, 38.826667, 38.831056, 38.843333, 
    38.843583, 38.865389, 38.874972, 38.881861, 38.893028, 38.90025, 
    38.91175, 38.916, 38.917694, 38.921556, 38.936722, 38.956139, 38.957889, 
    38.99925, 39.0025, 39.035139, 39.036722, 39.041972, 39.044472, 39.061389, 
    39.088389, 39.104167, 39.108417, 39.115444, 39.12275, 39.134111, 
    39.14075, 39.138833, 39.153361, 39.157444, 39.173472, 39.186889, 
    39.192667, 39.192, 39.198389, 39.201222, 39.212722, 39.215222, 39.223583, 
    39.227472, 39.231583, 39.239056, 39.252194, 39.258222, 39.271333, 
    39.269972, 39.279417, 39.29075, 39.291139, 39.298056, 39.300139, 
    39.301639, 39.299167, 39.306389, 39.311194, 39.313889, 39.318306, 
    39.323222, 39.327361, 39.32675, 39.333167, 39.33775, 39.348389, 
    39.354361, 39.361278, 39.361111, 39.366917, 39.376833, 39.3785, 
    39.388361, 39.405472, 39.416806, 39.423167, 39.428278, 39.430333, 
    39.438583, 39.441222, 39.452083, 39.473333, 39.485694, 39.490083, 
    39.489972, 39.504278, 39.558083, 39.568194, 39.572722, 39.582333, 
    39.591333, 39.601944, 39.611833, 39.620528, 39.625361, 39.65025, 
    39.659556, 39.665833, 39.687389, 39.708444, 39.723389, 39.734556, 
    39.738472, 39.740556, 39.754583, 39.792972, 39.805333, 39.830139, 
    39.845222, 39.85925, 39.907972, 39.911139, 39.922167, 39.960306, 
    39.967528, 39.984778, 39.988556, 39.996972, 40.015, 40.025056, 40.021639, 
    40.02475, 40.031778, 40.064167, 40.078694, 40.103639, 40.115722, 
    40.123333, 40.129972, 40.1565, 40.174333, 40.183417, 40.198722, 
    40.204111, 40.22975, 40.238278, 40.249861, 40.260361, 40.28325, 
    40.316389, 40.324028, 40.338361, 40.348389, 40.374833, 40.388194, 
    40.402528, 40.409722, 40.441667, 40.44975, 40.4715, 40.494944, 40.501861, 
    40.513083, 40.534139, 40.557444, 40.62625, 40.629194, 40.629639, 
    40.634917, 40.630611, 40.635806, 40.709222, 40.759333, 40.749833, 
    40.746278, 40.742861, 40.745028, 40.750639, 40.757667, 40.771889, 
    40.77425, 40.772778, 40.797056, 40.806583, 40.814889, 40.813722, 
    40.783861, 40.7685, 40.760028, 40.760333, 40.7685, 40.785028, 40.863222, 
    40.926861, 40.995306, 41.028861, 41.046583, 41.057472, 41.058278, 
    41.052778, 41.052472, 41.063389, 41.071972, 41.077861, 41.087139, 41.089, 
    41.103278, 41.106361, 41.117333, 41.131083, 41.140694, 41.144806, 
    41.143111, 41.147361, 41.227861, 41.234833, 41.2395, 41.243472, 
    41.265167, 41.319, 41.324194, 41.378417, 41.444694, 41.478222, 41.518972, 
    41.544056, 41.5535, 41.567667, 41.584917, 41.594917, 41.601694, 
    41.615056, 41.641778, 41.656556, 41.673472, 41.680194, 41.687528, 
    41.703278, 41.723111, 41.739417, 41.745833, 41.750028, 41.750833, 
    41.748472, 41.74425, 41.744278, 41.750083, 41.770917, 41.770611, 
    41.773167, 41.783917, 41.798167, 41.821639, 41.895972, 41.942861, 
    41.949944, 41.981222, 41.997917, 42.008583, 42.013444, 42.022361, 
    42.028056, 42.044361, 42.042306, 42.044694, 42.0415, 42.047389, 
    42.050222, 42.062472, 42.067361, 42.082333, 42.087639, 42.098833, 
    42.098139, 42.102194, 42.110972, 42.118111, 42.12175, 42.136361, 
    42.142361, 42.143389, 42.156583, 42.161306, 42.16925, 42.181028, 
    42.182861, 42.194167, 42.196639, 42.206833, 42.208778, 42.222333, 
    42.252278, 42.292139, 42.320639, 42.318417, 42.32925, 42.334806, 
    42.372972, 42.404194, 42.419111, 42.426, 42.428278, 42.427583, 42.420167, 
    42.438472, 42.459139, 42.463194, 42.466389, 42.474806, 42.476694, 
    42.490167, 42.496694, 42.528194, 42.569083, 42.575389, 42.577417, 42.583, 
    42.591333, 42.590722, 42.596028, 42.597194, 42.625389, 42.629111, 
    42.635583, 42.641472, 42.643611, 42.646556, 42.649972, 42.661528, 
    42.674694, 42.687389, 42.691694, 42.73325, 42.741722, 42.739167, 
    42.734167, 42.73525, 42.792417, 42.813333, 42.830806, 42.834111, 
    42.839167, 42.843222, 42.839889, 42.845194, 42.868444, 42.876389, 
    42.884028, 42.923722, 43.023611, 43.064667, 43.098694, 43.115167, 
    43.129667, 43.186778, 43.213, 43.230417, 43.269972, 43.277806, 43.291056, 
    43.303444, 43.301806, 43.306333, 43.324167, 43.330778, 43.335083, 
    43.341611, 43.34075, 43.344944, 43.344917, 43.352333, 43.349889, 
    43.351528, 43.345083, 43.340889, 43.359139, 43.364806, 43.364361, 
    43.375278, 43.383889, 43.397889, 43.415111, 43.418833, 43.425917, 
    43.426583, 43.423444, 43.38325, 43.374306, 43.372444, 43.383444, 
    43.388111, 43.388306, 43.395556, 43.401, 43.403528, 43.406806, 43.412389, 
    43.421556, 43.420889, 43.432167, 43.43325, 43.43625, 43.447889, 
    43.451111, 43.462306, 43.467056, 43.468139, 43.455944, 43.450667, 
    43.454694, 43.431722, 43.430806, 43.434167, 43.426, 43.424972, 43.421583, 
    43.412333, 43.400528, 43.382361, 43.363889, 43.356, 43.357472, 43.410389, 
    43.483833, 43.564972, 43.668667, 43.671861, 43.67975, 43.682333, 
    43.675833, 43.673889, 43.707583, 43.814083, 43.959194, 44.015417, 
    44.005389, 44.008306, 44.021667, 44.102472, 44.116667, 44.120778, 
    44.134167, 44.138333, 44.144167, 44.162472, 44.217472, 44.232444, 
    44.246639, 44.265, 44.273333, 44.281667, 44.294167, 44.304167, 44.307472, 
    44.31, 44.314944, 44.357472, 44.419111, 44.423694, 44.435417, 44.433278, 
    44.431194, 44.433778, 44.428722, 44.433722, 44.431222, 44.4375, 
    44.442917, 44.442056, 44.450389, 44.434556, 44.42375, 44.425833, 
    44.460833, 44.4975, 44.521639, 44.580833, 44.614167, 44.620389, 
    44.626222, 44.622472, 44.618306, 44.612917, 44.615417, 44.604167, 
    44.602889, 44.62, 44.62625, 44.62875, 44.6225, 44.622083, 44.632083, 
    44.621222, 44.666611, 44.672944, 44.672889, 44.6775, 44.679556, 
    44.677861, 44.682472, 44.732472, 44.741611, 44.746639, 44.767472, 
    44.771639, 44.786639, 44.789139, 44.790806, 44.798361, 44.804167, 
    44.8125, 44.8175, 44.820778, 44.826694, 44.832083, 44.831639, 44.849972, 
    44.927083, 44.892056, 44.897472, 44.909167, 44.915806, 44.926639, 
    44.929167, 44.95, 45.011389, 45.029778, 45.039444, 45.047389, 45.048278, 
    45.052306, 45.053778, 45.060611, 45.070556, 45.077056, 45.083444, 
    45.095333, 45.153528, 45.160667, 45.163083, 45.213222, 45.216861, 
    45.217444, 45.226833, 45.268778, 45.274528, 45.277639, 45.278361, 
    45.307111, 45.335028, 45.337833, 45.336528, 45.339972, 45.343556, 
    45.342333, 45.345028, 45.348278, 45.356167, 45.415972, 45.4155, 
    45.391417, 45.375306, 45.374861, 45.385778, 45.394472, 45.402861, 
    45.42625, 45.444, 45.463111, 45.480917, 45.489167, 45.498417, 45.511833, 
    45.504583, 45.507944, 45.505639, 45.494056, 45.472583, 45.482639, 
    45.483222, 45.488639, 45.490139, 45.498611, 45.502889, 45.501056, 
    45.505056, 45.509278, 45.51775, 45.527278, 45.535, 45.547556, 45.560806, 
    45.561194, 45.554667, 45.557472, 45.552778, 45.556861, 45.559306, 
    45.567722, 45.571278, 45.632333, 45.652222, 45.657056, 45.669944, 
    45.68975, 45.691833, 45.690361, 45.695611, 45.696222, 45.700361, 
    45.700556, 45.706917, 45.707528, 45.696861, 45.69175, 45.682, 45.670833, 
    45.658444, 45.661833, 45.704306, 45.731361, 45.742861, 45.763389, 
    45.760944, 45.767306, 45.782306, 45.803972, 45.814917, 45.843583, 
    45.880361, 45.886083, 45.893889, 45.907306, 45.914833, 45.91775, 
    45.929333, 45.937556, 45.947611, 45.95675, 45.971778, 45.979722, 
    46.009972, 46.014972, 46.018333, 46.074972, 46.125833, 46.205833, 
    46.224361, 46.226694, 46.229917, 46.233389, 46.233417, 46.229583, 
    46.225833, 46.22625, 46.222111, 46.208694, 46.212083, 46.207944, 
    46.203722, 46.185417, 46.167861, 46.165361, 46.160444, 46.15125, 
    46.167056, 46.164528, 46.170389, 46.152472, 46.150389, 46.16, 46.169556, 
    46.172917, 46.171222, 46.180417, 46.190417, 46.194583, 46.192028, 
    46.198722, 46.19625, 46.197917, 46.2025, 46.210389, 46.213722, 46.204139, 
    46.195833, 46.19375, 46.171222, 46.171611, 46.172083, 46.174556, 
    46.17375, 46.17125, 46.172083, 46.177083, 46.185361, 46.187083, 46.1875, 
    46.195417, 46.191222, 46.187056, 46.18875, 46.185361, 46.189972, 
    46.198333, 46.203278, 46.204972, 46.219583, 46.22625, 46.2325, 46.230806, 
    46.237056, 46.234556, 46.228306, 46.214583, 46.202056, 46.210778, 
    46.244167, 46.259583, 46.267889, 46.27375, 46.273722, 46.267056, 
    46.269583, 46.267056, 46.264583, 46.260389, 46.262056, 46.259556, 
    46.260444, 46.264556, 46.267056, 46.276667, 46.286694, 46.296667, 
    46.300806, 46.307444, 46.305417, 46.312056, 46.311667, 46.307444, 
    46.302056, 46.300806, 46.288722, 46.292083, 46.274528, 46.275444, 
    46.282917, 46.284556, 46.270389, 46.268722, 46.262861, 46.26125, 
    46.256611, 46.249583, 46.247917, 46.242056, 46.241222, 46.246222, 
    46.252056, 46.261278, 46.269556, 46.294139, 46.302944, 46.312917, 
    46.313889, 46.306722, 46.305778, 46.300222, 46.282833, 46.276389, 
    46.271694, 46.267694, 46.267611, 46.274083, 46.27425, 46.278472, 
    46.264194, 46.270639, 46.282444, 46.29275, 46.297306, 46.301889, 
    46.308111, 46.345611, 46.483139, 46.636306, 46.642444, 46.644222, 
    46.632944, 46.6275, 46.629306, 46.624139, 46.638722, 46.624528, 
    46.599667, 46.591028, 46.580833, 46.511889, 46.506778, 46.493833, 
    46.454167, 46.434861, 46.397444, 46.391139, 46.381333, 46.376028, 
    46.377889, 46.374556, 46.379528, 46.384556, 46.380389, 46.385417, 
    46.370778, 46.372028, 46.369611, 46.374139, 46.378333, 46.403306, 
    46.404556, 46.414139, 46.421667, 46.431667, 46.440806, 46.452528, 
    46.460444, 46.451667, 46.436667, 46.432889, 46.42875, 46.429556, 
    46.432472, 46.434556, 46.439944, 46.452472, 46.465389, 46.46625, 
    46.474139, 46.488306, 46.496694, 46.508278, 46.512028, 46.514556, 
    46.505833, 46.5125, 46.515, 46.53, 46.540833, 46.550417, 46.552056, 
    46.569111, 46.577472, 46.591667, 46.603306, 46.618306, 46.6375, 
    46.637083, 46.621222, 46.614611, 46.612889, 46.616278, 46.624194, 
    46.630389, 46.631639, 46.635417, 46.632056, 46.636639, 46.64375, 
    46.652444, 46.668333, 46.673778, 46.673694, 46.679583, 46.680361, 
    46.702889, 46.702056, 46.688722, 46.687917, 46.690833, 46.702444, 
    46.707056, 46.710417, 46.705833, 46.704556, 46.707472, 46.71625, 
    46.712056, 46.714167, 46.719583, 46.719528, 46.728722, 46.730389, 
    46.740389, 46.739556, 46.750389, 46.747083, 46.750389, 46.742917, 
    46.738306, 46.728306, 46.724583, 46.724583, 46.73875, 46.726639, 
    46.724139, 46.714194, 46.714972, 46.707917, 46.703722, 46.702889, 
    46.707083, 46.707833, 46.719056, 46.716611, 46.720667, 46.713917, 
    46.71325, 46.727667, 46.731028, 46.782167, 46.823111, 46.883028, 
    46.905528, 46.904972, 46.914056, 46.915, 46.907444, 46.904167, 46.894806, 
    46.881306, 46.88075, 46.869083, 46.865861, 46.8625, 46.864111, 46.858333, 
    46.857167, 46.859833, 46.864194, 46.861639, 46.863667, 46.877472, 
    46.890028, 46.897444, 46.902444, 46.905833, 46.903278, 46.910083, 
    46.914111, 46.914667, 46.909778, 46.924583, 46.922917, 46.931222, 
    46.942083, 46.952889, 46.957889, 46.971667, 46.97375, 46.96125, 
    46.970417, 46.96875, 46.971222, 46.972083, 46.968694, 46.971639, 
    46.97375, 46.975417, 46.977472, 46.982889, 46.980361, 46.984111, 
    46.993528, 46.997, 47.004, 47.008639, 47.015222, 47.029417, 47.034444, 
    47.032694, 47.037583, 47.03325, 47.033722, 47.040361, 47.041194, 
    47.032417, 47.021111, 47.008667, 47, 46.974556, 46.956361, 46.963611, 
    46.961778, 46.950194, 46.945806, 46.946444, 46.940778, 46.932639, 
    46.928306, 46.927333, 46.993056, 47.098389, 47.124972, 47.127333, 
    47.14375, 47.208194, 47.290917, 47.30275, 47.302861, 47.299361, 
    47.301917, 47.346639, 47.347917, 47.350194, 47.357444, 47.385444, 
    47.406556, 47.43025, 47.436528, 47.437556, 47.444833, 47.449556, 
    47.458778, 47.462139, 47.4645, 47.500556, 47.542778, 47.539194, 
    47.544639, 47.649917, 47.688611, 47.736167, 47.748056, 47.748778, 
    47.754722, 47.764694, 47.765528, 47.769444, 47.771472, 47.818472, 
    47.817917, 47.823111, 47.820361, 47.831028, 47.832972, 47.841667, 
    47.844139, 47.848722, 47.854444, 47.8655, 47.864972, 47.872778, 
    47.877167, 47.869778, 47.871194, 47.878028, 47.89125, 47.899694, 47.9085, 
    47.917111, 47.909056, 47.909361, 47.913444, 47.923694, 47.942222, 
    47.944611, 47.956111, 47.961, 47.9655, 47.969222, 47.981028, 48, 
    48.009167, 48.021667, 48.037472, 48.070778, 48.085833, 48.098306, 
    48.100806, 48.116639, 48.124972, 48.133306, 48.141639, 48.154194, 
    48.158722, 48.163306, 48.169556, 48.172861, 48.182056, 48.184556, 
    48.193333, 48.219944, 48.239139, 48.247889, 48.256639, 48.274972, 
    48.290806, 48.294167, 48.297917, 48.296194, 48.3, 48.315806, 48.319972, 
    48.325, 48.331667, 48.342472, 48.344583, 48.343722, 48.33875, 48.339611, 
    48.350417, 48.354139, 48.359972, 48.367083, 48.369972, 48.381667, 
    48.390417, 48.387028, 48.391222, 48.390389, 48.393694, 48.389528, 
    48.39125, 48.388722, 48.383278, 48.367917, 48.367028, 48.374583, 
    48.371194, 48.366194, 48.367889, 48.350361, 48.349528, 48.345389, 
    48.332889, 48.317889, 48.30875, 48.303722, 48.288722, 48.284611, 
    48.287917, 48.27625, 48.269556, 48.263306, 48.262889, 48.260389, 
    48.258722, 48.255361, 48.256222, 48.267111, 48.252889, 48.243694, 
    48.228722, 48.220417, 48.22125, 48.21875, 48.206611, 48.204583, 
    48.209583, 48.200361, 48.190361, 48.177056, 48.174528, 48.172056, 
    48.172917, 48.165333, 48.165333, 48.1695, 48.167, 48.167806, 48.162833, 
    48.160333, 48.161167, 48.156194, 48.157, 48.162806, 48.157, 48.156167, 
    48.157, 48.162861, 48.161222, 48.165333, 48.165333, 48.161167, 48.1595, 
    48.164889, 48.168639, 48.168667, 48.166167, 48.163667, 48.157, 48.150722, 
    48.146194, 48.139472, 48.136194, 48.152, 48.152, 48.136167, 48.132861, 
    48.135361, 48.143694, 48.142806, 48.139111, 48.137, 48.140333, 48.138694, 
    48.134944, 48.128694, 48.126167, 48.122806, 48.124556, 48.119472, 
    48.117028, 48.121194, 48.116139, 48.115333, 48.118667, 48.114528, 
    48.1145, 48.115333, 48.122833, 48.117833, 48.116167, 48.126167, 
    48.141194, 48.156194, 48.175361, 48.186167, 48.182028, 48.175333, 
    48.157028, 48.171611, 48.174528, 48.1695, 48.175333, 48.171194, 
    48.148222, 48.152, 48.160333, 48.152861, 48.151167, 48.153667, 48.153694, 
    48.126194, 48.121167, 48.08575, 48.082833, 48.091972, 48.08325, 
    48.081972, 48.085306, 48.082389, 48.064111, 48.057417, 48.038694, 
    48.030361, 48.024528, 48.026167, 48.029083, 48.044917, 48.052389, 
    48.061611, 48.069944, 48.078694, 48.082, 48.079472, 48.082, 48.098667, 
    48.096194, 48.074944, 48.063278, 48.057056, 48.047, 48.019917, 48.0045, 
    47.993722, 47.991278, 47.996222, 48.008694, 48.042444, 48.048667, 
    48.055333, 48.067, 48.076222, 48.076556, 48.089917, 48.10575, 48.122, 
    48.137861, 48.135333, 48.143667, 48.145306, 48.132417, 48.116611, 
    48.108667, 48.105361, 48.092028, 48.08575, 48.080361, 48.065333, 
    48.057417, 48.047417, 48.040333, 48.037, 48.027833, 48.033694, 48.025722, 
    48.026139, 48.023222, 48.024083, 48.019111, 47.999167, 47.991667, 
    47.975417, 47.97375, 47.969972, 47.958306, 47.942444, 47.924167, 
    47.920389, 47.923722, 47.920389, 47.916611, 47.91625, 47.918778, 
    47.915389, 47.917056, 47.927111, 47.932083, 47.923333, 47.905806, 
    47.894583, 47.89125, 47.891222, 47.8875, 47.877917, 47.88625, 47.868306, 
    47.863722, 47.867917, 47.868722, 47.862472, 47.851667, 47.831694, 
    47.825389, 47.812056, 47.809583, 47.803306, 47.793306, 47.783333, 
    47.776639, 47.773333, 47.768306, 47.759167, 47.745806, 47.742056, 
    47.723278, 47.704944, 47.692472, 47.688778, 47.685389, 47.681222, 
    47.691667, 47.71, 47.716667, 47.726667, 47.731667, 47.745778, 47.769139, 
    47.788306, 47.794139, 47.805861, 47.810833, 47.821639, 47.845389, 
    47.8375, 47.822472, 47.810028, 47.792472, 47.779528, 47.779556, 
    47.783333, 47.805833, 47.824111, 47.827056, 47.810833, 47.7925, 
    47.769972, 47.760806, 47.739972, 47.73625, 47.745417, 47.744556, 47.7325, 
    47.730389, 47.731667, 47.712472, 47.700806, 47.689167, 47.666667, 
    47.664139, 47.645806, 47.646278, 47.650389, 47.630389, 47.627889, 
    47.624583, 47.61875, 47.614583, 47.606639, 47.604139, 47.601222, 
    47.581528, 47.563139, 47.551917, 47.550778, 47.545639, 47.52925, 
    47.503972, 47.465111, 47.461611, 47.463139, 47.452528, 47.414778, 
    47.408278, 47.376194, 47.371556, 47.362472, 47.3535, 47.344778, 
    47.341611, 47.346, 47.346, 47.359278, 47.359278, 47.355083, 47.350833, 
    47.35275, 47.357611, 47.361611, 47.370806, 47.37, 47.375917, 47.373167, 
    47.373944, 47.391306, 47.449806, 47.455639, 47.453917, 47.458333, 
    47.465917, 47.489194, 47.502972, 47.510917, 47.529306, 47.544528, 
    47.558778, 47.561667, 47.566639, 47.568306, 47.58625, 47.587028, 
    47.59875, 47.61, 47.617472, 47.623694, 47.625417, 47.634583, 47.630389, 
    47.652083, 47.655444, 47.654167, 47.642472, 47.638694, 47.654583, 
    47.657917, 47.671222, 47.682472, 47.719972, 47.738333, 47.740833, 
    47.770389, 47.779972, 47.802917, 47.812889, 47.817083, 47.829556, 
    47.837056, 47.837028, 47.857889, 47.85875, 47.834139, 47.815389, 
    47.823278, 47.839972, 47.854972, 47.873306, 47.900833, 47.906639, 
    47.9125, 47.920417, 47.924583, 47.929167, 47.931639, 47.941222, 
    47.942028, 47.9275, 47.922083, 47.92125, 47.913722, 47.912472, 47.9025, 
    47.879972, 47.865, 47.855778, 47.834139, 47.826222, 47.817917, 47.813333, 
    47.797056, 47.796639, 47.790389, 47.780833, 47.769944, 47.766667, 
    47.756667, 47.747944, 47.743722, 47.746222, 47.731639, 47.703306, 
    47.697472, 47.690417, 47.69625, 47.705, 47.712056, 47.707917, 47.714139, 
    47.7175, 47.727056, 47.745417, 47.744167, 47.725, 47.72, 47.713694, 
    47.715389, 47.707889, 47.713306, 47.700806, 47.700389, 47.703306, 
    47.707083, 47.705389, 47.700861, 47.693306, 47.664167, 47.651667, 
    47.639556, 47.637528, 47.603306, 47.593306, 47.574528, 47.567889, 
    47.56875, 47.58125, 47.58375, 47.604139, 47.615417, 47.622472, 47.6375, 
    47.648722, 47.64875, 47.643306, 47.635, 47.614167, 47.60375, 47.60375, 
    47.610417, 47.608333, 47.599139, 47.5975, 47.593306, 47.584972, 
    47.576667, 47.585, 47.594139, 47.596194, 47.593722, 47.604556, 47.599972, 
    47.584972, 47.580389, 47.58875, 47.578722, 47.57875, 47.570833, 
    47.560389, 47.554583, 47.547083, 47.536194, 47.529167, 47.527889, 
    47.532083, 47.540389, 47.53875, 47.544611, 47.543778, 47.548722, 
    47.548722, 47.568778, 47.582917, 47.590417, 47.588333, 47.576667, 47.57, 
    47.569556, 47.565806, 47.558306, 47.545, 47.524944, 47.524583, 47.519528, 
    47.519583, 47.511667, 47.485833, 47.475833, 47.469972, 47.449139, 
    47.426639, 47.4075, 47.397444, 47.3875, 47.375, 47.326222, 47.340444, 
    47.336639, 47.328306, 47.313306, 47.288306, 47.275, 47.2585, 47.25, 
    47.281667, 47.294972, 47.315, 47.319583, 47.317889, 47.307083, 47.307056, 
    47.284556, 47.273722, 47.256194, 47.261639, 47.270417, 47.262944, 
    47.269972, 47.270417, 47.272472, 47.277028, 47.274167, 47.279167, 
    47.283722, 47.278778, 47.280806, 47.283778, 47.290417, 47.297917, 
    47.297111, 47.300417, 47.30625, 47.308778, 47.320389, 47.322056, 
    47.329583, 47.327917, 47.335417, 47.342917, 47.348306, 47.354167, 
    47.399167, 47.4175, 47.442056, 47.447083, 47.450833, 47.459944, 
    47.469167, 47.483278, 47.49, 47.502917, 47.515833, 47.524139, 47.529944, 
    47.535806, 47.555833, 47.569944, 47.575833, 47.596194, 47.585389, 
    47.585389, 47.57625, 47.587944, 47.59125, 47.57375, 47.6, 47.608722, 
    47.627917, 47.626222, 47.632083, 47.63125, 47.637083, 47.65375, 
    47.660806, 47.672917, 47.6675, 47.675, 47.684194, 47.695, 47.707028, 
    47.718306, 47.732472, 47.7475, 47.758333, 47.772472, 47.779167, 
    47.786667, 47.806694, 47.811278, 47.842917, 47.850806, 47.871639, 
    47.8825, 47.901667, 47.915806, 47.925861, 47.939111, 47.950389, 
    47.957889, 47.959556, 47.967083, 47.981667, 47.988333, 47.986194, 
    47.989139, 47.992111, 47.996639, 48, 48.005722, 48.012444, 48.017028, 
    48.019556, 48.018667, 48.012861, 48.002833, 48.00575, 48.014111, 
    48.023639, 48.021167, 48.022417, 48.030361, 48.034083, 48.037056, 
    48.040722, 48.0445, 48.045333, 48.038722, 48.030306, 48.032028, 
    48.045333, 48.052, 48.056167, 48.058667, 48.054056, 48.051194, 48.05325, 
    48.062833, 48.065361, 48.062861, 48.071194, 48.080333, 48.092806, 
    48.099083, 48.11075, 48.12325, 48.132444, 48.13575, 48.140722, 48.150778, 
    48.164944, 48.187417, 48.188278, 48.192444, 48.194944, 48.214083, 
    48.222028, 48.226583, 48.232, 48.2245, 48.234528, 48.2295, 48.226167, 
    48.227833, 48.235333, 48.232861, 48.227389, 48.219111, 48.215333, 
    48.214944, 48.209111, 48.193667, 48.193694, 48.199528, 48.205333, 
    48.195333, 48.19575, 48.189917, 48.177417, 48.172417, 48.167444, 
    48.162444, 48.150778, 48.144556, 48.129472, 48.126139, 48.117028, 
    48.114528, 48.093639, 48.067389, 48.063222, 48.057, 48.057, 48.063667, 
    48.078278, 48.085333, 48.091972, 48.103694, 48.106972, 48.130361, 
    48.128667, 48.121167, 48.121139, 48.128667, 48.132028, 48.166583, 
    48.170778, 48.183278, 48.19325, 48.205778, 48.247417, 48.252028, 
    48.258694, 48.253694, 48.252833, 48.258278, 48.270333, 48.271194, 
    48.260361, 48.258694, 48.2545, 48.247861, 48.254083, 48.256583, 48.26825, 
    48.266611, 48.260333, 48.272444, 48.280806, 48.292417, 48.301556, 
    48.299889, 48.314917, 48.308694, 48.31325, 48.317861, 48.314472, 
    48.322833, 48.327, 48.331222, 48.329528, 48.336194, 48.336194, 48.341139, 
    48.358278, 48.361972, 48.357833, 48.360361, 48.358694, 48.369528, 
    48.371194, 48.378694, 48.372861, 48.374472, 48.381167, 48.379944, 
    48.372444, 48.372, 48.38325, 48.390361, 48.383278, 48.371167, 48.372861, 
    48.375333, 48.374528, 48.391611, 48.406583, 48.419111, 48.41825, 
    48.421167, 48.422444, 48.44325, 48.452833, 48.444472, 48.444528, 
    48.447056, 48.445361, 48.429083, 48.422861, 48.423694, 48.413667, 
    48.412833, 48.415361, 48.4095, 48.410361, 48.407861, 48.412444, 
    48.414917, 48.417833, 48.4145, 48.420333, 48.426611, 48.443278, 
    48.443667, 48.449056, 48.452444, 48.455778, 48.472417, 48.47575, 
    48.484083, 48.4895, 48.494528, 48.490306, 48.490361, 48.49825, 48.509528, 
    48.505361, 48.522833, 48.522861, 48.519111, 48.511972, 48.516194, 
    48.513222, 48.486611, 48.482417, 48.479917, 48.465306, 48.463667, 
    48.466583, 48.47825, 48.48575, 48.492417, 48.490306, 48.492444, 
    48.500333, 48.501139, 48.47075, 48.459528, 48.459528, 48.452833, 
    48.463667, 48.458694, 48.457861, 48.461167, 48.458694, 48.458694, 48.452, 
    48.463694, 48.466194, 48.459889, 48.465722, 48.469083, 48.474917, 
    48.488278, 48.51325, 48.519917, 48.520778, 48.534917, 48.541583, 
    48.559083, 48.563667, 48.565333, 48.5745, 48.573667, 48.579917, 
    48.582389, 48.589528, 48.582028, 48.577861, 48.576194, 48.569917, 
    48.56575, 48.562, 48.566167, 48.5595, 48.5595, 48.556194, 48.556139, 
    48.55825, 48.562444, 48.562417, 48.567444, 48.567, 48.562833, 48.569111, 
    48.570306, 48.576167, 48.577, 48.59325, 48.594889, 48.612833, 48.622, 
    48.626167, 48.645361, 48.652861, 48.655361, 48.665722, 48.669472, 
    48.663667, 48.674083, 48.689917, 48.696583, 48.700722, 48.699528, 
    48.689111, 48.689528, 48.71575, 48.721194, 48.722444, 48.729917, 
    48.742417, 48.746583, 48.746167, 48.752417, 48.7645, 48.775361, 
    48.778667, 48.782, 48.778278, 48.776167, 48.7795, 48.773694, 48.773694, 
    48.76325, 48.757028, 48.739139, 48.715361, 48.7145, 48.719889, 48.731167, 
    48.731194, 48.738278, 48.754111, 48.767417, 48.772417, 48.784528, 
    48.786167, 48.801167, 48.800306, 48.803639, 48.801583, 48.789083, 
    48.788694, 48.819083, 48.849889, 48.860306, 48.881167, 48.885361, 
    48.894111, 48.897, 48.907028, 48.911167, 48.922444, 48.931583, 48.942028, 
    48.932806, 48.932028, 48.9395, 48.944944, 48.958694, 48.991972, 
    48.991556, 48.986139, 48.982861, 48.977444, 48.967806, 48.958667, 
    48.963667, 48.958694, 48.972417, 48.97325, 48.983694, 49, 49, 49, 49, 49, 
    49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 48.97825, 
    48.974556, 48.977, 48.971139, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 
    49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 
    49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 
    49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 
    49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 
    49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 
    49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 
    49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 
    49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 
    49, 49, 49, 49, 49, 49, 48.995778, 48.993778, 49, 49, 49, 49, 49, 49, 49, 
    49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 
    49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 
    49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 
    49, 49, 49, 49, 49, 49, 49, 49, 49, 48.996222, 45.871056, 43.552083, 
    44.509694, 41.162028, 38.104139, 37.694528, 34.928694, 28.016639, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28.001667, 28.000833, 28, 28, 28.001667, 28.005833, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28.031667, 30.374111, 29.1245, 28.004806, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28.011056, 28.003028, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 
    28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, 28, NaN, NaN, 
    48.999556, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 
    49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 
    49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 
    49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 
    49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 
    49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 
    49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 
    49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 
    49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 
    49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 
    49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 
    48.989917, 48.987417, 48.988639, 48.981167, 48.991167, 48.992028, 
    48.997861, 49, 49, 48.99825, 48.996972, 49, 49, 49, 49, 49, 49, 49, 49, 
    49, 49, 48.9995, 48.996167, 48.982028, 48.968667, 48.962861, 48.965333, 
    48.9595, 48.93825, 48.929528, 48.918667, 48.919083, 48.929083, 48.929556, 
    48.919111, 48.917417, 48.909944, 48.903639, 48.906167, 48.903278, 
    48.898306, 48.893694, 48.896167, 48.894083, 48.889528, 48.893278, 
    48.885361, 48.885333, 48.881139, 48.885333, 48.862833, 48.862861, 
    48.856194, 48.850361, 48.842417, 48.823278, 48.821167, 48.822, 48.814083, 
    48.792861, 48.803222, 48.808694, 48.799917, 48.789972, 48.779944, 
    48.779528, 48.768306, 48.744056, 48.745333, 48.752861, 48.752833, 
    48.767861, 48.757417, 48.755333, 48.7645, 48.764472, 48.76075, 48.758222, 
    48.759472, 48.75075, 48.747444, 48.733667, 48.718722, 48.7045, 48.694944, 
    48.660778, 48.654528, 48.655333, 48.659472, 48.657417, 48.649111, 
    48.633278, 48.615778, 48.598278, 48.582472, 48.569139, 48.561167, 
    48.557833, 48.549111, 48.536611, 48.52575, 48.516611, 48.509917, 
    48.507806, 48.515722, 48.547833, 48.553667, 48.577028, 48.575361, 
    48.568694, 48.571583, 48.579944, 48.589889, 48.597444, 48.599111, 
    48.602417, 48.61075, 48.627417, 48.629528, 48.627028, 48.635778, 
    48.642028, 48.654917, 48.662861, 48.664472, 48.668694, 48.667833, 
    48.6745, 48.677444, 48.681167, 48.68075, 48.687028, 48.689889, 48.694556, 
    48.699528, 48.691194, 48.688667, 48.682389, 48.680333, 48.682417, 
    48.674528, 48.674472, 48.680361, 48.677417, 48.6795, 48.675778, 48.67325, 
    48.670333, 48.667, 48.671194, 48.6695, 48.661139, 48.662444, 48.653278, 
    48.646611, 48.628278, 48.599944, 48.593667, 48.592, 48.598694, 48.597444, 
    48.564083, 48.559083, 48.516583, 48.496167, 48.4945, 48.498667, 
    48.497028, 48.489056, 48.477389, 48.464556, 48.452417, 48.450306, 
    48.458694, 48.45575, 48.449944, 48.437444, 48.437, 48.426583, 48.422389, 
    48.411194, 48.409528, 48.412861, 48.406167, 48.411167, 48.407833, 
    48.410333, 48.402806, 48.406167, 48.408667, 48.415333, 48.415778, 
    48.423667, 48.425361, 48.422861, 48.427833, 48.428722, 48.420722, 
    48.417028, 48.422028, 48.421167, 48.426167, 48.427833, 48.424528, 
    48.425306, 48.430778, 48.433722, 48.43325, 48.440333, 48.442444, 
    48.443278, 48.4495, 48.457, 48.448222, 48.442389, 48.439056, 48.432417, 
    48.429083, 48.39825, 48.392028, 48.392, 48.387444, 48.3845, 48.387, 
    48.382833, 48.3845, 48.3795, 48.354083, 48.342, 48.342389, 48.336194, 
    48.343278, 48.324972, 48.319528, 48.3095, 48.312833, 48.313694, 
    48.307833, 48.315333, 48.314556, 48.319917, 48.326194, 48.325361, 
    48.329111, 48.341167, 48.337833, 48.337, 48.333667, 48.335306, 48.32825, 
    48.324917, 48.323278, 48.316167, 48.312833, 48.316194, 48.3195, 
    48.334528, 48.338667, 48.336222, 48.338667, 48.337833, 48.35325, 
    48.357833, 48.361611, 48.362833, 48.36575, 48.375333, 48.377, 48.368667, 
    48.368639, 48.363667, 48.368694, 48.365333, 48.363667, 48.38325, 
    48.388222, 48.385306, 48.393667, 48.389111, 48.3895, 48.385389, 
    48.388639, 48.388667, 48.386583, 48.377, 48.383694, 48.378694, 48.372, 
    48.362417, 48.357028, 48.360333, 48.35825, 48.354472, 48.357889, 
    48.370361, 48.368667, 48.363639, 48.363694, 48.357056, 48.370306, 
    48.378694, 48.381139, 48.377028, 48.383694, 48.394528, 48.392833, 
    48.394889, 48.405361, 48.409556, 48.419556, 48.422083, 48.433694, 
    48.432083, 48.438694, 48.446222, 48.452056, 48.456222, 48.469528, 
    48.484556, 48.491639, 48.5045, 48.507833, 48.516194, 48.520333, 
    48.517833, 48.522833, 48.521972, 48.526194, 48.525333, 48.532444, 
    48.542028, 48.5545, 48.559889, 48.567417, 48.576167, 48.562861, 
    48.560306, 48.553667, 48.542833, 48.553667, 48.556972, 48.555333, 
    48.562833, 48.564528, 48.5695, 48.573639, 48.579472, 48.583667, 48.5895, 
    48.592833, 48.612028, 48.611139, 48.616972, 48.627861, 48.629472, 
    48.637028, 48.642, 48.660361, 48.661139, 48.657833, 48.666139, 48.681139, 
    48.669944, 48.668667, 48.675306, 48.675333, 48.681139, 48.699472, 
    48.700361, 48.7045, 48.705389, 48.712917, 48.722083, 48.720417, 48.72625, 
    48.730861, 48.739167, 48.747472, 48.757472, 48.757889, 48.761667, 
    48.764111, 48.774139, 48.788333, 48.792889, 48.797889, 48.7875, 48.7775, 
    48.77625, 48.771667, 48.770417, 48.775806, 48.777472, 48.78375, 
    48.787917, 48.783722, 48.786222, 48.78125, 48.785389, 48.781222, 
    48.784167, 48.789167, 48.789111, 48.791639, 48.798722, 48.79875, 
    48.802083, 48.802056, 48.806667, 48.81, 48.815389, 48.814583, 48.818722, 
    48.817861, 48.825361, 48.826278, 48.840389, 48.836639, 48.825806, 
    48.824556, 48.837472, 48.836639, 48.841611, 48.848361, 48.855417, 
    48.852083, 48.858306, 48.859139, 48.865, 48.868694, 48.878722, 48.881222, 
    48.885389, 48.887056, 48.884556, 48.877944, 48.885389, 48.883778, 
    48.886222, 48.892472, 48.896222, 48.899167, 48.902917, 48.907472, 
    48.915806, 48.915389, 48.919611, 48.917889, 48.922889, 48.921222, 
    48.925389, 48.91875, 48.919972, 48.928333, 48.929139, 48.934111, 
    48.935806, 48.940417, 48.939583, 48.944583, 48.947861, 48.945389, 
    48.938667, 48.952417, 48.953306, 48.959111, 48.961194, 48.966167, 
    48.973722, 48.976139, 48.978694, 48.975306, 48.979528, 48.989917, 
    48.996944, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 
    49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 
    49, 49, 49, 48.993639, 48.984528, 48.982861, 48.987, 48.983667, 
    48.987028, 48.983694, 48.981139, 48.984917, 48.989083, 48.992, 49, 49, 
    49, 49, 49, 49, 49, 49, 48.9975, 48.988722, 48.97825, 48.966222, 
    48.962083, 48.96375, 48.954528, 48.955833, 48.961639, 48.975806, 
    48.979556, 48.97375, 48.97375, 48.982889, 48.977917, 48.980389, 
    48.978306, 48.968722, 48.962889, 48.966222, 48.970833, 48.974167, 
    48.975417, 48.972889, 48.975389, 48.973722, 48.980389, 48.979972, 
    48.988333, 48.991639, 49, 49, 48.999528, 48.999167, 49, 49, 49, 49, 
    48.997472, 48.985389, 48.984583, 48.990417, 48.990417, 48.996222, 
    48.999556, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 
    49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 48.985, 48.979167, 
    48.974972, 48.970833, 48.96, 48.953333, 48.952889, 48.957083, 48.954139, 
    48.966222, 48.960806, 48.943722, 48.945806, 48.9525, 48.959167, 
    48.960417, 48.951222, 48.944556, 48.948278, 48.954556, 48.962028, 
    48.960806, 48.958333, 48.953722, 48.954972, 48.959528, 48.955417, 
    48.959139, 48.959611, 48.967056, 48.962889, 48.966222, 48.967917, 
    48.965389, 48.969583, 48.968694, 48.972028, 48.977083, 48.975833, 
    48.978306, 48.998306, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 
    49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 49, 48.999528, 
    48.985417, 48.98, 48.975389, 48.963694, 48.962889, 48.954556, 48.951194, 
    48.942889, 48.942056, 48.927472, 48.92125, 48.922083, 48.917917, 
    48.92625, 48.922528, 48.917056, 48.922889, 48.922111, 48.925389, 
    48.928278, 48.930833, 48.935417, 48.934583, 48.952917, 48.957056, 
    48.978778, 48.97875, 48.975806, 48.970806, 48.964944, 48.957889, 
    48.953333, 48.949556, 48.95125, 48.948722, 48.952083, 48.946222, 
    48.947028, 48.929972, 48.929972, 48.926667, 48.922083, 48.922083, 
    48.928306, 48.929167, 48.929972, 48.934583, 48.930361, 48.937056, 
    48.940389, 48.947056, 48.947056, 48.954583, 48.952917, 48.955028, 
    48.957028, 48.958306, 48.960861, 48.962472, 48.970833, 48.970417, 
    48.974944, 48.977861, 48.977444, 48.984972, 48.998694, 49, 49, 48.999194, 
    48.995389, 48.997028, 48.994556, 48.997889, 48.99625, 48.999556, NaN, 
    36.563611, 36.570556, 36.583889, 36.526667, 36.515278, 36.509167, 
    36.503889, 36.484167, 36.478889, 36.475833, 36.477778, 36.490833, 
    36.501667, 36.513611, 36.512778, 36.506944, 36.487222, 36.477222, 
    36.461389, 36.46, 36.4625, 36.459167, 36.451111, 36.435, 36.424444, 
    36.378889, 36.351667, 36.348611, 36.333611, 36.328611, 36.323611, 
    36.318056, 36.3075, 36.2975, 36.288333, 36.264722, 36.240833, 36.215278, 
    36.195, 36.171389, 36.166944, 36.164167, 36.169444, 36.169444, 36.155833, 
    36.160556, 36.146111, 36.142222, 36.146111, 36.153889, 36.155, 36.133889, 
    36.129444, 36.137222, 36.1275, 36.127222, 36.136944, 36.131667, 
    36.133056, 36.13, 36.125, 36.106667, 36.085556, 36.075556, 36.058056, 
    36.048333, 36.038056, 36.027222, 36.040278, 36.035833, 36.011667, 
    36.008889, 36.019444, 36.039722, 36.067778, 36.081389, 36.093333, 
    36.113611, 36.118889, 36.129444, 36.136111, 36.137778, 36.141667, 
    36.153056, 36.153056, 36.138333, 36.122778, 36.099167, 36.088889, 
    36.078889, 36.060556, 36.051667, 36.050556, 36.054167, 36.074444, 
    36.0775, 36.088889, 36.105, 36.111111, 36.112778, 36.101944, 36.113611, 
    36.135278, 36.136111, 36.113889, 36.11, 36.093056, 36.063889, 36.043056, 
    36.030556, 36.018333, 36.005833, 36.013889, 36.018333, 36.017778, 
    36.046111, 36.103889, 36.12, 36.123056, 36.181667, 36.191389, 36.188611, 
    36.195833, 36.1956272428, 36.178333, 36.167222, 36.123611, 36.117778, 
    36.116389, 36.116944, 36.126111, 36.124167, 36.116111, 36.100556, 
    36.086389, 36.067778, 36.056389, 36.049722, 36.048889, 36.042222, 
    36.030833, 36.057778, 36.065, 36.07, 36.095, 36.104722, 36.131944, 
    36.139444, 36.140833, 36.145278, 36.153056, 36.174167, 36.184444, 
    36.1975, 36.220833, 36.238056, 36.261018138893, 36.261944, 36.259444, 
    36.246667, 36.221667, 36.213333, 36.206111, 36.181111, 36.158889, 
    36.124167, 36.097222, 36.054444, 36.040833, 36.028889, 36.026667, 
    36.029444, 36.042222, 36.046667, 36.051667, 36.055278, 36.054444, 
    36.059444, 36.073611, 36.096667, 36.118333, 36.126111, 36.135556, 
    36.159444, 36.171389, 36.187222, 36.207778, 36.22, 36.280833, 36.334444, 
    36.350278, 36.381667, 36.402778, 36.417778, 36.433333, 36.450278, 
    36.461389, 36.47, 36.476944, 36.489444, 36.501944, 36.563611, NaN, 
    47.999556, 47.999556, 47.984139, 47.956639, 47.939139, 47.925028, 
    47.904583, 47.908333, 47.918333, 47.923722, 47.922083, 47.912083, 
    47.913694, 47.928278, 47.938306, 47.947472, 47.957472, 47.972056, 
    47.98875, 47.99125, 47.98875, 47.982083, 47.972056, 47.967083, 47.976639, 
    47.983306, 47.995, 48.007, 48.012, 48.028667, 48.03075, 48.037417, 
    48.051556, 48.059111, 48.073278, 48.110778, 48.151583, 48.1595, 
    48.162806, 48.161194, 48.156194, 48.1595, 48.155333, 48.155361, 
    48.180361, 48.193667, 48.200361, 48.211167, 48.213667, 48.217444, 
    48.23075, 48.259917, 48.279111, 48.304056, 48.333278, 48.364083, 
    48.374056, 48.402861, 48.405333, 48.40075, 48.397389, 48.397028, 48.412, 
    48.4095, 48.396972, 48.3945, 48.397444, 48.38825, 48.375778, 48.356194, 
    48.348694, 48.330333, 48.323694, 48.321194, 48.309111, 48.299111, 
    48.282861, 48.280361, 48.272028, 48.274083, 48.284083, 48.297028, 
    48.297889, 48.292, 48.289111, 48.279944, 48.267861, 48.267806, 48.273278, 
    48.281972, 48.28325, 48.287889, 48.287861, 48.276583, 48.264111, 
    48.251611, 48.242889, 48.238694, 48.237028, 48.231972, 48.233694, 
    48.226611, 48.224083, 48.215333, 48.215333, 48.222806, 48.222028, 
    48.225306, 48.223694, 48.227028, 48.223694, 48.220361, 48.222028, 
    48.20825, 48.194944, 48.194528, 48.184944, 48.159889, 48.146583, 
    48.133278, 48.117417, 48.10325, 48.079917, 48.075778, 48.054083, 
    48.051194, 48.044889, 48.017028, 48.017028, 48.021167, 48.037417, 
    48.06325, 48.076611, 48.09575, 48.098667, 48.096167, 48.097833, 
    48.052028, 48.045333, 48.042, 48.037, 48.034528, 47.999556, NaN, 
    48.456194, 48.456194, 48.457, 48.461167, 48.4595, 48.4695, 48.47325, 
    48.480806, 48.484111, 48.489528, 48.491139, 48.487806, 48.480333, 
    48.4845, 48.482028, 48.491167, 48.4895, 48.492028, 48.492, 48.498667, 
    48.50575, 48.513694, 48.515722, 48.519972, 48.529944, 48.549083, 
    48.550778, 48.567444, 48.572833, 48.568667, 48.569944, 48.577833, 
    48.570333, 48.573639, 48.57575, 48.589056, 48.591972, 48.5845, 48.583722, 
    48.580333, 48.586639, 48.59325, 48.594528, 48.604917, 48.608694, 
    48.599472, 48.600333, 48.5945, 48.591556, 48.59825, 48.599917, 48.607, 
    48.609528, 48.607028, 48.609944, 48.616611, 48.620722, 48.625361, 
    48.625361, 48.622861, 48.622444, 48.620333, 48.620306, 48.623694, 
    48.621194, 48.61325, 48.600333, 48.592861, 48.593667, 48.582833, 
    48.569528, 48.5645, 48.562056, 48.554056, 48.547417, 48.545306, 
    48.537889, 48.534528, 48.527028, 48.534917, 48.537028, 48.537028, 
    48.528667, 48.529083, 48.521194, 48.515361, 48.516167, 48.521139, 
    48.5195, 48.522, 48.517444, 48.509944, 48.505722, 48.503278, 48.494917, 
    48.484917, 48.475722, 48.472028, 48.461222, 48.463667, 48.461222, 
    48.468639, 48.465722, 48.450361, 48.456194, NaN, 48.477417, 48.478222, 
    48.517417, 48.522833, 48.523278, 48.520778, 48.515333, 48.509528, 
    48.501972, 48.507, 48.5045, 48.505333, 48.513278, 48.519917, 48.520778, 
    48.537444, 48.551556, 48.550361, 48.556167, 48.557833, 48.570722, 
    48.573639, 48.5545, 48.5545, 48.565333, 48.563278, 48.554944, 48.549917, 
    48.544083, 48.542028, 48.543667, 48.536583, 48.534083, 48.512444, 
    48.504111, 48.481556, 48.474083, 48.46575, 48.460778, 48.457861, 
    48.462833, 48.459917, 48.448278, 48.447, 48.4495, 48.460333, 48.461583, 
    48.464917, 48.469083, 48.466972, 48.47075, 48.478667, 48.471583, 
    48.457417, 48.453694, 48.452833, 48.44825, 48.442417, 48.431583, 
    48.431972, 48.426139, 48.422, 48.425333, 48.430361, 48.427, 48.431167, 
    48.424472, 48.430333, 48.427028, 48.42325, 48.423639, 48.419528, 
    48.421194, 48.417833, 48.420389, 48.422833, 48.42825, 48.432417, 
    48.435333, 48.438722, 48.4395, 48.434056, 48.433667, 48.442444, 
    48.446167, 48.445333, 48.450361, 48.446139, 48.448667, 48.446139, 
    48.447806, 48.441583, 48.440333, 48.451583, 48.455361, 48.455361, 
    48.460333, 48.466167, 48.458667, 48.456167, 48.457833, 48.477417, NaN, 
    48.939917, 48.941639, 48.942417, 48.946167, 48.937861, 48.9195, 
    48.915361, 48.893639, 48.892417, 48.897028, 48.894472, 48.887861, 
    48.853694, 48.843694, 48.859528, 48.860333, 48.867028, 48.866611, 
    48.866167, 48.860333, 48.844528, 48.840778, 48.840306, 48.850361, 
    48.844472, 48.849528, 48.858694, 48.855806, 48.854528, 48.857444, 
    48.846167, 48.841972, 48.845722, 48.846194, 48.841167, 48.833639, 
    48.828667, 48.812833, 48.812833, 48.803667, 48.798694, 48.797861, 
    48.790361, 48.787028, 48.778222, 48.774083, 48.766194, 48.768278, 
    48.759917, 48.752833, 48.753667, 48.757806, 48.754528, 48.757889, 
    48.7545, 48.766167, 48.770389, 48.756194, 48.749111, 48.732417, 48.7145, 
    48.714528, 48.733667, 48.745361, 48.761583, 48.767861, 48.772, 48.777444, 
    48.78575, 48.790333, 48.792028, 48.788667, 48.789889, 48.816167, 
    48.818667, 48.824944, 48.851194, 48.852, 48.857444, 48.865333, 48.862444, 
    48.876194, 48.886583, 48.888278, 48.896583, 48.901583, 48.913278, 
    48.920778, 48.925778, 48.939917, NaN, 48.614889, 48.61575, 48.631167, 
    48.61575, 48.609528, 48.616611, 48.631639, 48.63825, 48.657, 48.666167, 
    48.677833, 48.6845, 48.687417, 48.692, 48.693639, 48.704111, 48.712, 
    48.711167, 48.715333, 48.715333, 48.712, 48.713639, 48.705361, 48.704528, 
    48.697, 48.693694, 48.684528, 48.680361, 48.66075, 48.657, 48.649139, 
    48.642806, 48.639528, 48.641194, 48.638278, 48.6345, 48.632417, 
    48.624944, 48.619056, 48.601972, 48.606167, 48.5995, 48.602028, 
    48.600306, 48.621167, 48.617861, 48.620361, 48.618667, 48.646972, 
    48.642861, 48.65075, 48.689944, 48.694472, 48.688639, 48.693667, 
    48.68575, 48.683278, 48.671583, 48.65575, 48.649528, 48.646139, 
    48.637389, 48.622417, 48.612417, 48.601139, 48.591972, 48.595361, 
    48.588667, 48.592, 48.597028, 48.592861, 48.591139, 48.592861, 48.598694, 
    48.597, 48.617389, 48.625778, 48.631222, 48.6295, 48.642861, 48.632417, 
    48.632028, 48.624083, 48.619111, 48.600361, 48.601972, 48.610778, 
    48.614889, NaN, 48.04, 48.033889, 48.025, 48.015, 48.004444, 47.996944, 
    47.9925, 47.987222, 47.976389, 47.958889, 47.953889, 47.961111, 
    47.956944, 47.978056, 47.995, 48.013056, 48.023889, 48.04, 48.051944, 
    48.071944, 48.090556, 48.115556, 48.127222, 48.134444, 48.13, 48.135278, 
    48.149167, 48.151667, 48.145278, 48.150833, 48.161944, 48.176944, 48.18, 
    48.1775, 48.181111, 48.186944, 48.2075, 48.218333, 48.231944, 48.255833, 
    48.285278, 48.286944, 48.284167, 48.288611, 48.306111, 48.3125, 
    48.313056, 48.303333, 48.309722, 48.309444, 48.299167, 48.266944, 
    48.253611, 48.247222, 48.243611, 48.254167, 48.261944, 48.284167, 
    48.286667, 48.274167, 48.252778, 48.245278, 48.247222, 48.258056, 
    48.261111, 48.260556, 48.254444, 48.239722, 48.226667, 48.216667, 
    48.198889, 48.182778, 48.181667, 48.189444, 48.191111, 48.184167, 
    48.135556, 48.096111, 48.04, NaN, 33.989778, 33.99, 33.988111, 33.972306, 
    33.971444, 33.967111, 33.969056, 33.961472, 33.959833, 33.964, 33.963, 
    33.959639, 33.962278, 33.959694, 33.963139, 33.963861, 33.960389, 
    33.970667, 33.968028, 33.978917, 33.980611, 34.009556, 34.018333, 
    34.031889, 34.035778, 34.04925, 34.057611, 34.056, 34.059944, 34.061194, 
    34.070056, 34.075111, 34.078417, 34.078444, 34.074111, 34.075972, 
    34.071722, 34.072667, 34.060694, 34.053694, 34.054833, 34.051972, 
    34.054167, 34.057528, 34.058306, 34.056389, 34.060083, 34.054056, 
    34.054083, 34.047472, 34.0485, 34.044194, 34.035333, 34.030167, 
    34.021917, 34.021806, 34.018389, 34.021056, 34.01775, 34.015972, 
    34.018639, 34.030972, 34.036028, 34.041028, 34.05425, 34.052278, 
    34.057556, 34.05, 34.043417, 34.03675, 34.026861, 34.022444, 34.0065, 
    33.998083, 33.996472, 33.989778, NaN, 40.886389, 40.891111, 40.906389, 
    40.908333, 40.876389, 40.87, 40.865556, 40.829722, 40.808333, 40.781944, 
    40.771389, 40.768333, 40.771944, 40.79, 40.7975, 40.806944, 40.819444, 
    40.824167, 40.825833, 40.831111, 40.803056, 40.768611, 40.765, 40.779444, 
    40.781111, 40.762778, 40.749167, 40.741389, 40.7375, 40.733333, 
    40.730833, 40.718333, 40.716111, 40.721944, 40.735556, 40.741389, 
    40.758056, 40.755556, 40.743333, 40.748056, 40.756667, 40.757778, 
    40.744444, 40.74, 40.744444, 40.756111, 40.770833, 40.7775, 40.778333, 
    40.758056, 40.756389, 40.76, 40.760556, 40.764167, 40.769444, 40.783889, 
    40.788611, 40.793611, 40.794444, 40.7875, 40.773056, 40.769167, 
    40.769722, 40.7775, 40.794444, 40.803333, 40.825833, 40.843611, 
    40.863889, 40.886389, NaN, 47.728333, 47.725833, 47.714167, 47.705278, 
    47.717222, 47.715278, 47.704722, 47.707778, 47.711389, 47.723056, 
    47.746667, 47.763611, 47.789167, 47.792222, 47.788333, 47.778611, 
    47.7525, 47.747222, 47.745278, 47.750556, 47.758889, 47.7845465144821, 
    47.8185965432, 47.856944, 47.920833, 47.967778, 48.017222, 48.048056, 
    48.060556, 48.066944, 48.058056, 48.056389, 48.058333, 48.062222, 
    48.083611, 48.0875, 48.090278, 48.074444, 48.065278, 48.045833, 48.0225, 
    47.998056, 47.961111, 47.920833, 47.914722, 47.908611, 47.91, 47.907778, 
    47.878056, 47.870556, 47.865833, 47.849167, 47.841667, 47.838611, 
    47.8325, 47.825278, 47.813889, 47.823056, 47.824444, 47.818056, 
    47.807778, 47.806389, 47.8125, 47.8125, 47.801667, 47.795833, 47.784722, 
    47.771667, 47.751944, 47.728333, NaN, 28.99775, 29, 29.012417, 29.024667, 
    29.039944, 29.049806, 29.056694, 29.060917, 29.075111, 29.080056, 
    29.083472, 29.124306, 29.144611, 29.155722, 29.159611, 29.16275, 
    29.179528, 29.178639, 29.184306, 29.178722, 29.179361, 29.187583, 
    29.188417, 29.196194, 29.197028, 29.191972, 29.184333, 29.170028, 
    29.168417, 29.155694, 29.13575, 29.113722, 29.107833, 29.101778, 29.069, 
    29.014389, 29.002639, 28.985222, 28.980667, 28.968139, 28.942472, 
    28.929306, 28.917556, 28.897194, 28.896806, 28.892917, 28.886028, 
    28.886194, 28.890972, 28.886778, 28.883389, 28.884556, 28.889528, 
    28.894222, 28.899583, 28.909667, 28.918444, 28.922722, 28.935861, 
    28.9395, 28.941917, 28.950361, 28.957, 28.957694, 28.963, 28.973917, 
    28.985694, 28.99275, 28.99775, NaN, 42.613333, 42.620278, 42.628611, 
    42.631389, 42.628333, 42.603333, 42.590556, 42.587222, 42.585556, 
    42.578889, 42.555556, 42.550833, 42.544444, 42.540556, 42.521389, 
    42.505833, 42.501389, 42.501389, 42.498611, 42.485278, 42.481667, 
    42.476389, 42.4475, 42.421389, 42.410833, 42.407222, 42.417778, 
    42.419444, 42.413056, 42.389722, 42.390278, 42.399167, 42.404167, 
    42.397778, 42.366389, 42.355556, 42.352222, 42.342778, 42.318333, 
    42.308056, 42.303056, 42.316111, 42.317222, 42.299722, 42.28, 42.251667, 
    42.241667, 42.242222, 42.265278, 42.280556, 42.296389, 42.316667, 
    42.344722, 42.365833, 42.384722, 42.416389, 42.470556, 42.4725, 
    42.469722, 42.474167, 42.4925, 42.504722, 42.513333, 42.524444, 
    42.536389, 42.579167, 42.613333, NaN, 33.4775, 33.479111, 33.474583, 
    33.476222, 33.47375, 33.477917, 33.467889, 33.46625, 33.462083, 
    33.454583, 33.442056, 33.448778, 33.442917, 33.441222, 33.428722, 
    33.427917, 33.416222, 33.417889, 33.409583, 33.410417, 33.406694, 
    33.396694, 33.390028, 33.383306, 33.374583, 33.359139, 33.349139, 
    33.345806, 33.344583, 33.336694, 33.320833, 33.309139, 33.301222, 
    33.299583, 33.307917, 33.312889, 33.31875, 33.320444, 33.317083, 
    33.317056, 33.325361, 33.341667, 33.356639, 33.368278, 33.373361, 
    33.376694, 33.381194, 33.383333, 33.389944, 33.419194, 33.424528, 
    33.430833, 33.434528, 33.4275, 33.422056, 33.430389, 33.42875, 33.433722, 
    33.432889, 33.43625, 33.439139, 33.445806, 33.453722, 33.467056, 
    33.469556, 33.4775, NaN, 28.104083, 28.104194, 28.110833, 28.118306, 
    28.119167, 28.139306, 28.14, 28.148556, 28.173222, 28.220861, 28.232472, 
    28.244194, 28.247306, 28.270833, 28.279083, 28.298333, 28.305778, 
    28.329056, 28.349861, 28.353, 28.358139, 28.371083, 28.377528, 28.379139, 
    28.369111, 28.354778, 28.344917, 28.325611, 28.302472, 28.287278, 
    28.243167, 28.230667, 28.225861, 28.214833, 28.171472, 28.168194, 
    28.164889, 28.154028, 28.135833, 28.122333, 28.111667, 28.099639, 
    28.088639, 28.078222, 28.062861, 28.049583, 28.045417, 28.036389, 
    28.033389, 28.040806, 28.044222, 28.035, 28.043278, 28.041528, 28.043528, 
    28.053861, 28.061444, 28.083528, 28.096611, 28.105778, 28.107556, 
    28.10325, 28.104083, 28.095083, 28.104083, NaN, 33.982472, 33.982972, 
    33.985528, 33.983806, 33.970361, 33.942639, 33.942889, 33.936444, 
    33.930778, 33.917944, 33.914389, 33.912333, 33.90825, 33.907889, 
    33.901278, 33.896194, 33.893472, 33.902583, 33.9015, 33.911528, 
    33.912389, 33.916556, 33.915861, 33.922472, 33.923778, 33.945583, 
    33.950222, 33.969722, 33.979111, 33.986083, 33.990972, 33.996639, 
    33.996139, 34.000861, 34.004306, 34.009222, 34.011028, 34.005944, 
    34.004972, 34.008528, 34.006611, 34.009889, 34.01925, 34.025528, 
    34.027833, 34.024194, 34.020861, 34.020778, 34.025111, 34.039361, 34.037, 
    34.025944, 34.013222, 34, 33.993056, 33.9855, 33.981583, 33.982472, NaN, 
    47.6625, 47.664167, 47.675389, 47.674194, 47.664583, 47.67375, 47.673278, 
    47.68, 47.694167, 47.713361, 47.721194, 47.722083, 47.709556, 47.705, 
    47.699556, 47.70125, 47.697889, 47.692083, 47.69625, 47.697889, 
    47.708722, 47.707056, 47.709583, 47.694139, 47.6725, 47.661667, 
    47.651639, 47.634611, 47.624167, 47.620833, 47.619528, 47.625389, 
    47.620417, 47.622889, 47.620417, 47.627083, 47.624972, 47.616194, 
    47.618694, 47.61, 47.596694, 47.595806, 47.587889, 47.582056, 47.574583, 
    47.573722, 47.594972, 47.59625, 47.60375, 47.602944, 47.59125, 47.591222, 
    47.601639, 47.616667, 47.643306, 47.6625, NaN, 47.865556, 47.864167, 
    47.858056, 47.848056, 47.848056, 47.833611, 47.860833, 47.869444, 
    47.880278, 47.890833, 47.902778, 47.911667, 47.926944, 47.955, 47.973056, 
    47.995833, 48.008889, 48.029167, 48.037778, 48.048611, 48.053056, 
    48.074722, 48.098333, 48.134722, 48.191944, 48.204167, 48.22, 48.241667, 
    48.311389, 48.327222, 48.333056, 48.331111, 48.313889, 48.299167, 
    48.274167, 48.245, 48.218889, 48.211389, 48.204167, 48.170278, 48.150556, 
    48.114167, 48.09, 48.07, 48.059167, 48.045833, 48.0325, 48.010833, 
    48.000278, 47.989167, 47.965833, 47.948611, 47.902222, 47.884722, 
    47.865556, NaN, 46.895278, 46.893889, 46.884167, 46.859444, 46.86, 
    46.8775, 46.880556, 46.874444, 46.848333, 46.809444, 46.765, 46.734167, 
    46.670833, 46.641389, 46.630556, 46.623333, 46.629444, 46.643889, 
    46.645278, 46.639722, 46.630278, 46.610278, 46.586667, 46.575278, 
    46.540833, 46.523889, 46.518889, 46.521389, 46.547778, 46.551111, 
    46.559444, 46.565833, 46.599444, 46.610556, 46.62, 46.620833, 46.611389, 
    46.610833, 46.6175, 46.633056, 46.6425, 46.66, 46.726667, 46.761667, 
    46.798611, 46.82, 46.865556, 46.873333, 46.8725, 46.875, 46.882778, 
    46.890833, 46.892778, 46.895278, NaN, 48.999472, 49, 49, 49, 49, 
    48.984528, 48.958694, 48.950333, 48.947028, 48.937028, 48.925361, 
    48.920361, 48.920389, 48.911194, 48.906167, 48.896583, 48.892833, 48.892, 
    48.889528, 48.882, 48.885778, 48.887028, 48.881583, 48.876611, 48.87325, 
    48.861194, 48.861194, 48.865361, 48.866167, 48.859528, 48.858667, 
    48.866167, 48.870778, 48.876611, 48.885778, 48.887389, 48.892806, 
    48.897028, 48.897, 48.894083, 48.893694, 48.896583, 48.902028, 48.910361, 
    48.932833, 48.937861, 48.941194, 48.945306, 48.955333, 48.978667, 
    48.986583, 48.990778, 48.999472, NaN, 47.679167, 47.681389, 47.686944, 
    47.673056, 47.66, 47.6475, 47.635, 47.630278, 47.616944, 47.605, 
    47.598889, 47.596389, 47.598333, 47.596389, 47.585278, 47.55, 47.534444, 
    47.488889, 47.480278, 47.477778, 47.482778, 47.481389, 47.475278, 
    47.469722, 47.459167, 47.4575, 47.422778, 47.417222, 47.4225, 47.441389, 
    47.455, 47.476667, 47.476667, 47.471944, 47.4725, 47.478611, 47.491944, 
    47.503611, 47.513611, 47.530278, 47.553611, 47.558889, 47.591944, 
    47.612778, 47.632222, 47.636111, 47.638611, 47.6275, 47.628333, 
    47.633056, 47.651667, 47.679167, NaN, 47.344167, 47.3525, 47.366667, 
    47.375806, 47.380778, 47.391639, 47.399972, 47.414944, 47.423333, 47.455, 
    47.477889, 47.483333, 47.511639, 47.51125, 47.503278, 47.495778, 
    47.486639, 47.479556, 47.470389, 47.466639, 47.454167, 47.435806, 
    47.423306, 47.418333, 47.408306, 47.402028, 47.400389, 47.388333, 
    47.382083, 47.370417, 47.36875, 47.361667, 47.342917, 47.342889, 
    47.347472, 47.361639, 47.375417, 47.372056, 47.390806, 47.395806, 
    47.405417, 47.40125, 47.392056, 47.396278, 47.389167, 47.38375, 
    47.387056, 47.379972, 47.331222, 47.332861, 47.344167, NaN, 32.995472, 
    32.994972, 32.9855, 32.965556, 32.931, 32.911361, 32.89775, 32.879139, 
    32.837972, 32.818972, 32.815722, 32.820806, 32.824667, 32.820833, 
    32.812444, 32.811917, 32.799806, 32.804194, 32.816583, 32.814972, 
    32.820167, 32.819889, 32.842028, 32.844861, 32.850444, 32.851889, 
    32.863417, 32.868722, 32.878472, 32.885083, 32.888194, 32.907278, 
    32.906278, 32.917417, 32.919528, 32.925611, 32.948306, 32.968611, 
    33.009972, 33.014583, 33.014167, 33.032472, 33.03625, 33.029583, 
    33.033694, 33.026667, 33.007472, 33.007111, 33.002472, 32.995472, NaN, 
    47.698333, 47.708056, 47.729722, 47.761389, 47.764722, 47.765833, 
    47.763333, 47.76, 47.753611, 47.723889, 47.693056, 47.683333, 47.678333, 
    47.663611, 47.665833, 47.6625, 47.655278, 47.645556, 47.640556, 
    47.641111, 47.649444, 47.654722, 47.654167, 47.650833, 47.640278, 
    47.607778, 47.587778, 47.571389, 47.558889, 47.541111, 47.531389, 
    47.525556, 47.512222, 47.506389, 47.511667, 47.526944, 47.548889, 
    47.585556, 47.603611, 47.616111, 47.626944, 47.644444, 47.653889, 
    47.660278, 47.664444, 47.671389, 47.698333, NaN, 48.579083, 48.579639, 
    48.580333, 48.583694, 48.58325, 48.588667, 48.585361, 48.587806, 
    48.585361, 48.593694, 48.591167, 48.594944, 48.596139, 48.591167, 48.587, 
    48.580778, 48.573667, 48.576583, 48.579972, 48.584917, 48.587833, 
    48.5845, 48.579083, 48.565333, 48.566194, 48.562028, 48.565333, 
    48.563222, 48.558722, 48.561167, 48.553278, 48.547806, 48.547806, 
    48.552028, 48.548667, 48.555361, 48.552028, 48.558278, 48.562389, 
    48.563694, 48.558667, 48.559917, 48.564889, 48.568667, 48.565361, 
    48.569917, 48.579083, NaN, 39.647222, 39.656111, 39.665833, 39.672222, 
    39.689722, 39.691944, 39.687778, 39.666944, 39.661667, 39.658056, 
    39.654722, 39.646667, 39.62, 39.606667, 39.576389, 39.56, 39.541667, 
    39.538333, 39.538056, 39.525833, 39.521667, 39.522778, 39.533333, 
    39.534444, 39.520278, 39.519167, 39.521667, 39.529444, 39.533889, 
    39.540556, 39.5425, 39.545278, 39.551667, 39.560278, 39.571667, 
    39.575833, 39.580556, 39.576667, 39.566944, 39.564722, 39.57, 39.585556, 
    39.589167, 39.583056, 39.589444, 39.647222, NaN, 33.524167, 33.525278, 
    33.525, 33.517778, 33.511389, 33.5, 33.476389, 33.450833, 33.418889, 
    33.405278, 33.397778, 33.359444, 33.341944, 33.322222, 33.305278, 
    33.288056, 33.27, 33.237778, 33.211111, 33.176944, 33.174444, 33.163333, 
    33.116667, 33.107778, 33.110278, 33.123056, 33.126111, 33.121944, 33.125, 
    33.149167, 33.178056, 33.196389, 33.207778, 33.215278, 33.24, 33.280833, 
    33.3225, 33.333611, 33.342222, 33.348889, 33.348889, 33.357222, 
    33.496667, 33.513611, 33.524167, NaN, 39.22, 39.226111, 39.239722, 
    39.249444, 39.258611, 39.2525, 39.236111, 39.230278, 39.23, 39.236944, 
    39.233056, 39.206389, 39.180833, 39.166389, 39.151944, 39.133611, 
    39.103611, 39.090833, 39.081111, 39.075278, 39.074444, 39.068056, 39.025, 
    38.975278, 38.958333, 38.958056, 38.943056, 38.936944, 38.943333, 
    38.943056, 38.945833, 38.954722, 38.968611, 39.006111, 39.028333, 
    39.071389, 39.088889, 39.113056, 39.171944, 39.191111, 39.22, NaN, 
    39.1225, 39.125556, 39.127222, 39.123611, 39.119722, 39.106667, 
    39.066389, 39.053333, 39.043889, 39.0375, 39.035, 39.014444, 39.015556, 
    39.021389, 39.020556, 38.997778, 38.979444, 38.975278, 38.9675, 
    38.958333, 38.957222, 38.954167, 38.926667, 38.924722, 38.926667, 
    38.933333, 38.971667, 38.982222, 38.993056, 39.013056, 39.008333, 
    39.013611, 39.023611, 39.027222, 39.0275, 39.042222, 39.049444, 
    39.066667, 39.103056, 39.114722, 39.1225, NaN, 39.461389, 39.466389, 
    39.4725, 39.475278, 39.464167, 39.426111, 39.424722, 39.430278, 
    39.429722, 39.423611, 39.409167, 39.396944, 39.387222, 39.384167, 
    39.379167, 39.3725, 39.362778, 39.342222, 39.341944, 39.346389, 
    39.333333, 39.316389, 39.304167, 39.34, 39.351389, 39.355556, 39.374167, 
    39.380833, 39.398611, 39.408889, 39.416111, 39.418333, 39.408611, 
    39.409167, 39.412222, 39.428333, 39.435556, 39.439444, 39.443889, 
    39.461389, NaN, 34.013194, 34.014611, 34.016611, 34.024028, 34.031667, 
    34.031528, 34.027917, 34.024861, 34.0315, 34.028583, 34.030861, 
    34.032833, 34.038639, 34.039111, 34.048028, 34.054472, 34.0585, 
    34.060139, 34.054917, 34.051472, 34.05325, 34.064556, 34.071361, 
    34.073278, 34.077444, 34.074056, 34.065361, 34.057139, 34.054667, 
    34.048333, 34.047444, 34.049833, 34.041806, 34.025806, 34.022028, 
    34.019889, 34.017278, 34.019167, 34.013611, 34.013194, NaN, 47.083611, 
    47.088056, 47.098611, 47.101389, 47.096389, 47.085, 47.060833, 47.050833, 
    47.048889, 47.050833, 47.075, 47.099444, 47.100556, 47.0975, 47.0825, 
    47.072778, 47.066111, 47.059167, 47.051944, 47.047222, 47.023889, 47, 
    46.986111, 46.979722, 46.98, 46.981667, 46.996111, 46.997222, 46.992778, 
    46.994167, 46.997222, 47.003056, 47.008611, 47.010833, 47.010833, 
    47.005556, 47.011111, 47.026389, 47.061667, 47.083611, NaN, 48.746389, 
    48.746389, 48.730833, 48.726389, 48.725556, 48.722222, 48.72, 48.720556, 
    48.725, 48.743889, 48.743056, 48.7675, 48.773889, 48.788889, 48.795278, 
    48.814722, 48.870833, 48.877222, 48.903333, 48.929444, 48.948333, 
    48.975278, 48.986944, 49, 49, 49, 48.979444, 48.951111, 48.912778, 
    48.903611, 48.876944, 48.864444, 48.832778, 48.808611, 48.786111, 
    48.771111, 48.764722, 48.756111, 48.746389, NaN, 48.071611, 48.072417, 
    48.083694, 48.088694, 48.079944, 48.070778, 48.064111, 48.044889, 
    48.040778, 48.035778, 48.020361, 48.031583, 48.042417, 48.049111, 
    48.055306, 48.0545, 48.050333, 48.054944, 48.058222, 48.07075, 48.089111, 
    48.094111, 48.102861, 48.103667, 48.08825, 48.073278, 48.045722, 48.0395, 
    48.033278, 48.016556, 48.0095, 48.007806, 48.013667, 48.025389, 
    48.032306, 48.050806, 48.069111, 48.071611, NaN, 48.804083, 48.804944, 
    48.808694, 48.808278, 48.811583, 48.819111, 48.821972, 48.822, 48.817, 
    48.818639, 48.816194, 48.807417, 48.801194, 48.802861, 48.7945, 
    48.779944, 48.770778, 48.771194, 48.778694, 48.772861, 48.764889, 
    48.759917, 48.752, 48.747861, 48.743694, 48.739944, 48.736167, 48.742, 
    48.767861, 48.767833, 48.77075, 48.778278, 48.779917, 48.79075, 
    48.793278, 48.795389, 48.796611, 48.804083, NaN, 48.910556, 48.914722, 
    48.918333, 48.909444, 48.915833, 48.914444, 48.911944, 48.899444, 
    48.901111, 48.898889, 48.891111, 48.885833, 48.88, 48.871667, 48.865833, 
    48.855556, 48.855556, 48.849167, 48.837778, 48.809167, 48.804167, 
    48.798611, 48.798611, 48.803889, 48.809722, 48.824722, 48.824444, 
    48.831111, 48.843333, 48.850556, 48.860556, 48.8675, 48.873056, 
    48.884722, 48.889167, 48.895833, 48.910556, NaN, 39.723889, 39.724167, 
    39.722222, 39.724444, 39.713611, 39.709722, 39.710278, 39.700833, 
    39.703611, 39.696944, 39.703611, 39.701111, 39.675278, 39.672222, 
    39.679167, 39.679722, 39.675278, 39.665556, 39.649444, 39.641111, 
    39.655278, 39.655, 39.645, 39.627222, 39.624167, 39.63, 39.6525, 
    39.664722, 39.697222, 39.699722, 39.739167, 39.770556, 39.782222, 
    39.779444, 39.7525, 39.721667, 39.723889, NaN, 42.104444, 42.105278, 
    42.109167, 42.102222, 42.061389, 42.027222, 42.015556, 42.006944, 
    41.997222, 41.978611, 41.958333, 41.9525, 41.924444, 41.884444, 
    41.853889, 41.818333, 41.800833, 41.788056, 41.788333, 41.785, 41.772778, 
    41.77, 41.791389, 41.810833, 41.822222, 41.859722, 41.892778, 41.923889, 
    41.938056, 41.950833, 41.960278, 42.005833, 42.035556, 42.047222, 
    42.072778, 42.089722, 42.104444, NaN, 40.177778, 40.183333, 40.198056, 
    40.203889, 40.209444, 40.206111, 40.183056, 40.169722, 40.146111, 
    40.139722, 40.128333, 40.106111, 40.073611, 40.051389, 40.036389, 
    40.021111, 39.981111, 39.946944, 39.940833, 39.929722, 39.888333, 
    39.871389, 39.866944, 39.867222, 39.873611, 39.911389, 39.923333, 
    39.942778, 39.952778, 39.979444, 40.002778, 40.028056, 40.038056, 
    40.063889, 40.107778, 40.177778, NaN, 40.324722, 40.331944, 40.339722, 
    40.338889, 40.294444, 40.285, 40.280556, 40.269444, 40.258333, 40.230556, 
    40.191111, 40.180556, 40.150556, 40.141389, 40.140833, 40.143889, 
    40.1525, 40.164167, 40.169722, 40.176111, 40.173889, 40.1775, 40.183333, 
    40.195556, 40.226667, 40.2425, 40.244444, 40.21, 40.181389, 40.180278, 
    40.184167, 40.2, 40.223611, 40.269444, 40.324722, NaN, 31.670722, 
    31.672389, 31.676194, 31.690889, 31.676583, 31.695028, 31.709806, 
    31.730722, 31.750889, 31.764028, 31.784306, 31.8055, 31.803944, 31.78875, 
    31.763778, 31.748722, 31.7365, 31.746639, 31.713944, 31.682194, 
    31.671806, 31.666861, 31.661222, 31.658167, 31.658028, 31.661611, 
    31.663361, 31.668583, 31.682472, 31.689056, 31.684806, 31.695028, 
    31.687306, 31.6755, 31.670722, NaN, 48.668056, 48.671389, 48.678333, 
    48.663611, 48.645, 48.6275, 48.593889, 48.540278, 48.501944, 48.484722, 
    48.457778, 48.402222, 48.299722, 48.277778, 48.225833, 48.238333, 
    48.256944, 48.294722, 48.350278, 48.3875, 48.408889, 48.4275, 48.452222, 
    48.4575, 48.483889, 48.520833, 48.556111, 48.6075, 48.613333, 48.606944, 
    48.613333, 48.637222, 48.656389, 48.668056, NaN, 40.7225, 40.724444, 
    40.733611, 40.74, 40.733333, 40.720833, 40.701944, 40.693333, 40.688889, 
    40.695, 40.693333, 40.681111, 40.636389, 40.616111, 40.57, 40.558889, 
    40.551667, 40.549167, 40.554444, 40.6, 40.609444, 40.626944, 40.633889, 
    40.641944, 40.666389, 40.668333, 40.666667, 40.6525, 40.651389, 
    40.654722, 40.666111, 40.691389, 40.712778, 40.7225, NaN, 34.509722, 
    34.516111, 34.540556, 34.523889, 34.510556, 34.493889, 34.476667, 
    34.464167, 34.454722, 34.454722, 34.443333, 34.437222, 34.431111, 
    34.412222, 34.350278, 34.313056, 34.313889, 34.301944, 34.305833, 
    34.311667, 34.321389, 34.327778, 34.348611, 34.373333, 34.383056, 
    34.396389, 34.426389, 34.441667, 34.4525, 34.476389, 34.476389, 
    34.471111, 34.473611, 34.509722, NaN, 46.461528, 46.460222, 46.455389, 
    46.489167, 46.49875, 46.498694, 46.481611, 46.477917, 46.484583, 
    46.480806, 46.477444, 46.464583, 46.464944, 46.474972, 46.47625, 
    46.472472, 46.464611, 46.472889, 46.464139, 46.459972, 46.454167, 
    46.431667, 46.421639, 46.412056, 46.40875, 46.422472, 46.430806, 
    46.437472, 46.44625, 46.452917, 46.455889, 46.46075, 46.461528, NaN, 
    48.857444, 48.857833, 48.856194, 48.851194, 48.852028, 48.85825, 
    48.865778, 48.873639, 48.873722, 48.866139, 48.862861, 48.856611, 
    48.853694, 48.8595, 48.859917, 48.846611, 48.84575, 48.830722, 48.829111, 
    48.824528, 48.814083, 48.814528, 48.818694, 48.817806, 48.825361, 
    48.823694, 48.832861, 48.835333, 48.83575, 48.841583, 48.844083, 
    48.857444, NaN, 41.889444, 41.896944, 41.913333, 41.921667, 41.926389, 
    41.925556, 41.908611, 41.903889, 41.902222, 41.906944, 41.903611, 
    41.900833, 41.895278, 41.891389, 41.859444, 41.831389, 41.802778, 
    41.8025, 41.805278, 41.816667, 41.824722, 41.866389, 41.878611, 
    41.881944, 41.873611, 41.8625, 41.837222, 41.834444, 41.835556, 
    41.846944, 41.871389, 41.889444, NaN, 31.976667, 31.973132, 31.9675, 
    31.9475, 31.937778, 31.906111, 31.888611, 31.885556, 31.880278, 
    31.847778, 31.8425, 31.830556, 31.834444, 31.852222, 31.8675, 31.872778, 
    31.876944, 31.883333, 31.899444, 31.906389, 31.911944, 31.93, 31.931111, 
    31.934167, 31.977778, 31.980833, 31.971667, 31.972778, 31.9675, 
    31.965833, 31.966667, 31.976667, NaN, 38.665278, 38.668056, 38.685833, 
    38.689444, 38.688333, 38.683611, 38.645556, 38.63, 38.619722, 38.615278, 
    38.594722, 38.582778, 38.5575, 38.535278, 38.510556, 38.5, 38.523056, 
    38.5325, 38.537778, 38.535556, 38.504722, 38.5025, 38.516667, 38.506667, 
    38.506944, 38.514444, 38.518611, 38.551667, 38.569167, 38.608056, 
    38.647778, 38.665278, NaN, 43.380278, 43.383889, 43.383333, 43.378056, 
    43.376111, 43.381389, 43.378333, 43.342778, 43.333611, 43.322222, 
    43.319722, 43.308056, 43.302222, 43.301667, 43.305833, 43.300278, 
    43.286389, 43.288333, 43.296389, 43.279444, 43.280278, 43.291389, 
    43.313611, 43.326111, 43.336667, 43.341667, 43.349444, 43.361111, 
    43.379167, 43.381667, 43.380278, NaN, 33.265639, 33.265583, 33.257111, 
    33.229083, 33.225667, 33.217889, 33.218917, 33.215667, 33.21475, 
    33.218194, 33.218, 33.222389, 33.228167, 33.231472, 33.231417, 33.245944, 
    33.252556, 33.260389, 33.266417, 33.278306, 33.278222, 33.272639, 
    33.274167, 33.281472, 33.281667, 33.28575, 33.285861, 33.267611, 
    33.269222, 33.265639, NaN, 40.713611, 40.716389, 40.720278, 40.718333, 
    40.699167, 40.691944, 40.684722, 40.661111, 40.643611, 40.625833, 
    40.605556, 40.586111, 40.572778, 40.513611, 40.503333, 40.565556, 
    40.605556, 40.613611, 40.633333, 40.650278, 40.671667, 40.695556, 
    40.697222, 40.690556, 40.693056, 40.696944, 40.698611, 40.706389, 
    40.713611, NaN, 48.789944, 48.794056, 48.796972, 48.795333, 48.787806, 
    48.791583, 48.798667, 48.795333, 48.80575, 48.812028, 48.807, 48.813639, 
    48.796139, 48.7945, 48.789472, 48.784083, 48.781167, 48.7795, 48.778667, 
    48.773667, 48.769083, 48.763667, 48.765333, 48.762028, 48.762028, 
    48.762861, 48.773694, 48.780778, 48.789944, NaN, 35.574167, 35.580833, 
    35.595833, 35.614722, 35.623333, 35.588611, 35.563333, 35.551667, 
    35.526111, 35.513333, 35.500833, 35.471667, 35.433056, 35.415556, 
    35.381667, 35.346111, 35.3425, 35.3425, 35.354444, 35.388056, 35.415833, 
    35.440556, 35.489722, 35.503611, 35.520556, 35.534722, 35.54, 35.574167, 
    NaN, 48.904111, 48.904583, 48.907472, 48.914111, 48.915806, 48.920389, 
    48.919972, 48.925833, 48.9325, 48.934583, 48.937083, 48.94, 48.947889, 
    48.948722, 48.955417, 48.953722, 48.940833, 48.935833, 48.920806, 
    48.909556, 48.907861, 48.897028, 48.897056, 48.893722, 48.89375, 
    48.904111, NaN, 48.584083, 48.58575, 48.589083, 48.595778, 48.607861, 
    48.6095, 48.606167, 48.602, 48.597389, 48.590778, 48.589917, 48.569111, 
    48.563694, 48.565361, 48.55325, 48.551194, 48.554556, 48.553667, 
    48.544472, 48.540333, 48.555722, 48.562389, 48.570778, 48.584083, NaN, 
    40.269722, 40.274722, 40.281111, 40.278056, 40.272222, 40.263611, 
    40.251389, 40.233611, 40.231667, 40.294722, 40.294167, 40.300556, 
    40.301667, 40.292222, 40.265278, 40.259722, 40.244444, 40.225278, 
    40.206111, 40.191389, 40.195833, 40.2075, 40.238056, 40.269722, NaN, 
    37.084722, 37.0925, 37.098889, 37.070278, 37.055278, 37.049167, 
    37.039167, 37.016389, 37.009167, 36.994167, 36.977778, 36.976389, 
    36.981389, 36.99, 37.015278, 37.02, 37.026111, 37.020278, 37.021389, 
    37.025278, 37.045833, 37.058333, 37.076389, 37.084722, NaN, 48.729944, 
    48.734111, 48.747806, 48.745333, 48.735361, 48.735333, 48.714944, 48.707, 
    48.697, 48.698639, 48.694528, 48.692028, 48.682, 48.680333, 48.671972, 
    48.67075, 48.641194, 48.6495, 48.651167, 48.6795, 48.707417, 48.716194, 
    48.715361, 48.729944, NaN, 38.833333, 38.839722, 38.854167, 38.8375, 
    38.808333, 38.796667, 38.753333, 38.740278, 38.720833, 38.684167, 
    38.664167, 38.647222, 38.626111, 38.6025, 38.599722, 38.615833, 
    38.629722, 38.636667, 38.671389, 38.746944, 38.757222, 38.804444, 
    38.833333, NaN, 48.759889, 48.761611, 48.76075, 48.765333, 48.765778, 
    48.768694, 48.771194, 48.764083, 48.762833, 48.766972, 48.76325, 
    48.756167, 48.757833, 48.753694, 48.747, 48.747028, 48.753667, 48.752417, 
    48.747028, 48.750361, 48.752861, 48.75325, 48.759889, NaN, 48.653278, 
    48.654083, 48.637, 48.616139, 48.617028, 48.605306, 48.602417, 48.590361, 
    48.592833, 48.587833, 48.594917, 48.601556, 48.612861, 48.627417, 
    48.634083, 48.638667, 48.636639, 48.63325, 48.625333, 48.62575, 
    48.632417, 48.64075, 48.653278, NaN, 48.942472, 48.942889, 48.941222, 
    48.935389, 48.93875, 48.937083, 48.92875, 48.929556, 48.925417, 
    48.924583, 48.921667, 48.923722, 48.927917, 48.921222, 48.924583, 
    48.923722, 48.928694, 48.928361, 48.932083, 48.929528, 48.938333, 
    48.942472, NaN, 48.509944, 48.51075, 48.517028, 48.514111, 48.522833, 
    48.526194, 48.525333, 48.522028, 48.519944, 48.512444, 48.510389, 
    48.513694, 48.513278, 48.496167, 48.487, 48.480333, 48.482833, 48.481583, 
    48.492417, 48.49825, 48.509472, 48.509944, NaN, 42.691389, 42.694722, 
    42.710278, 42.716389, 42.723611, 42.732778, 42.731667, 42.727778, 
    42.716944, 42.690556, 42.640833, 42.616944, 42.601667, 42.580556, 
    42.538889, 42.533889, 42.531667, 42.540556, 42.584722, 42.633056, 
    42.666667, 42.691389, NaN, 48.684917, 48.688278, 48.690333, 48.690333, 
    48.688222, 48.685306, 48.684917, 48.680333, 48.6745, 48.682056, 
    48.681194, 48.674944, 48.67325, 48.665778, 48.664528, 48.670333, 
    48.677028, 48.667028, 48.660806, 48.658667, 48.667806, 48.684917, NaN, 
    48.589917, 48.594083, 48.607417, 48.612, 48.623667, 48.614944, 48.609944, 
    48.60825, 48.605333, 48.602389, 48.5995, 48.604472, 48.601583, 48.594917, 
    48.585722, 48.583667, 48.586583, 48.597028, 48.596556, 48.586167, 
    48.589917, NaN, 43.714444, 43.719444, 43.725278, 43.723333, 43.700278, 
    43.692778, 43.683889, 43.679167, 43.674444, 43.670556, 43.6675, 
    43.662222, 43.635, 43.631111, 43.639722, 43.663611, 43.671111, 43.685556, 
    43.6925, 43.708056, 43.714444, NaN, 38.800556, 38.803889, 38.819444, 
    38.821667, 38.813333, 38.794167, 38.780278, 38.725556, 38.714444, 
    38.695278, 38.694167, 38.7125, 38.7325, 38.751944, 38.757222, 38.760833, 
    38.737778, 38.738056, 38.742778, 38.787778, 38.800556, NaN, 43.294722, 
    43.295833, 43.2875, 43.266667, 43.255, 43.236667, 43.225, 43.203611, 
    43.201667, 43.203333, 43.19, 43.188056, 43.19, 43.201111, 43.250833, 
    43.270833, 43.2825, 43.288889, 43.295833, 43.294722, NaN, 46.198278, 
    46.199139, 46.202889, 46.204111, 46.206194, 46.205389, 46.207917, 
    46.207472, 46.214583, 46.214583, 46.217028, 46.217472, 46.210806, 
    46.201611, 46.185417, 46.185417, 46.188722, 46.18875, 46.198278, NaN, 
    48.843222, 48.843639, 48.840778, 48.848278, 48.850333, 48.832833, 48.832, 
    48.828222, 48.821194, 48.824083, 48.819917, 48.816139, 48.819917, 
    48.812028, 48.808667, 48.812833, 48.835778, 48.832444, 48.843222, NaN, 
    48.979111, 48.98075, 48.982833, 48.981222, 48.984528, 48.9795, 48.979972, 
    48.982861, 48.982444, 48.976611, 48.954889, 48.933694, 48.936167, 
    48.942833, 48.944472, 48.949083, 48.95825, 48.969056, 48.979111, NaN, 
    46.167222, 46.171111, 46.202778, 46.212778, 46.218889, 46.2025, 
    46.186667, 46.170833, 46.138056, 46.113889, 46.0825, 46.073889, 
    46.070278, 46.069167, 46.074167, 46.080278, 46.086667, 46.112778, 
    46.167222, NaN, 44.684722, 44.6925, 44.705, 44.701944, 44.652778, 
    44.620556, 44.614444, 44.615, 44.608056, 44.590278, 44.5725, 44.5425, 
    44.506389, 44.503333, 44.514167, 44.535833, 44.589167, 44.649167, 
    44.684722, NaN, 48.539944, 48.54325, 48.554944, 48.56075, 48.571583, 
    48.586611, 48.589556, 48.572861, 48.561167, 48.551167, 48.529889, 
    48.533667, 48.536972, 48.537833, 48.527, 48.526167, 48.529472, 48.539944, 
    NaN, 44.9725, 44.976667, 44.987778, 44.989167, 44.984444, 44.973611, 
    44.950833, 44.925, 44.9175, 44.915, 44.922222, 44.949444, 44.950278, 
    44.945833, 44.944722, 44.948611, 44.960278, 44.9725, NaN, 42.886667, 
    42.89, 42.901111, 42.903889, 42.902222, 42.875, 42.840833, 42.795556, 
    42.783611, 42.775, 42.770556, 42.771944, 42.787222, 42.810556, 42.849167, 
    42.871944, 42.886667, NaN, 48.571583, 48.573222, 48.583667, 48.584528, 
    48.587833, 48.588667, 48.582028, 48.560778, 48.546167, 48.537861, 
    48.539528, 48.532, 48.531139, 48.544944, 48.551611, 48.553278, 48.571583, 
    NaN, 37.663333, 37.669722, 37.678611, 37.673889, 37.630278, 37.625, 
    37.617778, 37.606111, 37.601111, 37.590278, 37.583889, 37.583056, 
    37.588611, 37.595833, 37.615556, 37.663333, NaN, 48.699944, 48.701583, 
    48.707028, 48.718694, 48.717833, 48.721139, 48.723667, 48.721611, 
    48.709944, 48.705722, 48.703278, 48.697444, 48.683667, 48.676194, 
    48.692861, 48.699944, NaN, 48.710722, 48.711583, 48.7095, 48.711194, 
    48.707, 48.707833, 48.714917, 48.719917, 48.721139, 48.714944, 48.704083, 
    48.697389, 48.692861, 48.692833, 48.697028, 48.710722, NaN, 48.924972, 
    48.925833, 48.929556, 48.929528, 48.925389, 48.925361, 48.916639, 
    48.915389, 48.91875, 48.915389, 48.914556, 48.917917, 48.922528, 
    48.92125, 48.924139, 48.924972, NaN, 47.294722, 47.2975, 47.307778, 
    47.3125, 47.299722, 47.300278, 47.2975, 47.264722, 47.257778, 47.217778, 
    47.190833, 47.225556, 47.236389, 47.258056, 47.273333, 47.294722, NaN, 
    48.998278, 49, 49, 49, 49, 49, 49, 49, 49, 48.989083, 48.98325, 
    48.969528, 48.969472, 48.980306, 48.981222, 48.998278, NaN, 42.987222, 
    42.985278, 42.978056, 42.9675, 42.948056, 42.9375, 42.930556, 42.926389, 
    42.923333, 42.927778, 42.934444, 42.951111, 42.974167, 42.984722, 
    42.987222, NaN, 48.76575, 48.767417, 48.767833, 48.762028, 48.757, 
    48.74325, 48.744472, 48.740778, 48.733667, 48.731194, 48.738722, 
    48.743639, 48.752833, 48.754528, 48.76575, NaN, 40.059722, 40.063889, 
    40.066111, 40.071667, 40.073056, 40.0625, 40.049444, 40.004722, 
    39.994444, 39.991389, 40.006667, 40.0325, 40.043333, 40.051111, 
    40.059722, NaN, 34.012167, 34.012528, 34.010917, 34.004167, 34.003389, 
    34.006806, 34.006833, 34.003278, 34.008306, 34.01475, 34.018444, 
    34.009111, 34.008694, 34.012167, NaN, 47.188333, 47.191667, 47.203056, 
    47.201944, 47.182222, 47.171944, 47.160278, 47.142778, 47.141944, 
    47.145278, 47.149167, 47.161667, 47.169722, 47.188333, NaN, 48.874139, 
    48.875, 48.882861, 48.883722, 48.890806, 48.89875, 48.897917, 48.892889, 
    48.893306, 48.880389, 48.882056, 48.874528, 48.874139, NaN, 46.175833, 
    46.1775, 46.182861, 46.179583, 46.181667, 46.184583, 46.182917, 
    46.184972, 46.189556, 46.187889, 46.181667, 46.172889, 46.175833, NaN, 
    48.989167, 48.99, 48.992917, 48.990389, 48.992056, 48.994583, 48.986667, 
    48.983694, 48.984556, 48.982111, 48.98125, 48.986222, 48.989167, NaN, 
    37.036667, 37.038611, 37.055556, 37.046111, 37.040278, 37.008056, 
    36.998611, 36.992222, 36.993333, 37.003889, 37.021111, 37.020833, 
    37.036667, NaN, 46.196667, 46.200833, 46.201194, 46.189111, 46.183306, 
    46.179611, 46.179583, 46.182889, 46.180417, 46.1825, 46.189194, 46.19625, 
    46.196667, NaN, 40.04, 40.0475, 40.052778, 40.055833, 40.042778, 
    40.026944, 40.001111, 39.993333, 39.996944, 40.000833, 40.006944, 40.04, 
    NaN, 48.71825, 48.721583, 48.727417, 48.731194, 48.731194, 48.72325, 
    48.714944, 48.704083, 48.702417, 48.6995, 48.707, 48.71825, NaN, 
    28.301472, 28.301639, 28.319111, 28.318778, 28.309083, 28.313028, 
    28.311583, 28.304917, 28.302417, 28.300583, 28.296333, 28.301472, NaN, 
    37.860806, 37.861667, 37.863306, 37.86875, 37.867917, 37.872083, 
    37.872056, 37.8675, 37.854167, 37.855417, 37.852861, 37.860806, NaN, 
    32.645278, 32.653056, 32.661111, 32.662778, 32.6425, 32.611389, 
    32.607778, 32.6125, 32.630278, 32.628611, 32.630556, 32.645278, NaN, 
    28.026528, 28.025889, 28.014833, 28.005611, 28.002833, 28.000917, 
    28.004583, 28.016944, 28.005, 28.004778, 28.011278, 28.026528, NaN, 
    48.617472, 48.618667, 48.617889, 48.607, 48.60325, 48.593667, 48.588639, 
    48.595778, 48.598694, 48.595778, 48.605361, 48.617472, NaN, 39.488333, 
    39.486944, 39.4725, 39.458611, 39.453889, 39.459167, 39.461111, 
    39.478611, 39.488889, 39.491111, 39.492778, 39.488333, NaN, 47.212778, 
    47.218889, 47.223611, 47.228333, 47.245556, 47.252778, 47.248889, 47.225, 
    47.220833, 47.206389, 47.206667, 47.212778, NaN, 31.728361, 31.728389, 
    31.730028, 31.742333, 31.745056, 31.753472, 31.756694, 31.754028, 
    31.749028, 31.745167, 31.731222, 31.728361, NaN, 45.540611, 45.537972, 
    45.532417, 45.518417, 45.524, 45.531806, 45.549833, 45.557056, 45.555222, 
    45.550667, 45.540611, NaN, 32.943611, 32.940833, 32.927778, 32.921667, 
    32.918611, 32.920556, 32.935278, 32.946944, 32.95, 32.949722, 32.943611, 
    NaN, 28.203611, 28.203972, 28.208222, 28.234694, 28.248222, 28.242694, 
    28.2225, 28.211806, 28.202056, 28.200722, 28.203611, NaN, 46.167222, 
    46.168611, 46.172778, 46.185278, 46.198611, 46.214167, 46.215, 46.208056, 
    46.195556, 46.169444, 46.167222, NaN, 48.908306, 48.910028, 48.910806, 
    48.915417, 48.912889, 48.914583, 48.907472, 48.904583, 48.907944, 
    48.906222, 48.908306, NaN, 48.831611, 48.833278, 48.831972, 48.814917, 
    48.812833, 48.816583, 48.81825, 48.821139, 48.821194, 48.818667, 
    48.831611, NaN, 29.824028, 29.824167, 29.817361, 29.806833, 29.811917, 
    29.808972, 29.818167, 29.819139, 29.822583, 29.820861, 29.824028, NaN, 
    29.969139, 29.9685, 29.963, 29.952472, 29.952444, 29.958389, 29.966472, 
    29.972722, 29.985556, 29.978333, 29.969139, NaN, 47.587222, 47.580833, 
    47.568611, 47.552778, 47.545278, 47.544722, 47.574444, 47.605833, 
    47.606389, 47.596944, 47.587222, NaN, 47.273611, 47.276944, 47.291944, 
    47.293611, 47.288056, 47.248889, 47.238889, 47.239444, 47.248333, 
    47.254444, 47.273611, NaN, 48.915778, 48.916639, 48.918333, 48.924611, 
    48.925389, 48.9225, 48.917889, 48.912889, 48.912111, 48.915778, NaN, 
    30.483306, 30.489167, 30.495417, 30.495417, 30.484167, 30.482472, 
    30.480417, 30.47625, 30.479583, 30.483306, NaN, 48.724944, 48.726611, 
    48.732, 48.737833, 48.734528, 48.7345, 48.726583, 48.71825, 48.7145, 
    48.724944, NaN, 30.091583, 30.093444, 30.093333, 30.083667, 30.081583, 
    30.082556, 30.089722, 30.087667, 30.089139, 30.091583, NaN, 48.822444, 
    48.824972, 48.835361, 48.832917, 48.837083, 48.834139, 48.827917, 
    48.822083, 48.820389, 48.822444, NaN, 41.846667, 41.856389, 41.860556, 
    41.846389, 41.840833, 41.812222, 41.810278, 41.812222, 41.822222, 
    41.846667, NaN, 37.086944, 37.089722, 37.096389, 37.0925, 37.086944, 
    37.063056, 37.051667, 37.051389, 37.06, 37.086944, NaN, 37.827444, 
    37.829167, 37.832944, 37.829972, 37.820833, 37.814194, 37.813333, 
    37.807056, 37.809167, 37.827444, NaN, 46.270917, 46.267722, 46.264694, 
    46.262417, 46.27075, 46.275639, 46.280972, 46.282472, 46.290861, 
    46.270917, NaN, 48.797417, 48.798278, 48.794472, 48.798694, 48.798694, 
    48.795333, 48.793278, 48.7895, 48.7895, 48.797417, NaN, 46.198333, 46.2, 
    46.20625, 46.205417, 46.209583, 46.209583, 46.205806, 46.198306, 
    46.187083, 46.198333, NaN, 46.245833, 46.246694, 46.24625, 46.248333, 
    46.252889, 46.24, 46.237917, 46.242861, 46.24125, 46.245833, NaN, 
    48.870806, 48.874167, 48.873722, 48.877472, 48.880806, 48.880417, 
    48.866639, 48.863722, 48.870806, NaN, 28.100083, 28.1005, 28.102528, 
    28.101806, 28.098556, 28.098472, 28.094167, 28.091694, 28.100083, NaN, 
    47.221667, 47.224444, 47.232778, 47.231667, 47.209444, 47.196111, 
    47.193889, 47.211944, 47.221667, NaN, 48.913306, 48.914167, 48.917917, 
    48.915806, 48.90875, 48.911222, 48.908722, 48.9125, 48.913306, NaN, 
    48.669111, 48.67075, 48.672833, 48.670333, 48.665361, 48.6645, 48.659889, 
    48.660333, 48.669111, NaN, 33.471417, 33.470722, 33.465361, 33.466083, 
    33.484472, 33.483361, 33.48925, 33.488333, 33.471417, NaN, 48.01825, 
    48.019056, 48.022861, 48.022861, 48.015306, 48.005778, 48.0045, 
    48.008667, 48.01825, NaN, 46.245806, 46.246667, 46.252083, 46.252056, 
    46.249583, 46.244972, 46.246222, 46.242861, 46.245806, NaN, 46.215, 
    46.215861, 46.227889, 46.227889, 46.223333, 46.218694, 46.209528, 
    46.214583, 46.215, NaN, 46.264972, 46.265833, 46.262889, 46.245806, 
    46.239556, 46.242083, 46.26, 46.260417, 46.264972, NaN, 47.541639, 
    47.542444, 47.547028, 47.543694, 47.540778, 47.5375, 47.530417, 47.53125, 
    47.541639, NaN, 48.620778, 48.622444, 48.630306, 48.620778, 48.609917, 
    48.607833, 48.610333, 48.617, 48.620778, NaN, 48.999167, 48.996639, 
    48.994139, 48.992083, 48.99375, 48.998333, 49, 49, 48.999167, NaN, 
    48.997833, 49, 49, 49, 49, 48.99325, 48.991167, 48.997028, 48.997833, 
    NaN, 48.846667, 48.849111, 48.851222, 48.84875, 48.848722, 48.830389, 
    48.841639, 48.847028, 48.846667, NaN, 48.619111, 48.619972, 48.622889, 
    48.618639, 48.621167, 48.612444, 48.612028, 48.619111, NaN, 46.235833, 
    46.236639, 46.241278, 46.24, 46.231194, 46.232472, 46.23625, 46.235833, 
    NaN, 48.64825, 48.650361, 48.642028, 48.637861, 48.637, 48.634083, 
    48.636194, 48.64825, NaN, 48.650722, 48.651139, 48.656583, 48.661167, 
    48.647417, 48.643667, 48.648694, 48.650722, NaN, 46.940111, 46.940139, 
    46.935361, 46.939639, 46.943278, 46.941889, 46.939139, 46.940111, NaN, 
    48.949167, 48.949972, 48.952861, 48.952917, 48.950361, 48.951667, 
    48.947083, 48.949167, NaN, 46.231639, 46.234139, 46.242917, 46.237917, 
    46.227528, 46.209556, 46.22125, 46.231639, NaN, 48.905778, 48.906639, 
    48.907083, 48.902917, 48.892028, 48.891222, 48.897056, 48.905778, NaN, 
    48.682444, 48.68325, 48.687417, 48.692, 48.685778, 48.678667, 48.677833, 
    48.682444, NaN, 48.954944, 48.956611, 48.947, 48.936167, 48.932, 48.942, 
    48.946167, 48.954944, NaN, 48.589944, 48.591556, 48.59325, 48.602, 
    48.598278, 48.591194, 48.587833, 48.589944, NaN, 48.424889, 48.42575, 
    48.430333, 48.429528, 48.42325, 48.423667, 48.4195, 48.424889, NaN, 
    38.103056, 38.104722, 38.098056, 38.086111, 38.083889, 38.085833, 
    38.090556, 38.103056, NaN, 28.312472, 28.312639, 28.318083, 28.318361, 
    28.312444, 28.31, 28.309833, 28.312472, NaN, 48.89575, 48.896611, 48.897, 
    48.893667, 48.87825, 48.873667, 48.882, 48.89575, NaN, 48.122417, 
    48.124472, 48.132028, 48.132, 48.127417, 48.126167, 48.121167, 48.122417, 
    NaN, 37.696389, 37.694444, 37.691528, 37.695639, 37.697194, 37.704, 
    37.703333, 37.696389, NaN, 48.683278, 48.684917, 48.684111, 48.682417, 
    48.677806, 48.680361, 48.683667, 48.683278, NaN, 48.601194, 48.601972, 
    48.601972, 48.595333, 48.592833, 48.5945, 48.599056, 48.601194, NaN, 
    48.863306, 48.86375, 48.865389, 48.863333, 48.861194, 48.857028, 
    48.863306, NaN, 38.058056, 38.065556, 38.057222, 38.0525, 38.045, 
    38.049167, 38.058056, NaN, 29.78825, 29.790083, 29.796639, 29.796611, 
    29.786389, 29.785083, 29.78825, NaN, 38.069167, 38.068056, 38.056944, 
    38.052778, 38.0625, 38.066667, 38.069167, NaN, 48.850833, 48.851639, 
    48.855361, 48.85625, 48.849139, 48.846222, 48.850833, NaN, 48.701583, 
    48.702444, 48.707806, 48.697417, 48.696611, 48.691194, 48.701583, NaN, 
    48.702417, 48.703222, 48.708667, 48.710361, 48.702444, 48.699472, 
    48.702417, NaN, 46.714222, 46.714972, 46.713444, 46.709778, 46.710083, 
    46.711917, 46.714222, NaN, 46.667333, 46.66675, 46.665472, 46.668083, 
    46.669583, 46.666611, 46.667333, NaN, 48.599056, 48.599917, 48.601194, 
    48.5945, 48.597, 48.5945, 48.599056, NaN, 48.464917, 48.468278, 
    48.471167, 48.464111, 48.457833, 48.457806, 48.464917, NaN, 31.812444, 
    31.811111, 31.804833, 31.808222, 31.808917, 31.812917, 31.812444, NaN, 
    48.663278, 48.664083, 48.666194, 48.666167, 48.663278, 48.661167, 
    48.663278, NaN, 48.524111, 48.524972, 48.528667, 48.528694, 48.522417, 
    48.5195, 48.524111, NaN, 48.514083, 48.517444, 48.517028, 48.509083, 
    48.507833, 48.512417, 48.514083, NaN, 28.30225, 28.303222, 28.312972, 
    28.316472, 28.304972, 28.295028, 28.30225, NaN, 46.701528, 46.701667, 
    46.704028, 46.710056, 46.704139, 46.701222, 46.701528, NaN, 48.476611, 
    48.477417, 48.4845, 48.488278, 48.4745, 48.473694, 48.476611, NaN, 
    28.855806, 28.855306, 28.853944, 28.849222, 28.851611, 28.855111, 
    28.855806, NaN, 48.487444, 48.488222, 48.494528, 48.4945, 48.491583, 
    48.4845, 48.487444, NaN, 48.873333, 48.874111, 48.877889, 48.876667, 
    48.872083, 48.873333, NaN, 46.199139, 46.199944, 46.202083, 46.200361, 
    46.194139, 46.199139, NaN, 46.665806, 46.666667, 46.673333, 46.675417, 
    46.664972, 46.665806, NaN, 48.363278, 48.364083, 48.367028, 48.363278, 
    48.359528, 48.363278, NaN, 48.396583, 48.398278, 48.402028, 48.402444, 
    48.397833, 48.396583, NaN, 48.883306, 48.884972, 48.88625, 48.880778, 
    48.879583, 48.883306, NaN, 46.2425, 46.243306, 46.251222, 46.249194, 
    46.242889, 46.2425, NaN, 48.613278, 48.614917, 48.614472, 48.607444, 
    48.606167, 48.613278, NaN, 46.2625, 46.265, 46.26375, 46.267083, 
    46.262472, 46.2625, NaN, 48.566611, 48.570778, 48.570361, 48.562417, 
    48.560333, 48.566611, NaN, 48.784944, 48.786194, 48.788694, 48.784917, 
    48.780361, 48.784944, NaN, 30.021333, 30.02075, 30.013972, 30.012194, 
    30.018306, 30.021333, NaN, 33.951694, 33.953083, 33.949611, 33.946639, 
    33.948972, 33.951694, NaN, 31.806639, 31.806528, 31.804111, 31.789056, 
    31.804417, 31.806639, NaN, 48.903306, 48.904167, 48.907917, 48.909556, 
    48.902917, 48.903306, NaN, 32.420556, 32.420806, 32.414917, 32.388111, 
    32.393417, 32.420556, NaN, 48.910806, 48.911667, 48.907056, 48.903722, 
    48.904583, 48.910806, NaN, 46.211667, 46.213333, 46.21625, 46.215, 
    46.210417, 46.211667, NaN, 28.876333, 28.875083, 28.86925, 28.87375, 
    28.881056, 28.876333, NaN, 48.929111, 48.93075, 48.932028, 48.925722, 
    48.921167, 48.929111, NaN, 48.436611, 48.438278, 48.442, 48.435778, 
    48.432056, 48.436611, NaN, 48.367444, 48.369944, 48.370333, 48.365778, 
    48.362, 48.367444, NaN, 34.019306, 34.019389, 34.017722, 34.014167, 
    34.013667, 34.019306, NaN, 46.242472, 46.242889, 46.243722, 46.239194, 
    46.238722, 46.242472, NaN, 46.963361, 46.966667, 46.966222, 46.96, 
    46.957917, 46.963361, NaN, 48.309889, 48.31075, 48.314528, 48.317833, 
    48.312, 48.309889, NaN, 48.891583, 48.894917, 48.894583, 48.88825, 
    48.886194, 48.891583, NaN, 48.435778, 48.436583, 48.444556, 48.431167, 
    48.430306, 48.435778, NaN, 48.858333, 48.859167, 48.862917, 48.855, 
    48.855417, 48.858333, NaN, 48.877444, 48.878722, 48.877056, 48.872889, 
    48.872083, 48.877444, NaN, 48.948278, 48.95, 48.952889, 48.950833, 
    48.94625, 48.948278, NaN, 48.972417, 48.974111, 48.9595, 48.955333, 
    48.959528, 48.972417, NaN, 28.114028, 28.114194, 28.115861, 28.112222, 
    28.110111, 28.114028, NaN, 48.747417, 48.748694, 48.749528, 48.74575, 
    48.742833, 48.747417, NaN, 48.36075, 48.361611, 48.366972, 48.36825, 
    48.359528, 48.36075, NaN, 28.036861, 28.037444, 28.039389, 28.042556, 
    28.039972, 28.036861, NaN, 28.035333, 28.033778, 28.030889, 28.036028, 
    28.037639, 28.035333, NaN, 34.058306, 34.057083, 34.054167, 34.056556, 
    34.061028, 34.058306, NaN, 48.971583, 48.974889, 48.97325, 48.970361, 
    48.972861, 48.971583, NaN, 48.888306, 48.889972, 48.892889, 48.889139, 
    48.887111, 48.888306, NaN, 46.669972, 46.668944, 46.664139, 46.666361, 
    46.671694, 46.669972, NaN, 37.9, 37.90125, 37.901222, 37.895, 37.895389, 
    37.9, NaN, 48.677444, 48.67825, 48.681167, 48.677417, 48.674556, 
    48.677444, NaN, 48.984083, 48.985778, 48.9845, 48.979889, 48.979528, 
    48.984083, NaN, 48.646556, 48.647417, 48.650333, 48.649944, 48.646167, 
    48.646556, NaN, 28.143333, 28.144194, 28.146778, 28.143, 28.140861, 
    28.143333, NaN, 47.906389, 47.907139, 47.907861, 47.902472, 47.903389, 
    47.906389, NaN, 48.50325, 48.504111, 48.507833, 48.507028, 48.502861, 
    48.50325, NaN, 48.306611, 48.30825, 48.312028, 48.306583, 48.304472, 
    48.306611, NaN, 48.540333, 48.539417, 48.536222, 48.539083, 48.542, 
    48.540333, NaN, 30.052639, 30.053056, 30.056333, 30.058806, 30.052806, 
    30.052639, NaN, 48.950028, 48.951639, 48.955389, 48.953333, 48.948722, 
    48.950028, NaN, 48.747417, 48.748278, 48.751222, 48.749917, 48.746194, 
    48.747417, NaN, 46.202444, 46.204972, 46.204556, 46.198722, 46.19875, 
    46.202444, NaN, 48.972444, 48.973306, 48.976222, 48.975, 48.969556, 
    48.972444, NaN, 32.418778, 32.42025, 32.419194, 32.414889, 32.414806, 
    32.418778, NaN, 48.535778, 48.536583, 48.538694, 48.537417, 48.5345, 
    48.535778, NaN, 48.392472, 48.393278, 48.395361, 48.391667, 48.389556, 
    48.392472, NaN, 46.873389, 46.877472, 46.880056, 46.88, 46.874, 
    46.873389, NaN, 48.829111, 48.829972, 48.830806, 48.82625, 48.829111, 
    NaN, 48.953306, 48.954528, 48.9525, 48.949556, 48.953306, NaN, 48.537444, 
    48.539944, 48.542861, 48.533667, 48.537444, NaN, 28, 28, 28.002111, 28, 
    28, NaN, 48.900778, 48.907472, 48.894917, 48.895333, 48.900778, NaN, 
    48.866667, 48.867444, 48.869944, 48.86625, 48.866667, NaN, 46.2075, 
    46.209167, 46.209972, 46.206222, 46.2075, NaN, 46.253333, 46.254139, 
    46.254139, 46.250389, 46.253333, NaN, 48.863333, 48.864111, 48.860778, 
    48.859556, 48.863333, NaN, 46.662472, 46.663306, 46.664556, 46.660806, 
    46.662472, NaN, 48.384139, 48.385, 48.382889, 48.377889, 48.384139, NaN, 
    48.157472, 48.158333, 48.160417, 48.155028, 48.157472, NaN, 48.684917, 
    48.687389, 48.686611, 48.681194, 48.684917, NaN, 48.799944, 48.80075, 
    48.798222, 48.797028, 48.799944, NaN, 34.040056, 34.040056, 34.045083, 
    34.040889, 34.040056, NaN, 48.084944, 48.08575, 48.093667, 48.085722, 
    48.084944, NaN, 48.696583, 48.697389, 48.704528, 48.696583, 48.696583, 
    NaN, 28.114139, 28.115361, 28.126583, 28.118694, 28.114139, NaN, 
    48.965778, 48.966639, 48.969528, 48.961611, 48.965778, NaN, 38.802556, 
    38.802333, 38.80075, 38.798778, 38.802556, NaN, 48.757028, 48.758222, 
    48.753694, 48.750333, 48.757028, NaN, 48.956639, 48.9575, 48.959972, 
    48.954611, 48.956639, NaN, 48.60325, 48.604083, 48.607861, 48.60325, 
    48.60325, NaN, 48.432417, 48.43325, 48.436194, 48.434083, 48.432417, NaN, 
    34.057667, 34.057444, 34.053333, 34.057444, 34.057667, NaN, 28.039167, 
    28.039972, 28.046083, 28.0485, 28.039167, NaN, 48.616583, 48.617444, 
    48.617861, 48.61575, 48.616583, NaN, 48.989917, 48.991583, 48.992889, 
    48.98825, 48.989917, NaN, 47.799778, 47.799667, 47.794889, 47.796194, 
    47.799778, NaN, 48.591583, 48.592444, 48.591583, 48.589528, 48.591583, 
    NaN, 48.396611, 48.399917, 48.402833, 48.394944, 48.396611, NaN, 
    48.554944, 48.559111, 48.561167, 48.557389, 48.554944, NaN, 48.412417, 
    48.414056, 48.414889, 48.411139, 48.412417, NaN, 48.697417, 48.699944, 
    48.702028, 48.695722, 48.697417, NaN, 48.844111, 48.846167, 48.843667, 
    48.841167, 48.844111, NaN, 48.82575, 48.826556, 48.82325, 48.822, 
    48.82575, NaN, 46.976972, 46.979806, 46.974139, 46.974028, 46.976972, 
    NaN, 48.919944, 48.920806, 48.9225, 48.918722, 48.919944, NaN, 29.375139, 
    29.374972, 29.37925, 29.377056, 29.375139, NaN, 48.939972, 48.941694, 
    48.937889, 48.933722, 48.939972, NaN, 48.965722, 48.967028, 48.964056, 
    48.958667, 48.965722, NaN, 37.697194, 37.695833, 37.697889, 37.700639, 
    37.697194, NaN, 48.442389, 48.44325, 48.441583, 48.437833, 48.442389, 
    NaN, 48.829944, 48.83075, 48.834528, 48.826583, 48.829944, NaN, 
    48.331583, 48.332389, 48.333667, 48.3295, 48.331583, NaN, 48.92, 
    48.921639, 48.921667, 48.91625, 48.92, NaN, 29.613861, 29.614139, 
    29.613306, 29.610861, 29.613861, NaN, 46.251667, 46.252472, 46.252028, 
    46.248722, 46.251667, NaN, 28.155139, 28.155361, 28.155667, 28.153472, 
    28.155139, NaN, 48.978306, 48.979111, 48.982083, 48.979167, 48.978306, 
    NaN, 48.966667, 48.9675, 48.967444, 48.963694, 48.966667, NaN, 48.932472, 
    48.932889, 48.935806, 48.930361, 48.932472, NaN, 48.903278, 48.904083, 
    48.90075, 48.8995, 48.903278, NaN, 28.667111, 28.668472, 28.667333, 
    28.665361, 28.667111, NaN, 29.984361, 29.98275, 29.98325, 29.986806, 
    29.984361, NaN, 48.671611, 48.673278, 48.674528, 48.666556, 48.671611, 
    NaN, 48.664083, 48.664944, 48.6645, 48.658694, 48.664083, NaN, 48.981556, 
    48.981972, 48.981167, 48.975333, 48.981556, NaN, 48.865833, 48.868333, 
    48.87375, 48.865389, 48.865833, NaN, 48.906667, 48.908278, 48.910417, 
    48.905, 48.906667, NaN, 28.138389, 28.1385, 28.138972, 28.136583, 
    28.138389, NaN, 32.446361, 32.446417, 32.432389, 32.438861, 32.446361, 
    NaN, 28.144194, 28.144556, 28.146056, 28.143972, 28.144194, NaN, 
    46.221639, 46.2225, 46.222083, 46.2175, 46.221639, NaN, 46.177472, 46.18, 
    46.176694, 46.174583, 46.177472, NaN, 37.727306, 37.727639, 37.729944, 
    37.72725, 37.727306, NaN, 46.264972, 46.265833, 46.258306, 46.248722, 
    46.264972, NaN, 28.139083, 28.139306, 28.138361, 28.136722, 28.139083, 
    NaN, 29.27925, 29.279222, 29.277333, 29.276639, 29.27925, NaN, 48.922472, 
    48.924139, 48.925417, 48.922528, 48.922472, NaN, 48.904167, 48.906667, 
    48.907889, 48.904972, 48.904167, NaN, 37.964972, 37.965417, 37.964944, 
    37.962056, 37.964972, NaN, 37.827528, 37.829111, 37.825833, 37.824583, 
    37.827528, NaN, 48.719111, 48.719917, 48.720778, 48.717028, 48.719111, 
    NaN, 48.569972, 48.571556, 48.571583, 48.567806, 48.569972, NaN, 
    48.864111, 48.864972, 48.868694, 48.863722, 48.864111, NaN, 48.949167, 
    48.950806, 48.952111, 48.949972, 48.949167, NaN, 48.939944, 48.940806, 
    48.941222, 48.937861, 48.939944, NaN, 47.830833, 47.831, 47.834806, 
    47.831722, 47.830833, NaN, 48.725778, 48.726583, 48.728694, 48.727417, 
    48.725778, NaN, 28.625944, 28.626556, 28.628917, 28.627333, 28.625944, 
    NaN, 48.662417, 48.663222, 48.664556, 48.662444, 48.662417, NaN, 
    45.495111, 45.494306, 45.492556, 45.494444, 45.495111, NaN, 48.851667, 
    48.852472, 48.852889, 48.849972, 48.851667, NaN, 48.531583, 48.53325, 
    48.536167, 48.53325, 48.531583, NaN, 48.639917, 48.641583, 48.642, 
    48.639083, 48.639917, NaN, 48.916611, 48.918333, 48.919583, 48.916639, 
    48.916611, NaN, 48.925806, 48.927472, 48.927472, 48.924583, 48.925806, 
    NaN, 48.840833, 48.841639, 48.841222, 48.838694, 48.840833, NaN, 
    48.894167, 48.895806, 48.897083, 48.894139, 48.894167, NaN, 48.941639, 
    48.943278, 48.944583, 48.9425, 48.941639, NaN, 48.912472, 48.914139, 
    48.911667, 48.910389, 48.912472, NaN, 48.699056, 48.699917, 48.701167, 
    48.698278, 48.699056, NaN, 47.576639, 47.578306, 47.58125, 47.574972, 
    47.576639, NaN, 33.46525, 33.466028, 33.463556, 33.461611, 33.46525, NaN, 
    48.509083, 48.5095, 48.509083, 48.506167, 48.509083, NaN, 29.730944, 
    29.729972, 29.727833, 29.730806, 29.730944, NaN, 48.326556, 48.327417, 
    48.328639, 48.326583, 48.326556, NaN, 32.4265, 32.426611, 32.4225, 
    32.421333, 32.4265, NaN, 47.888944, 47.888972, 47.885361, 47.888944, NaN, 
    29.971444, 29.971722, 29.969139, 29.971444, NaN, 29.749056, 29.749167, 
    29.746583, 29.749056, NaN, 29.162861, 29.163667, 29.160167, 29.162861, 
    NaN, 29.752278, 29.752556, 29.749972, 29.752278, NaN, 29.743444, 
    29.744028, 29.741139, 29.743444, NaN, 29.731139, 29.731889, 29.729167, 
    29.731139, NaN, 29.746139, 29.746694, 29.744222, 29.746139, NaN, 
    45.212583, 45.211833, 45.213361, 45.212583, NaN, 28.144028, 28.144194, 
    28.146556, 28.144028, NaN, 47.9945, 47.993417, 47.99, 47.9945, NaN, 
    48.421556, 48.423278, 48.421583, 48.421556, NaN, 29.742972, 29.744111, 
    29.74575, 29.742972, NaN, 29.750583, 29.750972, 29.748389, 29.750583, 
    NaN, 29.745889, 29.745889, 29.742556, 29.745889, NaN, 29.783, 29.783111, 
    29.779861, 29.783, NaN, 48.941694, 48.942472, 48.944167, 48.941694, NaN, 
    48.9075, 48.910833, 48.906639, 48.9075, NaN, 48.621583, 48.622444, 
    48.619889, 48.621583, NaN, 48.634917, 48.635778, 48.632417, 48.634917, 
    NaN, 48.841556, 48.843278, 48.840722, 48.841556, NaN, 48.36075, 
    48.363278, 48.364083, 48.36075, NaN, 47.715639, 47.715639, 47.712056, 
    47.715639, NaN, 48.915833, 48.91875, 48.917472, 48.915833, NaN, 48.935, 
    48.935806, 48.936611, 48.935, NaN, 47.864917, 47.864806, 47.860333, 
    47.864917, NaN, 46.254167, 46.255833, 46.254139, 46.254167, NaN, 
    48.860806, 48.862083, 48.859944, 48.860806, NaN, 48.894972, 48.895778, 
    48.896611, 48.894972, NaN, 48.899139, 48.9, 48.901639, 48.899139, NaN, 
    45.460583, 45.460139, 45.460722, 45.460583, NaN, 45.510361, 45.509778, 
    45.509917, 45.510361, NaN, 48.910833, 48.911639, 48.912444, 48.910833, 
    NaN, 48.901667, 48.902472, 48.9025, 48.901667, NaN, 38.75325, 38.753361, 
    38.751028, 38.75325, NaN, 48.88575, 48.887417, 48.883667, 48.88575, NaN, 
    48.88825, 48.889111, 48.886167, 48.88825, NaN, 48.91075, 48.911194, 
    48.907833, 48.91075, NaN, 48.882417, 48.883222, 48.881583, 48.882417, 
    NaN, 48.684972, 48.685778, 48.682, 48.684972, NaN, 48.649944, 48.65075, 
    48.649111, 48.649944, NaN, 37.108306, 37.110833, 37.106611, 37.108306, 
    NaN, 48.676583, 48.676972, 48.674528, 48.676583, NaN, 48.902417, 
    48.903278, 48.900778, 48.902417, NaN, 48.669056, 48.669917, 48.670806, 
    48.669056, NaN, 48.419917, 48.421583, 48.420722, 48.419917, NaN, 
    28.907472, 28.907806, 28.91325, 28.907472, NaN, 48.755778, 48.756194, 
    48.752861, 48.755778, NaN, 48.536556, 48.538278, 48.537417, 48.536556, 
    NaN, 48.846583, 48.847444, 48.846611, 48.846583, NaN, 48.807417, 
    48.808694, 48.806583, 48.807417, NaN, 48.657417, 48.658278, 48.656583, 
    48.657417, NaN, 48.575778, 48.576194, 48.573667, 48.575778, NaN, 
    48.332444, 48.333306, 48.334056, 48.332444, NaN, 48.939167, 48.939583, 
    48.939139, 48.939167, NaN, 46.159139, 46.16, 46.162083, 46.159139, NaN, 
    46.740833, 46.741639, 46.740806, 46.740833, NaN, 48.921667, 48.9225, 
    48.92375, 48.921667, NaN, 48.961667, 48.962528, 48.963278, 48.961667, 
    NaN, 29.983611, 29.984167, 29.980861, 29.983611, NaN, 29.974, 29.974278, 
    29.971694, 29.974, NaN, 37.769083, 37.768917, 37.773167, 37.769083, NaN, 
    46.2375, 46.240833, 46.239139, 46.2375, NaN, 46.227472, 46.229139, 
    46.229972, 46.227472, NaN, 29.723472, 29.723472, 29.725861, 29.723472, 
    NaN, 48.669917, 48.670778, 48.669139, 48.669917, NaN, 48.906639, 48.9075, 
    48.908306, 48.906639, NaN, 37.7675, 37.768472, 37.770944, 37.7675, NaN, 
    46.216667, 46.218306, 46.219167, 46.216667, NaN, 46.221639, 46.2225, 
    46.223333, 46.221639, NaN, 46.252472, 46.253722, 46.249583, 46.252472, 
    NaN, 45.465194, 45.463611, 45.463333, 45.465194, NaN, 47.929639, 
    47.929944, 47.933167, 47.929639, NaN, 28.867611, 28.868306, 28.866417, 
    28.867611, NaN, 29.728806, 29.7285, 29.726917, 29.728806, NaN, 47.994722, 
    47.99475, 47.998083, 47.994722, NaN, 48.903333, 48.904139, 48.9025, 
    48.903333, NaN, 48.831611, 48.83325, 48.83075, 48.831611, NaN, 48.416583, 
    48.417444, 48.415778, 48.416583, NaN, 28.251556, 28.251917, 28.255778, 
    28.251556, NaN, 48.874972, 48.876639, 48.877472, 48.874972, NaN, 28.877, 
    28.877417, 28.879167, 28.877, NaN, 38.431917, 38.431583, 38.434611, 
    38.431917, NaN, 38.683194, 38.683194, 38.680667, 38.683194, NaN, 
    38.297611, 38.297556, 38.294056, 38.297611, NaN, 33.034139, 33.035, 
    33.033333, 33.034139, NaN, 29.744917, 29.745028, 29.748333, 29.744917, 
    NaN, 46.720833, 46.722472, 46.717889, 46.720833, NaN, 30.131861, 
    30.131111, 30.128222, 30.131861, NaN, 28.767889, 28.769694, 28.767222, 
    28.767889, NaN, 48.830722, 48.831194, 48.827028, 48.830722, NaN, 
    37.763028, 37.764917, 37.76325, 37.763028, NaN, 37.964972, 37.966639, 
    37.964972, 37.964972, NaN, 29.961556, 29.962167, 29.959028, 29.961556, 
    NaN, 29.727722, 29.726861, 29.728056, 29.727722, NaN, 29.605639, 
    29.606528, 29.604222, 29.605639, NaN, 48.651583, 48.652861, 48.65075, 
    48.651583, NaN, 48.908306, 48.909167, 48.908333, 48.908306, NaN, 
    48.36825, 48.368694, 48.367417, 48.36825, NaN, 33.037528, 33.038333, 
    33.038306, 33.037528, NaN, 48.426611, 48.427389, 48.426611, 48.426611, 
    NaN, 48.679111, 48.68075, 48.678278, 48.679111, NaN, 48.428278, 
    48.429056, 48.427417, 48.428278, NaN, 48.842417, 48.843667, 48.841556, 
    48.842417, NaN, 48.73325, 48.734111, 48.732444, 48.73325, NaN, 48.809917, 
    48.810778, 48.809944, 48.809917, NaN, 48.899056, 48.8995, 48.897028, 
    48.899056, NaN, 48.175806, 48.176667, 48.174944, 48.175806, NaN, 
    48.173306, 48.174972, 48.174167, 48.173306, NaN, 48.774111, 48.776639, 
    48.775833, 48.774111, NaN, 48.919972, 48.921611, 48.920833, 48.919972, 
    NaN, 48.854972, 48.855833, 48.855, 48.854972, NaN, 48.996694, 48.998278, 
    48.996639, 48.996694, NaN, 48.830806, 48.831667, 48.829528, 48.830806, 
    NaN, 48.925778, 48.926639, 48.927889, 48.925778, NaN, 48.919972, 
    48.920417, 48.919972, 48.919972, NaN, 48.8925, 48.893278, 48.891639, 
    48.8925, NaN, 48.871639, 48.874167, 48.873333, 48.871639, NaN, 46.300861, 
    46.301667, 46.301611, 46.300861, NaN, 29.950861, 29.951889, 29.951528, 
    29.950861, NaN, 29.976167, 29.976722, 29.974444, 29.976167, NaN, 
    29.748667, 29.748306, 29.7485, 29.748667, NaN, 45.076333, 45.077833, 
    45.078833, 45.076333, NaN, 45.806944, 45.805389, 45.807861, 45.806944, 
    NaN, 28.309889, 28.310111, 28.309917, 28.309889, NaN, 48.916639, 
    48.917028, 48.910333, 48.916639, NaN, 28.293361, 28.293611, 28.293111, 
    28.293361, NaN, 28.312444, 28.312611, 28.31075, 28.312444, NaN, 28.309, 
    28.309306, 28.308917, 28.309, NaN, 28.307361, 28.307611, 28.307278, 
    28.307361, NaN, 28.314806, 28.315028, 28.314389, 28.314806, NaN, 
    28.141556, 28.141722, 28.141806, 28.141556, NaN, 28.310694, 28.310972, 
    28.310667, 28.310694, NaN, 28.298417, 28.298583, 28.298194, 28.298417, 
    NaN, 28.299028, 28.299444, 28.298833, 28.299028, NaN, 29.747389, 
    29.748528, 29.746778, 29.747389, NaN, 48.852417, 48.853278, 48.849111, 
    48.852417, NaN, 28.094056, 28.094222, 28.093806, 28.094056, NaN, 
    28.306361, 28.306583, 28.306722, 28.306361, NaN, 28.308111, 28.308556, 
    28.308083, 28.308111, NaN, 28.144028, 28.144194, 28.142667, 28.144028, 
    NaN, 37.9, 37.900778, 37.900778, 37.9, NaN, 46.743306, 46.745444, 
    46.743278, 46.743306, NaN, 46.739972, 46.740833, 46.740806, 46.739972, 
    NaN, 48.929944, 48.930417, 48.929139, 48.929944, NaN, 48.896639, 
    48.897056, 48.895417, 48.896639, NaN, 48.592444, 48.593222, 48.591611, 
    48.592444, NaN, 48.669917, 48.670778, 48.670778, 48.669917, NaN, 
    48.744944, 48.74575, 48.744944, 48.744944, NaN, 48.969083, 48.969472, 
    48.967, 48.969083, NaN, 48.434972, 48.43575, 48.43575, 48.434972, NaN, 
    48.419889, 48.420361, 48.418694, 48.419889, NaN, 28.318194, 28.318417, 
    28.319028, 28.318194, NaN, 28.304833, 28.305, 28.30475, 28.304833, NaN, 
    48.657444, 48.65825, 48.657444, 48.657444, NaN, 48.891583, 48.892, 
    48.8895, 48.891583, NaN, 48.892444, 48.892861, 48.8895, 48.892444, NaN, 
    48.869972, 48.870389, 48.869972, 48.869972, NaN, 28.05225, 28.052583, 
    28.053778, 28.05225, NaN, 28.145556, 28.145722, 28.145667, 28.145556, 
    NaN, 28.154111, 28.154278, 28.154194, 28.154111, NaN, 28.100361, 
    28.100611, 28.100833, 28.100361, NaN, 28.051944, 28.052194, 28.051389, 
    28.051944, NaN, 28.144806, 28.144972, 28.147, 28.144806, NaN, 28.151389, 
    28.151556, 28.151417, 28.151389, NaN, 28.106667, 28.106972, 28.106389, 
    28.106667, NaN ;
}
