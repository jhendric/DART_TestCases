netcdf f3coerr {
dimensions:
	local_time = 25 ;
	latitude = 37 ;
	altitude = 15 ;
variables:
	float altitude(altitude) ;
		altitude:units = "km" ;
	float latitude(latitude) ;
		latitude:long_name = "local time of day" ;
		latitude:units = "degrees" ;
	float local_time(local_time) ;
		local_time:units = "hours" ;
	float percent(local_time, latitude, altitude) ;
		percent:usage = "observation_error_variance = max(some_floor, percent(k,j,t)*observation_value)" ;

// global attributes:
		:supporting_material_1 = "X. Yue et. al; 2010 https://www.ann-geophys.net/28/217/2010" ;
		:supporting_material_2 = "J. Y. Liu et. al; 2010 doi:10.1029/2009JA015079" ;
data:

 altitude = 100, 150, 200, 250, 300, 350, 400, 450, 500, 550, 600, 650, 700, 
    750, 800 ;

 latitude = -90, -85, -80, -75, -70, -65, -60, -55, -50, -45, -40, -35, -30, 
    -25, -20, -15, -10, -5, 0, 5, 10, 15, 20, 25, 30, 35, 40, 45, 50, 55, 60, 
    65, 70, 75, 80, 85, 90 ;

 local_time = 0, 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12, 13, 14, 15, 16, 17, 
    18, 19, 20, 21, 22, 23, 24 ;

 percent =
  -375.714, -499.778, -499.788, -749.25, -686.83, -499.565, -499.499, 
    -499.493, -499.539, -499.519, -499.51, -499.469, -749.25, -749.25, 
    -561.938,
  -0.284, -0.452, -0.493, -249.821, -187.384, -0.115, -0.082, -0.083, -0.091, 
    -0.032, -0.011, 0.045, -249.712, -249.733, -187.373,
  0.781, 0.309, 0.123, 0.042, 0.02, -0.023, -0.026, -0.053, -0.079, -0.092, 
    -0.096, -0.116, -0.1, -0.097, -0.087,
  3.178, 1.004, 0.909, 0.201, 0.091, 0.088, 0.065, 0.065, 0.07, 0.037, 0.032, 
    -0.005, -0.045, -0.047, -0.048,
  3.887, 1.08, 0.945, 0.198, 0.092, 0.079, 0.085, 0.081, 0.07, 0.066, 0.057, 
    0.039, 0.016, -0.031, -0.066,
  4.141, 1.343, 1.179, 0.233, 0.106, 0.095, 0.095, 0.091, 0.085, 0.072, 
    0.058, 0.025, 0.003, -0.018, -0.054,
  4.936, 1.536, 1.263, 0.275, 0.113, 0.103, 0.096, 0.095, 0.091, 0.076, 
    0.064, 0.052, 0.021, -0.027, -0.065,
  4.215, 1.372, 1.081, 0.223, 0.09, 0.08, 0.085, 0.078, 0.07, 0.059, 0.038, 
    0.018, -0.002, -0.018, -0.048,
  3.095, 1.049, 0.737, 0.146, 0.056, 0.043, 0.034, 0.028, 0.021, 0.011, 
    0.002, -0.012, -0.027, -0.044, -0.037,
  3.168, 0.895, 0.702, 0.113, 0.034, 0.027, 0.023, 0.025, 0.023, 0.018, 
    0.017, 0.002, -0.024, -0.039, -0.057,
  2.612, 0.897, 0.593, 0.096, 0.019, 0.015, 0.014, 0.005, -0.001, -0.01, 
    -0.016, -0.029, -0.039, -0.032, -0.023,
  5.035, 1.509, 0.874, 0.145, 0.034, 0.009, 0.01, 0.005, -0.003, -0.007, 
    -0.009, -0.009, -0.001, -0.004, 0.034,
  8.182, 2.498, 1.436, 0.195, 0.056, 0.043, 0.037, 0.023, 0.02, 0.03, 0.029, 
    0.022, 0.028, 0.053, 0.03,
  9.827, 3.695, 1.801, 0.311, 0.102, 0.085, 0.079, 0.071, 0.067, 0.056, 
    0.051, 0.05, 0.049, 0.037, 0.017,
  8.839, 3.665, 1.929, 0.352, 0.137, 0.114, 0.097, 0.084, 0.075, 0.073, 
    0.063, 0.056, 0.046, 0.031, 0.022,
  5.052, 2.792, 1.377, 0.246, 0.094, 0.074, 0.06, 0.063, 0.058, 0.03, 0.037, 
    0.032, 0.036, 0.055, 0.031,
  -0.489, -0.375, -0.124, -0.055, -0.032, -0.021, -0.001, -0.005, -0.021, 
    0.004, 0.022, -0.016, -0.009, -0.006, 0.013,
  -7.133, -1.836, -0.404, -0.056, -0.019, -0.013, -0.021, -0.018, -0.011, 
    -0.022, -0.013, -0.019, -0.01, 0.03, 0.046,
  -2.834, -1.441, -0.323, -0.077, -0.035, -0.02, -0.031, -0.036, -0.039, 
    -0.027, -0.024, -0.004, 0.021, 0.045, 0.014,
  -6.271, -1.918, -0.682, -0.145, -0.068, -0.074, -0.089, -0.09, -0.083, 
    -0.066, -0.043, -0.023, -0.004, -0.006, -0.012,
  -2.943, -1.032, -0.136, -0.018, -0.024, -0.024, -0.021, -0.019, -0.025, 
    -0.035, -0.025, -0.018, -0.027, -0.019, -0.029,
  1.143, 1.145, 1.008, 0.283, 0.119, 0.098, 0.082, 0.067, 0.056, 0.045, 
    0.032, 0.021, 0.011, -0.037, -0.026,
  7.162, 3.615, 1.468, 0.27, 0.094, 0.077, 0.07, 0.061, 0.054, 0.058, 0.046, 
    0.036, 0.008, -0.044, -0.017,
  4.635, 1.673, 1.014, 0.237, 0.068, 0.058, 0.061, 0.069, 0.071, 0.064, 
    0.057, 0.039, 0.011, -0.055, 0.011,
  3.16, 1.501, 0.947, 0.146, 0.039, 0.02, 0.02, 0.014, 0.014, -0.002, -0.003, 
    -0.011, -0.027, -0.032, 0.006,
  1.424, 0.299, 0.061, -0.035, -0.029, -0.024, -0.02, -0.023, -0.024, -0.032, 
    -0.024, -0.02, -0.034, -0.031, 0.019,
  0.478, -0.023, -0.158, -0.027, -0.015, -0.025, -0.033, -0.04, -0.048, 
    -0.041, -0.04, -0.05, -0.041, -0.01, -0.011,
  0.592, 0.036, 0.031, -0.002, -0.004, 0.001, 0.002, -0.003, -0.014, -0.026, 
    -0.021, -0.011, -0.018, -0.012, -0.047,
  2.905, 0.917, 0.59, 0.11, 0.044, 0.036, 0.03, 0.027, 0.029, 0.029, 0.026, 
    0.017, 0.006, 0.005, -0.071,
  5.623, 1.552, 1.087, 0.207, 0.094, 0.091, 0.091, 0.087, 0.071, 0.06, 0.05, 
    0.029, 0.01, 0.01, -0.073,
  5.288, 1.649, 1.092, 0.204, 0.099, 0.092, 0.095, 0.092, 0.086, 0.099, 
    0.101, 0.06, 0.02, -0.029, -0.18,
  3.799, 0.745, 0.619, 0.166, 0.085, 0.076, 0.077, 0.081, 0.092, 0.09, 0.067, 
    0.027, 0.013, -0.033, -0.232,
  1.967, 0.522, 0.531, 0.161, 0.095, 0.082, 0.085, 0.087, 0.077, 0.059, 
    0.039, -0.008, -0.031, -0.087, -0.014,
  1.378, 0.415, 0.198, 0.079, 0.065, 0.065, 0.059, 0.052, 0.042, 0.044, 
    0.016, 0.063, 0.021, 0.054, -125.047,
  0.538, 0.111, -0.015, -0.015, 0.006, -0.012, -0.016, -0.007, 0.012, 0.023, 
    -0.017, 0.017, 0.001, 0.016, -249.782,
  -187.774, -249.942, -249.764, -62.47, -0.033, -0.033, -0.03, -0, -0.029, 
    -0.042, -0.104, -0.16, -0.159, -62.69, -686.801,
  -561.938, -749.25, -749.25, -561.945, -499.516, -499.513, -499.509, 
    -499.505, -499.499, -499.492, -499.511, -499.527, -0.239, -561.998, 
    -561.938,
  -374.417, 0.36, 0.24, 0.064, 0.01, 0.016, 0.01, -374.622, 0.039, 0.022, 
    -124.823, -499.494, -499.496, -499.599, -561.938,
  0.626, 0.07, -0.114, -0.082, -0.061, -0.061, -0.05, -0.034, -0.014, 0.004, 
    -0.018, -0.036, -0.017, -0.118, -187.33,
  0.207, -0.053, -0.319, -0.098, -0.068, -0.073, -0.087, -0.097, -0.132, 
    -0.156, -0.128, -0.069, -0.035, -0.019, 0.02,
  2.094, 0.551, 0.416, 0.05, 0.02, 0.02, 0.039, 0.032, 0.021, 0.01, 0.002, 
    -0.009, -0.035, 0.009, 0.016,
  3.005, 0.844, 0.768, 0.161, 0.073, 0.075, 0.067, 0.061, 0.057, 0.047, 
    0.031, 0.011, -0.013, -0.03, -0.05,
  3.881, 1.188, 1.062, 0.227, 0.104, 0.094, 0.092, 0.094, 0.09, 0.082, 0.067, 
    0.048, 0.02, -0.012, -0.06,
  4.178, 1.317, 1.088, 0.205, 0.086, 0.082, 0.089, 0.091, 0.089, 0.075, 
    0.061, 0.038, 0.014, -0.019, -0.065,
  3.599, 1.134, 0.909, 0.175, 0.072, 0.071, 0.068, 0.068, 0.057, 0.05, 0.039, 
    0.029, 0.012, -0.017, -0.045,
  3.203, 1.066, 0.97, 0.198, 0.076, 0.068, 0.07, 0.071, 0.069, 0.06, 0.058, 
    0.035, 0.011, -0.013, -0.033,
  3.145, 0.981, 0.702, 0.131, 0.049, 0.042, 0.039, 0.034, 0.033, 0.03, 0.022, 
    0.013, 0.001, 0.002, 0.007,
  2.207, 0.683, 0.408, 0.073, 0.02, 0.013, 0.016, 0.015, 0.014, 0.007, 0.004, 
    0.003, 0.008, 0.016, 0.014,
  2.532, 0.767, 0.449, 0.07, 0.02, 0.013, 0.008, 0.006, 0.006, 0.006, 0.014, 
    0.015, 0.017, 0.014, 0.009,
  3.714, 1.111, 0.524, 0.068, 0.025, 0.024, 0.024, 0.027, 0.025, 0.031, 
    0.028, 0.025, 0.024, 0.03, 0.035,
  5.083, 1.907, 0.979, 0.148, 0.054, 0.044, 0.045, 0.039, 0.041, 0.036, 
    0.032, 0.033, 0.037, 0.035, 0.024,
  5.004, 2.245, 1.15, 0.205, 0.083, 0.064, 0.057, 0.054, 0.054, 0.045, 0.042, 
    0.034, 0.033, 0.025, 0.024,
  3.441, 1.367, 0.582, 0.108, 0.045, 0.036, 0.03, 0.031, 0.025, 0.025, 0.026, 
    0.027, 0.029, 0.036, 0.027,
  -0.258, -0.226, -0.114, -0.047, -0.025, -0.026, -0.034, -0.032, -0.038, 
    -0.029, -0.026, -0.021, -0.016, -0.001, 0.026,
  -4.648, -1.593, -0.352, -0.068, -0.036, -0.031, -0.019, -0.018, -0.012, 
    -0.023, -0.024, -0.018, -0.009, 0.001, 0.027,
  -7.922, -2.264, -0.442, -0.067, -0.032, -0.006, -0.001, -0.007, -0.017, 
    -0.018, -0.023, -0.013, -0.004, 0.011, 0.02,
  -5.038, -2.158, -0.569, -0.132, -0.072, -0.073, -0.086, -0.092, -0.098, 
    -0.094, -0.071, -0.065, -0.047, -0.031, 0.003,
  -3.149, -1.269, -0.345, -0.057, -0.037, -0.034, -0.04, -0.042, -0.042, 
    -0.037, -0.039, -0.037, -0.035, -0.026, -0.06,
  0.159, 0.387, 0.236, 0.073, 0.042, 0.039, 0.039, 0.043, 0.051, 0.037, 
    0.026, 0.02, 0.006, -0.009, -0.096,
  3.703, 2.17, 1.198, 0.183, 0.08, 0.069, 0.072, 0.071, 0.072, 0.071, 0.05, 
    0.032, 0.006, -0.04, -0.159,
  2.997, 0.97, 0.441, 0.07, 0.018, 0.015, 0.015, 0.012, 0.008, 0.002, -0.006, 
    -0.008, -0.027, -0.058, -0.089,
  0.33, 0.145, -0.006, -0.033, -0.026, -0.025, -0.02, -0.016, -0.014, -0.012, 
    -0.016, -0.027, -0.05, -0.054, -0.042,
  -1.252, -0.445, -0.349, -0.087, -0.04, -0.036, -0.041, -0.048, -0.054, 
    -0.059, -0.057, -0.051, -0.046, -0.027, -0.076,
  -0.344, -0.269, -0.151, -0.043, -0.023, -0.03, -0.034, -0.039, -0.043, 
    -0.044, -0.043, -0.037, -0.035, -0.009, -0.053,
  1.634, 0.491, 0.328, 0.065, 0.013, 0.009, 0.005, 0.002, -0.003, -0.007, 
    -0.004, -0.002, -0.004, -0, -0.055,
  4.662, 1.494, 1.3, 0.288, 0.096, 0.074, 0.067, 0.061, 0.052, 0.043, 0.03, 
    0.016, 0, -0.003, -0.058,
  6.742, 1.891, 1.615, 0.332, 0.128, 0.105, 0.1, 0.089, 0.08, 0.076, 0.077, 
    0.056, 0.029, -0.021, -0.105,
  5.961, 1.647, 1.402, 0.365, 0.159, 0.142, 0.145, 0.151, 0.135, 0.129, 
    0.111, 0.084, 0.045, 0.001, -0.121,
  3.285, 0.837, 0.685, 0.23, 0.118, 0.105, 0.102, 0.103, 0.104, 0.095, 0.076, 
    0.061, 0.028, -0.001, -0.073,
  3.223, 0.598, 0.392, 0.128, 0.081, 0.077, 0.074, 0.078, 0.069, 0.071, 
    0.065, 0.073, 0.032, 0.015, -0.053,
  1.406, 0.319, 0.193, 0.093, 0.061, 0.067, 0.077, 0.081, 0.091, 0.091, 
    0.109, 0.123, 0.092, 0.129, -0.119,
  0.989, -0, -0.028, -0.006, -0.002, 0.004, 0.008, 0.009, 0.029, 0.021, 
    0.002, -0.006, -0.007, -0.085, -125.125,
  -0.942, -0.331, -0.187, -0.095, -0.06, -0.066, -0.083, -0.079, -0.081, 
    -0.093, -0.098, -0.086, -62.492, -0.159, -686.818,
  -374.986, -499.621, -499.521, -499.509, -499.509, -499.514, -499.559, 
    -499.543, -499.523, -374.65, -124.907, -499.503, -561.911, -499.616, 
    -561.938,
  -375.136, -499.695, -499.694, -499.543, -499.522, -499.526, -374.649, 
    -0.063, -0.056, -0.048, -0.054, -499.487, -499.528, -374.657, -187.361,
  -1.012, -0.419, -0.556, -0.16, -0.085, -0.082, -0.093, -0.092, -0.087, 
    -0.072, -0.061, -0.079, -0.04, -0.026, -187.289,
  -0.049, -0.161, -0.338, -0.087, -0.075, -0.087, -0.107, -0.135, -0.134, 
    -0.157, -0.166, -0.143, -0.079, -0.041, 0.01,
  2.192, 0.548, 0.411, 0.047, 0.031, 0.001, 0.006, 0.004, -0.02, -0.045, 
    -0.043, -0.075, -0.104, -0.138, -0.127,
  2.716, 0.77, 0.622, 0.124, 0.054, 0.057, 0.05, 0.041, 0.029, 0.011, -0.015, 
    -0.05, -0.065, -0.089, -0.138,
  3.221, 0.976, 0.816, 0.159, 0.079, 0.071, 0.074, 0.069, 0.063, 0.049, 
    0.032, 0.005, -0.024, -0.055, -0.12,
  3.628, 1.105, 0.915, 0.177, 0.085, 0.079, 0.078, 0.077, 0.076, 0.068, 
    0.051, 0.039, 0.012, -0.005, -0.078,
  2.845, 0.947, 0.8, 0.157, 0.071, 0.066, 0.066, 0.067, 0.061, 0.052, 0.039, 
    0.019, -0.003, -0.019, -0.061,
  3.155, 1.085, 0.864, 0.156, 0.064, 0.061, 0.064, 0.064, 0.067, 0.063, 0.05, 
    0.037, 0.012, -0.011, -0.035,
  1.716, 0.629, 0.467, 0.095, 0.041, 0.037, 0.038, 0.038, 0.034, 0.034, 0.03, 
    0.024, 0.004, -0.004, -0.006,
  0.151, 0.037, 0.027, 0.009, -0.004, -0.004, -0.005, -0.005, -0.007, -0.012, 
    -0.011, -0.009, -0.007, 0.012, 0.044,
  -1.316, -0.573, -0.38, -0.072, -0.035, -0.033, -0.029, -0.028, -0.023, 
    -0.016, -0.007, 0.008, 0.019, 0.045, 0.038,
  -2.304, -0.929, -0.606, -0.119, -0.061, -0.052, -0.051, -0.044, -0.032, 
    -0.022, -0.013, -0.004, 0.015, 0.03, 0.045,
  -1.137, -0.398, -0.247, -0.058, -0.027, -0.019, -0.014, -0.008, -0.007, 
    -0.001, 0.002, 0.012, 0.024, 0.039, 0.054,
  -0.484, 0.003, 0.078, 0.016, 0, -0.004, -0.002, 0.004, 0.008, 0.01, 0.021, 
    0.026, 0.036, 0.048, 0.051,
  -1.629, -0.273, 0.017, 0.002, 0.004, 0.001, -0.005, -0.005, -0.006, -0.003, 
    0.001, 0.006, 0.01, 0.019, 0.066,
  -4.731, -1.757, -0.59, -0.118, -0.075, -0.077, -0.074, -0.073, -0.065, 
    -0.06, -0.054, -0.045, -0.028, 0.022, 0.032,
  -6.229, -1.934, -0.543, -0.103, -0.064, -0.052, -0.06, -0.06, -0.052, 
    -0.049, -0.041, -0.024, 0.013, 0.024, 0.019,
  -8.001, -2.457, -0.514, -0.058, -0.03, -0.026, -0.014, -0.018, -0.022, 
    -0.015, -0.012, 0.004, 0.016, 0.022, 0.049,
  -5.602, -1.781, -0.452, -0.082, -0.053, -0.05, -0.053, -0.048, -0.047, 
    -0.047, -0.045, -0.056, -0.054, -0.042, -0.009,
  -2.214, -0.835, -0.214, -0.035, -0.014, -0.016, -0.014, -0.025, -0.033, 
    -0.035, -0.033, -0.035, -0.042, -0.057, -0.027,
  -1.323, 0.213, 0.308, 0.061, 0.043, 0.051, 0.052, 0.056, 0.041, 0.048, 
    0.038, 0.026, 0.017, -0.013, -0.068,
  2.031, 1.083, 0.448, 0.073, 0.039, 0.029, 0.023, 0.02, 0.032, 0.025, 0.036, 
    0.038, 0.019, -0.025, -0.086,
  0.829, 0.324, 0.142, 0.019, 0.006, 0.009, 0.01, 0.024, 0.026, 0.019, 0.004, 
    -0.009, -0.026, -0.059, -0.064,
  -2.31, -0.934, -0.562, -0.119, -0.053, -0.049, -0.04, -0.044, -0.044, 
    -0.052, -0.055, -0.058, -0.069, -0.078, -0.067,
  -1.852, -0.677, -0.589, -0.151, -0.071, -0.065, -0.075, -0.081, -0.081, 
    -0.074, -0.065, -0.061, -0.057, -0.041, -0.013,
  0.577, 0.142, 0.138, 0, -0.024, -0.032, -0.033, -0.037, -0.045, -0.044, 
    -0.047, -0.04, -0.032, -0.003, -0.075,
  2.867, 0.945, 0.813, 0.176, 0.048, 0.03, 0.016, 0.007, 0.003, -0.004, 
    0.002, 0.002, -0.005, 0.001, -0.072,
  5.496, 1.491, 1.529, 0.346, 0.097, 0.071, 0.067, 0.057, 0.043, 0.045, 
    0.037, 0.03, 0.018, 0.002, -0.11,
  7.174, 2.099, 2.075, 0.484, 0.159, 0.129, 0.124, 0.115, 0.105, 0.091, 
    0.071, 0.047, 0.024, -0.003, -0.107,
  6.213, 1.816, 1.799, 0.473, 0.173, 0.15, 0.143, 0.135, 0.125, 0.108, 0.096, 
    0.069, 0.035, -0.012, -0.126,
  4.903, 1.048, 0.899, 0.294, 0.141, 0.128, 0.126, 0.114, 0.098, 0.082, 
    0.053, 0.019, -0.01, -0.062, -0.119,
  4.491, 1.086, 0.766, 0.215, 0.093, 0.084, 0.078, 0.085, 0.087, 0.076, 
    0.058, 0.053, 0.026, 0.013, -0.154,
  2.155, 0.409, 0.225, 0.054, 0.021, 0.024, 0.036, 0.041, 0.044, 0.048, 
    0.057, 0.036, 0.048, 0.046, -0.003,
  1.285, 0.173, 0.025, 0.003, 0.013, 0.028, 0.047, 0.056, 0.063, 0.058, 
    0.061, 0.048, 0.085, 0.162, -124.854,
  0.538, -0.025, -0.205, -0.098, -0.043, -0.039, -0.033, -0.01, 0.011, 0.028, 
    0.056, 0.112, -249.638, -249.683, -686.823,
  -375.02, -499.623, -499.654, -499.55, -499.522, -499.517, -0.035, -0.021, 
    -499.503, -499.496, -499.481, -499.458, -749.25, -749.25, -561.938,
  1.021, -124.695, -499.507, -499.506, -374.62, 0.017, 0.017, 0.018, -499.49, 
    -499.482, -499.517, -499.542, -499.529, -499.528, -374.625,
  1.372, 0.289, -0.054, -0.119, -0.071, -0.1, -0.107, -0.112, -0.087, -0.05, 
    -0.038, -0.032, 0, -0.001, -0.002,
  1.289, 0.227, 0.164, 0.037, 0.007, -0.004, -0.03, -0.033, -0.041, -0.056, 
    -0.022, 0.004, -0.003, -0.015, 0.032,
  2.547, 0.759, 0.631, 0.122, 0.079, 0.079, 0.074, 0.058, 0.046, 0.004, 
    -0.052, -0.061, -0.052, -0.053, -0.067,
  2.309, 0.666, 0.637, 0.122, 0.067, 0.067, 0.066, 0.063, 0.045, 0.036, 0.04, 
    0.011, -0.035, -0.052, -0.086,
  2.776, 0.894, 0.803, 0.152, 0.083, 0.077, 0.078, 0.08, 0.087, 0.076, 0.059, 
    0.044, 0.028, 0.012, -0.07,
  3.486, 1.131, 1.031, 0.189, 0.096, 0.091, 0.091, 0.089, 0.083, 0.078, 
    0.062, 0.037, -0.003, -0.033, -0.079,
  2.981, 0.899, 0.752, 0.152, 0.072, 0.068, 0.071, 0.073, 0.075, 0.065, 
    0.043, 0.022, -0.005, -0.038, -0.076,
  1.587, 0.518, 0.428, 0.078, 0.034, 0.035, 0.037, 0.035, 0.029, 0.025, 
    0.026, 0.009, -0.009, -0.029, -0.054,
  0.386, 0.173, 0.157, 0.028, 0.008, 0.007, 0.007, 0.008, 0.006, 0.003, 
    -0.009, -0.018, -0.031, -0.05, -0.047,
  -1.294, -0.381, -0.218, -0.043, -0.022, -0.021, -0.023, -0.022, -0.025, 
    -0.023, -0.024, -0.018, -0.019, -0.019, -0.013,
  -3.319, -1.263, -0.794, -0.135, -0.067, -0.061, -0.057, -0.055, -0.05, 
    -0.046, -0.039, -0.037, -0.03, -0.018, 0.005,
  -3.823, -1.42, -0.875, -0.161, -0.078, -0.073, -0.075, -0.076, -0.073, 
    -0.069, -0.064, -0.052, -0.044, -0.03, -0.002,
  -3.421, -1.249, -0.726, -0.133, -0.071, -0.067, -0.066, -0.063, -0.059, 
    -0.055, -0.048, -0.042, -0.025, -0.009, 0.014,
  -2.581, -0.85, -0.325, -0.054, -0.032, -0.03, -0.032, -0.037, -0.035, 
    -0.032, -0.025, -0.014, -0.002, 0.014, 0.032,
  -3.249, -0.702, -0.246, -0.032, -0.025, -0.035, -0.046, -0.05, -0.049, 
    -0.044, -0.039, -0.022, -0.004, 0.029, 0.051,
  -3.093, -1.5, -0.643, -0.14, -0.083, -0.085, -0.079, -0.071, -0.069, 
    -0.068, -0.06, -0.058, -0.04, -0.026, -0.011,
  -4.867, -1.596, -0.464, -0.08, -0.063, -0.054, -0.049, -0.052, -0.044, 
    -0.044, -0.037, -0.041, -0.027, -0.025, -0.011,
  -5.359, -1.52, -0.272, -0.015, -0.007, -0.019, -0.024, -0.024, -0.03, 
    -0.021, -0.006, -0.01, 0.009, 0.001, -0.003,
  -0.703, -0.541, -0.276, -0.042, -0.026, -0.026, -0.029, -0.032, -0.039, 
    -0.054, -0.057, -0.074, -0.063, -0.118, -0.061,
  1.006, 0.229, 0.016, 0.008, 0.014, 0.017, 0.008, 0, 0.001, -0.011, -0.037, 
    -0.05, -0.078, -0.126, -0.08,
  -0.438, 0.192, 0.27, 0.053, 0.043, 0.047, 0.051, 0.05, 0.042, 0.036, 0.014, 
    0.001, -0.021, -0.097, -0.078,
  0.248, 0.323, 0.153, 0.014, 0.008, 0.002, 0.004, 0.009, 0.007, 0, -0.003, 
    -0.014, -0.05, -0.105, -0.091,
  -0.464, -0.225, -0.111, -0.043, -0.024, -0.017, -0.008, -0.005, 0.004, 
    0.003, -0.005, -0.024, -0.054, -0.098, 0.021,
  -2.136, -0.856, -0.688, -0.16, -0.068, -0.06, -0.065, -0.072, -0.086, 
    -0.094, -0.077, -0.07, -0.059, -0.032, 0.05,
  -1.279, -0.61, -0.54, -0.14, -0.073, -0.072, -0.07, -0.073, -0.071, -0.069, 
    -0.063, -0.049, -0.035, 0, 0.022,
  0.748, 0.189, 0.172, 0.028, -0.009, -0.02, -0.029, -0.035, -0.037, -0.034, 
    -0.033, -0.024, -0.019, 0.002, -0.008,
  3.423, 1.049, 0.986, 0.211, 0.058, 0.045, 0.037, 0.033, 0.027, 0.014, 
    0.004, 0.002, -0.019, 0.002, -0.014,
  5.511, 1.504, 1.492, 0.324, 0.107, 0.092, 0.093, 0.087, 0.086, 0.085, 0.08, 
    0.063, 0.046, -0.009, -0.052,
  7.162, 2.004, 2.184, 0.507, 0.174, 0.158, 0.15, 0.149, 0.139, 0.126, 0.114, 
    0.09, 0.051, -0.007, -0.021,
  6.303, 1.712, 1.65, 0.434, 0.186, 0.17, 0.165, 0.16, 0.155, 0.139, 0.113, 
    0.076, 0.032, -0.033, -0.077,
  4.112, 0.912, 0.816, 0.262, 0.145, 0.126, 0.132, 0.134, 0.128, 0.116, 
    0.096, 0.061, 0.022, -0.015, -0.104,
  3.442, 0.871, 0.715, 0.213, 0.112, 0.116, 0.106, 0.105, 0.099, 0.092, 
    0.087, 0.074, 0.057, 0.032, -0.079,
  2.21, 0.457, 0.395, 0.102, 0.048, 0.046, 0.052, 0.049, 0.055, 0.06, 0.052, 
    0.05, 0.055, 0.052, 0.016,
  0.795, 0.14, 0.051, 0.003, -0.008, -0.009, -0.01, -0.003, -0.002, -0.005, 
    -0.006, 0.013, 0.014, 0.061, -0.023,
  -0.037, -0.039, -0.101, -0.075, -0.056, -0.051, -0.043, -0.032, -0.029, 
    -0.016, 0.002, -0.028, -0.035, -249.77, -561.921,
  -0.727, -0.192, -0.096, -499.515, -499.509, -499.508, -499.512, -499.524, 
    -499.534, -499.535, -499.535, -499.545, -499.535, -749.25, -561.938,
  -1.764, -0.68, -0.704, -0.121, -499.514, -499.512, -499.512, -499.473, 
    -499.456, -499.453, -499.449, -749.25, -749.25, -749.25, -561.938,
  1.544, 0.342, 0.204, 0.001, 0.001, 0.012, 0.023, 0.019, 0.022, 0.039, 
    0.047, -249.699, -249.689, -249.639, -187.268,
  1.176, 0.167, 0.169, 0.006, 0.011, 0.02, 0.022, 0.031, 0.035, 0.018, 0.022, 
    0.007, 0.03, 0.059, -0.033,
  2.728, 0.772, 0.637, 0.101, 0.049, 0.039, 0.045, 0.024, 0.022, 0.029, 
    0.025, 0.023, 0.031, -0.003, -0.064,
  3.152, 0.927, 0.857, 0.168, 0.104, 0.097, 0.077, 0.07, 0.058, 0.041, 0.014, 
    0.001, -0.029, -0.033, -0.056,
  3.282, 0.944, 0.86, 0.178, 0.098, 0.097, 0.093, 0.085, 0.081, 0.076, 0.073, 
    0.064, 0.039, 0.033, -0.06,
  3.205, 0.93, 0.853, 0.156, 0.075, 0.066, 0.061, 0.054, 0.051, 0.046, 0.035, 
    0.024, -0.001, -0.017, -0.045,
  2.688, 0.773, 0.717, 0.13, 0.06, 0.059, 0.057, 0.056, 0.051, 0.047, 0.039, 
    0.019, 0.001, -0.013, -0.038,
  1.792, 0.57, 0.507, 0.094, 0.048, 0.045, 0.047, 0.047, 0.05, 0.045, 0.031, 
    0.017, -0.002, -0.023, -0.044,
  0.406, 0.207, 0.207, 0.032, 0.017, 0.023, 0.028, 0.026, 0.022, 0.014, 
    0.008, -0.008, -0.023, -0.026, -0.061,
  -0.482, -0.149, -0.158, -0.043, -0.027, -0.029, -0.031, -0.03, -0.032, 
    -0.026, -0.024, -0.018, -0.015, -0.024, -0.033,
  -2.372, -0.886, -0.64, -0.126, -0.074, -0.066, -0.06, -0.056, -0.053, 
    -0.05, -0.042, -0.028, -0.025, -0.01, -0.003,
  -3.096, -1.163, -0.782, -0.14, -0.075, -0.072, -0.071, -0.067, -0.064, 
    -0.062, -0.054, -0.041, -0.039, -0.027, 0.005,
  -1.562, -0.598, -0.404, -0.079, -0.052, -0.052, -0.053, -0.053, -0.047, 
    -0.041, -0.042, -0.041, -0.019, 0.01, 0.049,
  0.81, 0.33, 0.192, 0.033, 0.017, 0.009, -0.001, -0.018, -0.021, -0.015, 
    -0.018, 0.001, 0.006, 0.002, 0.007,
  0.865, 0.329, 0.218, 0.055, 0.031, 0.027, 0.015, 0.01, -0.001, -0.018, 
    -0.028, -0.044, -0.031, -0.035, -0.02,
  2.116, 0.707, 0.291, 0.038, 0.02, -0.001, -0.02, -0.036, -0.052, -0.055, 
    -0.062, -0.053, -0.042, -0.084, -0.085,
  1.516, 0.331, 0.067, -0.013, -0.003, -0.007, -0.012, -0.009, -0.009, 
    -0.026, -0.049, -0.107, -0.121, -0.176, -0.128,
  3.292, 1.067, 0.515, 0.112, 0.08, 0.052, 0.025, 0, -0.027, -0.034, -0.08, 
    -0.068, -0.039, -0.15, -0.195,
  5.465, 1.791, 0.709, 0.14, 0.102, 0.096, 0.077, 0.066, 0.054, 0.016, -0.03, 
    -0.093, -0.146, -0.285, -0.236,
  4.884, 1.53, 0.73, 0.135, 0.108, 0.113, 0.099, 0.073, 0.031, -0.027, -0.08, 
    -0.158, -0.189, -0.296, -0.22,
  4.455, 1.372, 0.728, 0.111, 0.079, 0.076, 0.068, 0.065, 0.05, 0.029, -0.03, 
    -0.061, -0.136, -0.217, -0.174,
  2.216, 0.795, 0.423, 0.056, 0.038, 0.039, 0.046, 0.047, 0.039, 0.022, 
    0.013, 0.001, -0.026, -0.062, -0.018,
  0.73, 0.07, -0.013, -0.026, -0.016, -0.015, -0.014, -0.015, -0.008, -0.006, 
    -0.017, -0.025, -0.055, -0.101, -0.064,
  -0.905, -0.412, -0.438, -0.118, -0.066, -0.06, -0.059, -0.061, -0.068, 
    -0.068, -0.064, -0.061, -0.065, -0.066, 0,
  -0.031, -0.205, -0.311, -0.096, -0.05, -0.054, -0.058, -0.061, -0.063, 
    -0.067, -0.061, -0.049, -0.032, 0.002, 0.049,
  1.295, 0.4, 0.252, 0.031, -0.004, -0.01, -0.01, -0.016, -0.023, -0.033, 
    -0.036, -0.035, -0.02, 0.003, 0.031,
  2.601, 0.668, 0.557, 0.109, 0.035, 0.032, 0.031, 0.034, 0.04, 0.034, 0.028, 
    0.019, 0.005, 0.005, -0.035,
  3.944, 1.101, 1.026, 0.244, 0.098, 0.089, 0.089, 0.095, 0.095, 0.098, 
    0.094, 0.082, 0.054, 0.002, -0.016,
  3.465, 0.896, 0.729, 0.246, 0.132, 0.121, 0.122, 0.122, 0.127, 0.123, 
    0.117, 0.104, 0.082, 0.029, -0.008,
  3.44, 0.753, 0.576, 0.226, 0.143, 0.137, 0.134, 0.126, 0.117, 0.108, 0.091, 
    0.072, 0.058, 0.02, 0.052,
  3.056, 0.647, 0.447, 0.178, 0.115, 0.113, 0.121, 0.128, 0.125, 0.118, 0.1, 
    0.08, 0.076, 0.053, 0.112,
  1.859, 0.393, 0.228, 0.121, 0.095, 0.093, 0.09, 0.083, 0.081, 0.084, 0.097, 
    0.104, 0.109, 0.061, 0.023,
  1.266, 0.206, 0.103, 0.064, 0.05, 0.046, 0.043, 0.046, 0.044, 0.048, 0.051, 
    0.054, 0.059, 0.062, 0.128,
  0.735, 0.083, 0.022, 0.001, -0.004, -0.013, -0.01, -0.013, -0.018, -0.007, 
    0.001, -0.005, 0.01, 0.036, -0.008,
  -0.415, -0.23, -0.223, -0.125, -0.084, -0.091, -0.096, -0.092, -0.083, 
    -0.089, -0.066, -0.039, -0.02, -62.408, -187.284,
  -1.002, -0.361, -0.289, -0.136, -0.093, -0.084, -0.082, -499.527, -499.538, 
    -499.524, -499.51, -499.508, -499.503, -561.936, -561.938,
  0.226, -0.055, -249.707, -249.763, -499.518, -499.511, -499.509, -0.028, 
    -187.363, -62.521, -0.12, -499.552, -561.989, -749.25, -561.938,
  -0.499, -0.464, -250.086, -249.831, -0.057, -0.05, -0.053, -0.076, 
    -187.349, -62.472, -0.046, -0.05, -62.524, -249.898, -561.938,
  1.95, 0.489, 0.43, 0.064, 0.022, 0.01, 0.003, 0.005, 0.004, -0.009, -0.014, 
    -0.016, 0.01, 0.023, 0.014,
  2.447, 0.678, 0.577, 0.105, 0.064, 0.061, 0.055, 0.048, 0.041, 0.03, 0.018, 
    0.008, 0.005, -0.011, -0.032,
  3.193, 0.92, 0.783, 0.145, 0.083, 0.078, 0.077, 0.07, 0.07, 0.062, 0.049, 
    0.035, 0.003, -0.048, -0.016,
  3.74, 1.025, 0.839, 0.161, 0.1, 0.096, 0.094, 0.083, 0.081, 0.067, 0.06, 
    0.053, 0.036, 0.02, -0.049,
  3.484, 0.978, 0.801, 0.146, 0.085, 0.074, 0.068, 0.065, 0.068, 0.068, 0.06, 
    0.056, 0.057, 0.039, 0.016,
  2.539, 0.733, 0.557, 0.089, 0.055, 0.05, 0.052, 0.051, 0.045, 0.041, 0.037, 
    0.026, 0.015, -0.004, -0.007,
  1.805, 0.499, 0.367, 0.058, 0.026, 0.026, 0.026, 0.023, 0.021, 0.014, 
    0.006, -0.002, -0.018, -0.038, -0.036,
  1.466, 0.399, 0.278, 0.034, 0.019, 0.014, 0.016, 0.011, 0.009, 0.003, 
    -0.003, -0.01, -0.022, -0.029, -0.041,
  0.455, 0.168, 0.115, 0.013, -0.001, -0.001, -0.004, -0.009, -0.009, -0.007, 
    -0.009, -0.011, -0.022, -0.024, -0.034,
  0.029, -0.081, -0.115, -0.038, -0.031, -0.035, -0.033, -0.03, -0.034, 
    -0.028, -0.023, -0.038, -0.042, -0.063, -0.04,
  0.42, -0.064, -0.066, -0.024, -0.02, -0.024, -0.032, -0.04, -0.044, -0.062, 
    -0.07, -0.087, -0.094, -0.088, -0.056,
  2.042, 0.576, 0.276, 0.04, 0.026, 0.018, 0.003, -0.014, -0.018, -0.022, 
    -0.025, -0.031, -0.034, -0.066, -0.054,
  3.694, 1.079, 0.614, 0.136, 0.095, 0.094, 0.07, 0.056, 0.05, 0.029, 0.007, 
    -0.011, -0.062, -0.101, -0.103,
  5.848, 1.921, 1.074, 0.263, 0.181, 0.156, 0.118, 0.093, 0.072, 0.07, 0.012, 
    -0.059, -0.064, -0.114, -0.048,
  6.383, 1.736, 0.92, 0.202, 0.155, 0.15, 0.128, 0.103, 0.057, 0.022, 0.009, 
    -0.009, -0.05, -0.134, -0.145,
  5.657, 1.53, 0.677, 0.108, 0.084, 0.076, 0.074, 0.055, 0.034, -0.015, 
    -0.089, -0.142, -0.167, -0.227, -0.276,
  5.677, 1.494, 0.716, 0.153, 0.126, 0.116, 0.106, 0.088, 0.052, 0.009, 
    -0.031, -0.106, -0.139, -0.225, -0.297,
  7.267, 1.914, 0.849, 0.218, 0.204, 0.197, 0.193, 0.176, 0.17, 0.103, 0.045, 
    -0.073, -0.178, -0.294, -0.316,
  7.009, 2.027, 0.91, 0.217, 0.195, 0.208, 0.215, 0.205, 0.172, 0.128, 0.048, 
    -0.05, -0.168, -0.265, -0.355,
  5.409, 1.519, 0.742, 0.183, 0.164, 0.171, 0.174, 0.178, 0.171, 0.13, 0.066, 
    -0.011, -0.082, -0.153, -0.137,
  3.244, 1.013, 0.53, 0.111, 0.091, 0.089, 0.092, 0.092, 0.081, 0.061, 0.036, 
    0.008, -0.053, -0.151, -0.097,
  2.074, 0.601, 0.244, 0.019, 0.013, 0.013, 0.009, -0.002, -0.009, -0.02, 
    -0.033, -0.043, -0.038, -0.05, -0.036,
  0.632, 0.03, -0.118, -0.056, -0.042, -0.039, -0.038, -0.036, -0.037, 
    -0.041, -0.043, -0.039, -0.045, -0.072, -0.017,
  0.131, -0.014, -0.074, -0.053, -0.044, -0.045, -0.048, -0.055, -0.057, 
    -0.059, -0.059, -0.063, -0.064, -0.073, -0.004,
  0.185, 0.024, -0.067, -0.055, -0.04, -0.043, -0.047, -0.053, -0.054, 
    -0.053, -0.047, -0.032, -0.042, -0.037, -0.009,
  0.466, 0.137, 0.087, 0.007, -0.004, -0.007, -0.011, -0.012, -0.019, -0.025, 
    -0.021, -0.016, -0.012, -0.01, -0.007,
  0.88, 0.177, 0.131, 0.047, 0.029, 0.027, 0.029, 0.03, 0.029, 0.028, 0.02, 
    0.013, -0.006, -0.018, 0.024,
  1.56, 0.365, 0.24, 0.104, 0.077, 0.073, 0.072, 0.069, 0.068, 0.063, 0.053, 
    0.045, 0.019, -0.012, 0.003,
  2.092, 0.435, 0.234, 0.123, 0.099, 0.091, 0.086, 0.081, 0.075, 0.061, 
    0.046, 0.033, 0.021, 0.011, 0.007,
  1.81, 0.398, 0.201, 0.129, 0.11, 0.1, 0.095, 0.087, 0.079, 0.068, 0.058, 
    0.045, 0.035, 0.023, 0.053,
  1.39, 0.308, 0.135, 0.08, 0.07, 0.061, 0.05, 0.037, 0.029, 0.019, 0.015, 
    0.024, 0.03, 0.033, 0.06,
  0.637, 0.09, 0.026, 0.02, 0.017, 0.017, 0.008, 0.015, 0.016, 0.033, 0.024, 
    0.039, 0.01, 0.04, 0.035,
  0.239, -0.004, -0.044, -0.025, -0.021, -0.02, -0.022, -0.025, -0.025, 
    -0.029, -0.015, -0.003, 0.021, 0.046, 0.043,
  -0.589, -0.309, -0.117, -0.065, -0.05, -0.059, -0.07, -0.072, -0.066, 
    -0.052, -0.058, 0, -0.002, -374.629, -561.932,
  -374.872, -499.597, -499.54, -499.525, -499.519, -499.519, -0.015, -0.023, 
    -499.53, -499.53, -0.108, -0.041, -499.508, -749.25, -561.938,
  -374.221, -499.387, -499.297, -499.462, -499.488, -499.488, -499.499, 
    -499.511, -374.632, 0.022, -374.606, -499.462, -749.25, -749.25, -561.938,
  2.83, 0.837, 0.822, 0.134, 0.05, 0.043, 0.029, 0.049, 0.061, 0.064, 0.067, 
    0.018, -249.73, -749.227, -561.91,
  2.548, 0.662, 0.572, 0.08, 0.05, 0.048, 0.06, 0.074, 0.067, 0.064, 0.056, 
    0.063, 0.072, 0.065, -0.013,
  3.736, 1.061, 0.866, 0.125, 0.076, 0.068, 0.064, 0.057, 0.059, 0.055, 0.04, 
    0.031, 0.019, -0.001, -0.005,
  3.92, 1.031, 0.759, 0.141, 0.084, 0.079, 0.073, 0.068, 0.061, 0.051, 0.043, 
    0.032, 0.016, -0.008, -0.021,
  3.627, 1.048, 0.743, 0.125, 0.081, 0.068, 0.067, 0.061, 0.042, 0.027, 
    0.018, 0.008, -0.007, -0.026, -0.061,
  3.382, 0.838, 0.551, 0.095, 0.056, 0.046, 0.038, 0.03, 0.032, 0.033, 0.021, 
    0.01, -0.003, -0.023, -0.011,
  3.285, 0.905, 0.584, 0.105, 0.066, 0.056, 0.048, 0.033, 0.014, 0.002, 
    -0.009, -0.024, -0.034, -0.087, -0.096,
  2.896, 0.77, 0.414, 0.051, 0.028, 0.03, 0.023, 0.021, 0.011, -0.01, -0.03, 
    -0.056, -0.077, -0.085, -0.099,
  2.148, 0.597, 0.351, 0.055, 0.031, 0.019, 0.015, 0.008, 0.003, -0.002, 
    -0.027, -0.044, -0.066, -0.059, -0.068,
  1.42, 0.409, 0.16, 0.021, 0.009, 0.006, -0.002, -0.012, -0.018, -0.034, 
    -0.046, -0.067, -0.094, -0.116, -0.074,
  1.508, 0.246, 0.086, -0.003, 0, 0, -0.005, -0.012, -0.018, -0.022, -0.047, 
    -0.051, -0.071, -0.052, -0.058,
  0.834, 0.225, 0.081, 0, -0.01, -0.017, -0.019, -0.024, -0.034, -0.047, 
    -0.05, -0.079, -0.086, -0.12, -0.037,
  2.327, 0.481, 0.16, 0.027, 0.021, 0.017, 0.008, -0.001, -0.01, -0.023, 
    -0.035, -0.043, -0.035, -0.058, 0.014,
  2.829, 0.726, 0.302, 0.087, 0.079, 0.077, 0.076, 0.066, 0.065, 0.047, 0.03, 
    -0.009, -0.054, -0.156, -0.012,
  2.548, 0.971, 0.401, 0.123, 0.11, 0.106, 0.087, 0.075, 0.068, 0.059, 0.032, 
    0, -0.032, -0.122, -0.007,
  1.611, 0.726, 0.399, 0.113, 0.097, 0.086, 0.082, 0.081, 0.055, 0.024, 0.02, 
    -0.001, -0.023, -0.038, -0.007,
  1.253, 0.579, 0.171, 0.015, 0.006, 0.005, 0.004, 0.004, -0.012, -0.014, 
    -0.02, -0.006, 0.003, 0.017, -0,
  0.603, 0.367, 0.113, 0.014, 0.012, 0.005, -0, -0.013, -0.005, 0.007, 0.029, 
    0.033, 0.008, -0.022, 0.03,
  0.504, 0.407, 0.193, 0.061, 0.053, 0.061, 0.072, 0.07, 0.069, 0.043, 0.027, 
    0.011, 0.002, -0.02, -0.019,
  0.821, 0.466, 0.268, 0.098, 0.096, 0.097, 0.095, 0.092, 0.083, 0.074, 
    0.061, 0.046, 0.031, -0.013, -0.019,
  0.662, 0.371, 0.269, 0.112, 0.1, 0.097, 0.099, 0.105, 0.114, 0.108, 0.097, 
    0.071, 0.048, 0.028, 0.008,
  0.637, 0.215, 0.14, 0.058, 0.059, 0.06, 0.059, 0.062, 0.055, 0.055, 0.053, 
    0.042, 0.038, 0.012, 0.039,
  0.445, 0.158, 0.079, 0.032, 0.025, 0.027, 0.029, 0.027, 0.03, 0.026, 0.021, 
    0.02, 0.035, 0.021, 0.041,
  -0.017, -0.02, -0.033, -0.018, -0.014, -0.014, -0.012, -0.011, -0.01, 
    -0.009, -0.008, -0.004, -0, 0.001, 0.027,
  -0.132, -0.028, -0.033, -0.026, -0.024, -0.027, -0.032, -0.034, -0.032, 
    -0.028, -0.024, -0.013, -0.008, 0.011, 0.008,
  -0.166, -0.052, -0.048, -0.037, -0.036, -0.039, -0.038, -0.039, -0.04, 
    -0.04, -0.034, -0.025, -0.016, 0.01, 0.02,
  0.276, 0.045, 0.019, -0.003, -0.015, -0.02, -0.028, -0.035, -0.034, -0.029, 
    -0.025, -0.016, -0.015, 0.004, 0.018,
  0.503, 0.112, 0.059, 0.029, 0.02, 0.012, 0.008, 0.003, -0.001, -0.002, 
    -0.002, -0.002, -0.012, -0.008, 0.041,
  1.099, 0.229, 0.104, 0.064, 0.054, 0.045, 0.037, 0.032, 0.03, 0.028, 0.023, 
    0.023, -0.006, -0.015, 0.043,
  1.57, 0.338, 0.154, 0.093, 0.07, 0.06, 0.048, 0.041, 0.032, 0.023, 0.019, 
    0.019, 0.014, 0.015, 0.041,
  1.26, 0.292, 0.125, 0.075, 0.058, 0.048, 0.037, 0.03, 0.023, 0.006, -0.001, 
    0, -0.015, -0.011, 0.01,
  1.103, 0.277, 0.111, 0.053, 0.034, 0.016, 0.008, -0.005, -0.014, -0.019, 
    -0.027, -0.029, -0.044, -0.025, -0.03,
  0.758, 0.216, 0.061, 0.011, -0.007, -0.029, -0.043, -0.046, -0.055, -0.037, 
    -0.028, -0.005, 0.018, 0.026, 0.012,
  0.221, 0.072, -0.039, -0.056, -0.054, -0.053, -0.061, -0.07, -0.068, 
    -0.059, -0.05, -0.028, -0.014, 0.054, 0.007,
  -0.191, -0.077, -0.105, -0.092, -0.083, -0.103, -0.107, -0.102, -0.104, 
    -0.093, -0.083, -0.088, -0.012, -62.382, -187.297,
  -1.299, -0.295, -0.107, -124.911, -499.516, -499.526, -499.532, -499.544, 
    -499.549, -125.021, -499.54, -499.533, -499.484, -561.916, -561.938,
  3.908, 1.04, 0.988, -374.532, -499.48, -499.481, -499.478, -749.25, 
    -499.52, -499.555, -499.558, -499.519, 0.171, -561.879, -561.938,
  4.011, 1.014, 0.862, 0.118, 0.024, -0.026, -0.03, -249.809, -0.074, -0.072, 
    -0.076, -0.104, -0.037, -62.491, -187.459,
  2.96, 0.728, 0.488, 0.056, 0.025, 0.035, 0.013, 0.015, 0.037, -0.025, 
    -0.041, -0.064, -0.028, -0.109, -0.053,
  2.824, 0.727, 0.511, 0.109, 0.073, 0.063, 0.065, 0.059, 0.052, 0.037, 
    -0.009, 0.022, -0.022, -0.109, -0.061,
  3.486, 0.933, 0.666, 0.116, 0.075, 0.071, 0.073, 0.081, 0.072, 0.06, 0.027, 
    0.017, -0.03, -0.022, -0.013,
  3.25, 0.799, 0.493, 0.1, 0.07, 0.061, 0.058, 0.046, 0.023, 0, -0.021, 
    -0.043, -0.087, -0.137, -0.089,
  3.288, 0.69, 0.377, 0.078, 0.058, 0.054, 0.05, 0.037, 0.03, 0.017, -0.007, 
    -0.026, -0.052, -0.117, -0.098,
  2.877, 0.637, 0.279, 0.067, 0.049, 0.046, 0.049, 0.052, 0.049, 0.034, 0.01, 
    -0.023, -0.053, -0.066, -0.073,
  1.026, 0.238, 0.138, 0.032, 0.024, 0.021, 0.016, -0.001, -0.013, -0.028, 
    -0.042, -0.049, -0.082, -0.106, -0.094,
  1.416, 0.244, 0.05, -0.003, -0.006, -0.004, -0.004, -0.006, -0.015, -0.03, 
    -0.05, -0.078, -0.112, -0.094, -0.111,
  0.844, 0.102, 0.011, -0.006, -0.008, -0.012, -0.013, -0.02, -0.026, -0.037, 
    -0.049, -0.052, -0.063, -0.044, -0.08,
  1, 0.194, 0.063, 0.013, 0.004, 0.003, 0.001, -0.002, -0.013, -0.016, 
    -0.021, -0.024, -0.017, -0.068, -0.014,
  0.397, 0.107, 0.052, 0.021, 0.019, 0.016, 0.012, 0.01, 0.012, -0, -0.014, 
    -0.033, -0.027, -0.065, -0.016,
  0.997, 0.155, 0.056, 0.029, 0.034, 0.043, 0.05, 0.046, 0.035, 0.031, 0.016, 
    0.003, -0.01, -0.038, -0.054,
  0.738, 0.191, 0.121, 0.066, 0.064, 0.066, 0.072, 0.08, 0.079, 0.074, 0.059, 
    0.019, 0.005, -0.065, 0.016,
  0.517, 0.21, 0.14, 0.087, 0.088, 0.092, 0.098, 0.103, 0.116, 0.125, 0.116, 
    0.108, 0.084, 0.002, 0.067,
  0.018, 0.011, 0.015, 0.044, 0.053, 0.054, 0.058, 0.071, 0.073, 0.073, 
    0.073, 0.055, 0.062, 0.022, 0.042,
  -0.092, -0.057, -0.041, -0.026, -0.018, -0.012, -0.005, 0.001, 0.009, 
    0.017, 0.025, 0.045, 0.058, 0.086, 0.031,
  -0.144, -0.12, -0.118, -0.052, -0.044, -0.038, -0.033, -0.032, -0.021, 
    -0.009, 0, 0.011, 0.041, 0.085, 0.06,
  -0.212, -0.152, -0.122, -0.041, -0.027, -0.019, -0.018, -0.009, 0.002, 
    0.004, 0.016, 0.036, 0.063, 0.067, 0.122,
  -0.102, -0.048, -0.022, 0.002, 0.005, 0.004, 0.011, 0.017, 0.026, 0.034, 
    0.037, 0.051, 0.072, 0.086, 0.11,
  0.017, 0.013, 0.027, 0.02, 0.023, 0.022, 0.026, 0.023, 0.022, 0.031, 0.045, 
    0.062, 0.071, 0.075, 0.095,
  0.06, 0.016, 0.018, 0.011, 0.015, 0.017, 0.016, 0.027, 0.037, 0.047, 0.05, 
    0.068, 0.066, 0.047, 0.145,
  0.154, 0.034, 0.028, 0.03, 0.027, 0.032, 0.036, 0.039, 0.046, 0.053, 0.058, 
    0.06, 0.058, 0.065, 0.098,
  0.159, 0.038, 0.036, 0.024, 0.03, 0.026, 0.028, 0.033, 0.036, 0.038, 0.048, 
    0.065, 0.066, 0.082, 0.069,
  0.162, 0.005, 0.005, 0.002, 0, 0.003, 0.007, 0.01, 0.015, 0.025, 0.032, 
    0.046, 0.055, 0.071, 0.071,
  0.127, -0, -0.009, -0.015, -0.018, -0.018, -0.016, -0.011, -0.002, 0.005, 
    0.019, 0.026, 0.022, 0.04, 0.05,
  0.293, 0.064, 0.021, 0.009, 0.006, 0.003, 0.001, -0.001, -0.002, 0.002, 
    0.002, 0.019, 0.015, 0.024, 0.034,
  0.499, 0.09, 0.047, 0.032, 0.025, 0.019, 0.017, 0.017, 0.019, 0.015, 0.019, 
    0.02, 0.019, 0.03, 0.027,
  1.013, 0.206, 0.083, 0.057, 0.051, 0.051, 0.053, 0.056, 0.05, 0.051, 0.049, 
    0.047, 0.034, 0.028, 0.026,
  1.358, 0.326, 0.117, 0.089, 0.078, 0.079, 0.074, 0.07, 0.073, 0.067, 0.066, 
    0.062, 0.05, 0.05, 0.035,
  1.201, 0.305, 0.113, 0.079, 0.065, 0.061, 0.061, 0.061, 0.056, 0.055, 
    0.052, 0.045, 0.031, 0.016, 0.034,
  0.711, 0.191, 0.075, 0.049, 0.033, 0.025, 0.019, 0.016, 0.014, 0.021, 
    0.021, 0.027, 0.041, 0.048, 0.043,
  0.4, 0.118, 0.029, 0.007, -0.009, -0.018, -0.022, -0.019, -0.014, -0.007, 
    0.02, 0.028, 0.025, 0.041, 0.016,
  -0.196, -0.047, -0.032, -0.035, -0.041, -0.051, -0.053, -0.056, -0.047, 
    -0.022, -0.012, -0.008, 0.003, 0.021, 0.012,
  -0.709, -0.143, -0.055, -0.09, -0.085, -0.083, -0.087, -0.081, -0.088, 
    -62.503, -0.085, -0.032, 0.033, -187.235, -187.306,
  -374.969, -499.597, -124.939, -0.033, -0.025, -0.03, -499.517, -499.512, 
    -374.653, -62.505, -0.059, -499.492, -499.474, -686.794, -561.938,
  -378.09, -499.9, -499.807, -499.559, -499.534, -499.534, -499.553, 
    -686.826, -561.943, -499.503, -499.503, 0.088, -499.478, -749.25, -561.938,
  0.319, 0.713, 0.573, 0.077, 0.019, 0.017, -0.02, -187.381, -62.535, -0.126, 
    -499.543, -499.5, 0.19, -374.556, -561.932,
  3.104, 0.579, 0.428, 0.07, 0.105, 0.134, 0.077, 0.05, 0.033, 0.006, -0.052, 
    -0.081, -0.082, -0.077, -0.062,
  1.695, 0.513, 0.373, 0.096, 0.079, 0.074, 0.078, 0.084, 0.07, 0.06, 0.045, 
    0.013, 0.009, -0.107, -0.018,
  3.862, 0.954, 0.515, 0.124, 0.102, 0.103, 0.104, 0.109, 0.108, 0.039, 
    0.004, 0.013, -0.089, -0.19, -0.108,
  2.362, 0.523, 0.223, 0.072, 0.057, 0.063, 0.065, 0.062, 0.053, 0.058, 
    0.028, 0.002, -0.017, -0.054, -0.027,
  2.427, 0.527, 0.172, 0.062, 0.056, 0.058, 0.062, 0.06, 0.055, 0.041, 0.029, 
    0.013, -0.014, -0.081, -0.017,
  2.077, 0.409, 0.14, 0.057, 0.05, 0.05, 0.046, 0.047, 0.048, 0.046, 0.032, 
    0.021, 0.013, -0.013, -0.007,
  1.797, 0.372, 0.11, 0.037, 0.034, 0.033, 0.032, 0.027, 0.017, 0.012, 0.006, 
    -0.007, -0.017, -0.012, -0.002,
  1.072, 0.167, 0.042, 0.015, 0.013, 0.012, 0.014, 0.012, 0.012, 0.009, 
    -0.004, -0.001, -0.002, -0.01, -0.027,
  1.502, 0.282, 0.079, 0.043, 0.04, 0.037, 0.034, 0.028, 0.018, 0.009, 0.006, 
    -0.011, -0.015, -0.016, -0.001,
  1.307, 0.221, 0.072, 0.042, 0.04, 0.043, 0.048, 0.053, 0.056, 0.057, 0.05, 
    0.03, 0.03, -0.076, -0.007,
  1.524, 0.251, 0.092, 0.053, 0.052, 0.053, 0.059, 0.062, 0.065, 0.061, 
    0.061, 0.054, 0.07, -0.002, 0.07,
  1.166, 0.21, 0.092, 0.069, 0.069, 0.076, 0.082, 0.087, 0.093, 0.098, 0.093, 
    0.071, 0.08, -0.001, 0.047,
  0.423, 0.123, 0.085, 0.067, 0.07, 0.071, 0.084, 0.098, 0.102, 0.106, 0.102, 
    0.093, 0.1, 0.033, 0.064,
  -0.096, -0.026, 0.03, 0.062, 0.079, 0.094, 0.106, 0.118, 0.13, 0.141, 
    0.134, 0.139, 0.138, 0.083, 0.125,
  -0.302, -0.169, -0.111, -0.021, 0.016, 0.035, 0.056, 0.074, 0.096, 0.118, 
    0.125, 0.144, 0.166, 0.105, 0.014,
  -0.264, -0.162, -0.137, -0.074, -0.047, -0.036, -0.027, -0.014, 0.003, 
    0.011, 0.037, 0.062, 0.124, 0.119, 0.077,
  -0.241, -0.18, -0.166, -0.099, -0.076, -0.07, -0.07, -0.056, -0.048, -0.03, 
    -0.016, 0.03, 0.096, 0.121, 0.188,
  -0.259, -0.209, -0.197, -0.098, -0.069, -0.06, -0.051, -0.047, -0.034, 
    -0.021, -0.004, 0.02, 0.069, 0.104, 0.179,
  -0.243, -0.148, -0.119, -0.054, -0.028, -0.019, -0.011, -0.008, -0.004, 
    0.006, 0.016, 0.042, 0.066, 0.074, 0.167,
  -0.126, -0.064, -0.053, -0.018, -0.006, -0.006, -0.01, -0.007, -0.012, 
    -0.005, 0.01, 0.02, 0.032, 0.034, 0.117,
  -0.048, -0.024, 0.011, 0.019, 0.021, 0.009, 0.008, 0.014, 0.019, 0.021, 
    0.027, 0.043, 0.039, 0.033, 0.07,
  0.066, 0.022, 0.029, 0.035, 0.042, 0.049, 0.051, 0.049, 0.053, 0.06, 0.054, 
    0.042, 0.037, 0.029, 0.049,
  0.371, 0.052, 0.03, 0.032, 0.031, 0.033, 0.039, 0.044, 0.047, 0.043, 0.045, 
    0.043, 0.039, 0.024, 0.023,
  0.613, 0.095, 0.039, 0.023, 0.023, 0.023, 0.022, 0.02, 0.019, 0.02, 0.02, 
    0.012, 0.022, 0.003, 0.046,
  0.584, 0.09, 0.028, 0.013, 0.008, 0.005, 0.006, 0.004, 0.002, 0.001, 
    -0.001, 0.005, 0.001, 0.011, 0.017,
  0.684, 0.119, 0.033, 0.02, 0.016, 0.011, 0.011, 0.011, 0.009, 0.009, 0.005, 
    -0.004, -0.01, -0.021, 0.01,
  0.741, 0.165, 0.053, 0.039, 0.038, 0.04, 0.044, 0.043, 0.037, 0.028, 0.018, 
    0.009, -0.009, -0.034, 0.001,
  0.84, 0.239, 0.087, 0.068, 0.07, 0.07, 0.069, 0.068, 0.072, 0.074, 0.063, 
    0.058, 0.047, -0.007, -0.007,
  0.934, 0.238, 0.079, 0.066, 0.062, 0.068, 0.073, 0.078, 0.076, 0.072, 
    0.068, 0.061, 0.046, 0.051, 0.007,
  0.711, 0.189, 0.07, 0.058, 0.05, 0.052, 0.057, 0.063, 0.067, 0.067, 0.059, 
    0.054, 0.036, 0.02, 0.009,
  0.551, 0.142, 0.051, 0.046, 0.042, 0.042, 0.042, 0.041, 0.043, 0.05, 0.057, 
    0.039, 0.019, 0.005, 0.006,
  0.111, 0.038, 0.015, 0.018, 0.022, 0.028, 0.039, 0.051, 0.059, 0.059, 
    0.051, 0.048, 0.028, -0.013, 0.025,
  -0.092, -0.056, -0.019, -0.009, -0.016, -0.021, -0.016, -0.013, -0.008, 
    -0.006, 0.015, 0.036, 0.065, 0.068, 0.08,
  -0.679, -0.192, -0.063, -0.045, -0.047, -0.053, -0.052, -0.052, -0.043, 
    -0.025, 0.014, 0.028, 0.064, -249.647, -187.267,
  -0.45, -0.052, 0.217, -0.045, -0.039, -0.044, -499.52, -0.027, 0.035, 
    0.015, 0.01, -499.482, -499.461, -749.25, -561.938,
  -249.981, 0.268, 0.25, -0.023, -249.724, -249.725, -249.721, -374.601, 
    -499.476, -499.467, -499.466, -499.48, -499.51, -499.516, -561.938,
  2.784, 0.28, 0.33, -0.018, -249.755, -249.731, -249.732, 0.04, 0.089, 0.08, 
    0.031, 0.089, 0.083, 0.035, -187.276,
  2.233, 0.385, 0.402, 0.096, 0.063, 0.074, 0.087, 0.098, 0.12, 0.13, 0.132, 
    0.11, 0.136, 0.131, 0.075,
  3.041, 0.526, 0.461, 0.122, 0.093, 0.104, 0.128, 0.145, 0.144, 0.134, 0.11, 
    0.12, 0.107, 0.059, 0.062,
  2.061, 0.471, 0.205, 0.091, 0.094, 0.107, 0.108, 0.113, 0.121, 0.122, 
    0.119, 0.109, 0.105, 0.09, 0.063,
  1.56, 0.385, 0.123, 0.059, 0.054, 0.055, 0.057, 0.052, 0.049, 0.058, 0.055, 
    0.061, 0.057, 0.079, 0.04,
  1.546, 0.342, 0.092, 0.049, 0.043, 0.046, 0.051, 0.051, 0.063, 0.061, 
    0.059, 0.046, 0.037, 0.015, 0.041,
  1.404, 0.253, 0.069, 0.046, 0.04, 0.046, 0.046, 0.053, 0.048, 0.043, 0.044, 
    0.059, 0.068, 0.102, 0.051,
  1.193, 0.237, 0.069, 0.041, 0.041, 0.046, 0.049, 0.05, 0.056, 0.055, 0.046, 
    0.046, 0.056, 0.08, 0.047,
  1.441, 0.277, 0.084, 0.054, 0.054, 0.057, 0.065, 0.07, 0.071, 0.076, 0.076, 
    0.079, 0.069, 0.056, 0.018,
  2.028, 0.402, 0.115, 0.07, 0.064, 0.069, 0.076, 0.08, 0.094, 0.092, 0.092, 
    0.08, 0.085, 0.059, 0.039,
  1.731, 0.32, 0.109, 0.068, 0.065, 0.065, 0.069, 0.068, 0.061, 0.055, 0.055, 
    0.05, 0.045, 0.018, 0.007,
  1.582, 0.301, 0.103, 0.07, 0.065, 0.063, 0.067, 0.068, 0.074, 0.075, 0.071, 
    0.044, 0.039, -0.013, -0.02,
  0.797, 0.193, 0.077, 0.06, 0.057, 0.057, 0.063, 0.075, 0.079, 0.08, 0.076, 
    0.065, 0.074, -0.005, -0.059,
  -0.001, 0.012, 0.033, 0.049, 0.062, 0.069, 0.071, 0.063, 0.062, 0.064, 
    0.063, 0.044, 0.047, 0.008, -0.128,
  -0.703, -0.265, -0.114, -0.018, 0.019, 0.031, 0.046, 0.061, 0.075, 0.083, 
    0.073, 0.067, 0.057, 0.032, -0.075,
  -0.428, -0.251, -0.184, -0.093, -0.037, -0.01, 0.002, 0.018, 0.017, 0.03, 
    0.052, 0.062, 0.086, 0.093, -0.043,
  -0.264, -0.156, -0.138, -0.106, -0.08, -0.068, -0.056, -0.046, -0.033, 
    -0.024, -0.018, 0.013, 0.078, 0.1, 0.028,
  -0.168, -0.11, -0.069, -0.048, -0.045, -0.047, -0.05, -0.053, -0.051, 
    -0.04, -0.022, -0.002, 0.036, 0.097, 0.071,
  -0.119, -0.062, -0.06, -0.056, -0.051, -0.048, -0.049, -0.053, -0.046, 
    -0.039, -0.022, -0.002, 0.037, 0.123, 0.106,
  -0.12, -0.071, -0.062, -0.058, -0.045, -0.04, -0.041, -0.032, -0.024, 
    -0.015, 0, 0.015, 0.035, 0.095, 0.084,
  -0.075, -0.052, -0.05, -0.025, -0.01, -0.002, 0.008, 0.01, 0.036, 0.049, 
    0.06, 0.075, 0.079, 0.093, 0.056,
  0.041, 0.004, 0.036, 0.041, 0.055, 0.053, 0.054, 0.064, 0.067, 0.079, 
    0.086, 0.086, 0.084, 0.064, 0.059,
  0.398, 0.093, 0.064, 0.059, 0.068, 0.077, 0.086, 0.092, 0.089, 0.082, 
    0.081, 0.083, 0.075, 0.047, 0.016,
  0.792, 0.166, 0.089, 0.078, 0.082, 0.087, 0.09, 0.094, 0.099, 0.094, 0.091, 
    0.082, 0.072, 0.036, 0.039,
  1.03, 0.191, 0.085, 0.057, 0.052, 0.05, 0.049, 0.043, 0.043, 0.046, 0.041, 
    0.038, 0.026, 0.005, 0.045,
  0.908, 0.195, 0.054, 0.041, 0.035, 0.034, 0.032, 0.028, 0.026, 0.015, 
    0.008, -0, 0.007, 0.011, 0.023,
  0.958, 0.209, 0.058, 0.036, 0.032, 0.03, 0.031, 0.033, 0.026, 0.022, 0.018, 
    0.013, 0.01, 0.025, 0.001,
  0.843, 0.208, 0.057, 0.041, 0.038, 0.039, 0.038, 0.037, 0.039, 0.034, 
    0.031, 0.014, 0.015, 0.012, 0.013,
  0.971, 0.277, 0.082, 0.061, 0.055, 0.052, 0.052, 0.052, 0.048, 0.046, 
    0.035, 0.034, 0.028, 0.011, -0.002,
  0.901, 0.265, 0.079, 0.063, 0.057, 0.055, 0.052, 0.05, 0.049, 0.047, 0.052, 
    0.048, 0.037, 0.022, 0.005,
  0.645, 0.21, 0.058, 0.042, 0.032, 0.027, 0.028, 0.025, 0.025, 0.024, 0.017, 
    0.016, 0.017, 0.009, 0.004,
  0.376, 0.116, 0.038, 0.031, 0.025, 0.024, 0.026, 0.028, 0.031, 0.033, 
    0.032, 0.024, 0.015, 0.012, 0.009,
  0.02, 0.012, 0.013, 0.015, 0.011, 0.016, 0.022, 0.025, 0.025, 0.028, 0.03, 
    0.032, 0.021, -0.013, 0.015,
  -0.452, -0.118, -0.03, -0.024, -0.012, -0.015, -0.014, -0.002, 0.007, 
    0.005, 0.003, 0.002, 0.022, 0.037, 0.035,
  -0.69, -0.222, -0.069, -0.052, -0.051, -0.052, -0.054, -0.058, -0.064, 
    -0.058, -0.059, -0.047, -0.013, 0.017, -187.239,
  -0.636, -0.255, -0.044, -0.035, -0.049, -0.054, -0.057, -0.085, -0.071, 
    -0.083, -124.95, -499.527, -499.509, -499.496, -561.938,
  -374.674, -499.469, -499.491, -499.484, -0.004, -0.006, -0.013, -0.019, 
    -124.904, -499.513, -499.526, -499.53, -749.25, -749.25, -561.938,
  1.763, 0.178, 0.103, 0.018, 0.017, 0.042, 0.06, 0.073, 0.09, 0.043, 0.028, 
    0.005, -249.759, -249.744, -187.26,
  2.789, 0.54, 0.277, 0.069, 0.053, 0.048, 0.036, 0.028, 0.043, 0.047, 0.05, 
    0.072, 0.057, 0.006, 0.055,
  1.233, 0.274, 0.106, 0.04, 0.033, 0.036, 0.046, 0.046, 0.034, 0.008, 
    -0.002, -0.008, 0.025, 0.043, 0.031,
  1.408, 0.339, 0.11, 0.04, 0.039, 0.051, 0.059, 0.06, 0.062, 0.064, 0.063, 
    0.049, 0.033, 0.037, 0.022,
  1.508, 0.295, 0.094, 0.048, 0.043, 0.042, 0.047, 0.049, 0.055, 0.047, 
    0.041, 0.04, 0.036, 0.021, 0.02,
  0.678, 0.138, 0.049, 0.031, 0.03, 0.042, 0.041, 0.044, 0.039, 0.036, 0.035, 
    0.04, 0.041, 0.052, 0.027,
  1.149, 0.251, 0.062, 0.034, 0.032, 0.03, 0.032, 0.033, 0.036, 0.047, 0.046, 
    0.046, 0.04, 0.04, 0.014,
  0.897, 0.194, 0.054, 0.035, 0.035, 0.038, 0.042, 0.038, 0.035, 0.021, 
    0.017, 0.017, 0.022, 0.024, 0.016,
  1.168, 0.186, 0.058, 0.042, 0.038, 0.04, 0.042, 0.043, 0.035, 0.032, 0.023, 
    0.01, -0.009, -0.028, -0.02,
  1.654, 0.299, 0.102, 0.064, 0.058, 0.053, 0.055, 0.054, 0.055, 0.049, 
    0.036, 0.018, -0.018, -0.06, -0.045,
  1.83, 0.334, 0.128, 0.093, 0.08, 0.081, 0.08, 0.079, 0.07, 0.066, 0.066, 
    0.052, 0.05, 0.002, -0.049,
  1.2, 0.274, 0.116, 0.078, 0.072, 0.074, 0.075, 0.073, 0.067, 0.055, 0.048, 
    0.029, 0.014, -0.007, -0.035,
  0.436, 0.122, 0.056, 0.041, 0.042, 0.047, 0.063, 0.063, 0.059, 0.058, 
    0.038, 0.01, -0.027, -0.059, -0.061,
  -0.839, -0.179, -0.043, 0.012, 0.033, 0.043, 0.037, 0.049, 0.046, 0.044, 
    0.037, 0.033, -0.006, -0.062, -0.1,
  -0.568, -0.232, -0.133, -0.057, -0.019, 0.005, 0.01, 0.005, 0.001, -0, 
    -0.005, -0.008, -0.01, 0.003, -0.071,
  -0.291, -0.169, -0.134, -0.087, -0.054, -0.039, -0.029, -0.015, -0.003, 
    -0.01, -0.002, 0.013, 0.008, 0, -0.034,
  -0.174, -0.093, -0.081, -0.082, -0.068, -0.058, -0.053, -0.047, -0.039, 
    -0.028, -0.017, -0.005, 0.012, 0.04, -0.01,
  -0.057, 0.002, 0.015, -0.019, -0.034, -0.047, -0.049, -0.052, -0.049, 
    -0.035, -0.017, 0.003, 0.038, 0.102, 0.028,
  0.004, 0.013, 0.019, 0.015, -0.025, -0.033, -0.033, -0.029, -0.026, -0.022, 
    -0.01, 0.011, 0.044, 0.085, 0.082,
  -0.081, -0.044, -0.071, -0.091, -0.069, -0.053, -0.05, -0.051, -0.045, 
    -0.024, -0.012, 0.007, 0.045, 0.12, 0.081,
  -0.166, -0.137, -0.128, -0.096, -0.036, -0.014, -0.003, 0.012, 0.014, 
    0.019, 0.027, 0.045, 0.061, 0.098, 0.109,
  -0.14, -0.077, -0.054, -0.016, 0.024, 0.044, 0.055, 0.064, 0.081, 0.088, 
    0.092, 0.084, 0.076, 0.083, 0.08,
  0.243, 0.076, 0.065, 0.052, 0.071, 0.078, 0.091, 0.095, 0.1, 0.105, 0.112, 
    0.102, 0.102, 0.108, 0.098,
  0.605, 0.149, 0.109, 0.103, 0.117, 0.126, 0.128, 0.131, 0.131, 0.137, 
    0.131, 0.126, 0.113, 0.091, 0.068,
  1.645, 0.396, 0.16, 0.12, 0.113, 0.113, 0.126, 0.136, 0.139, 0.127, 0.115, 
    0.099, 0.075, 0.042, 0.046,
  1.951, 0.452, 0.138, 0.096, 0.089, 0.089, 0.087, 0.085, 0.08, 0.079, 0.068, 
    0.049, 0.049, 0.044, 0.032,
  1.458, 0.363, 0.102, 0.069, 0.06, 0.055, 0.05, 0.049, 0.044, 0.041, 0.042, 
    0.038, 0.039, 0.044, 0.024,
  1.112, 0.278, 0.074, 0.048, 0.044, 0.043, 0.044, 0.043, 0.038, 0.034, 
    0.027, 0.025, 0.024, 0.028, 0.023,
  0.995, 0.28, 0.077, 0.057, 0.05, 0.046, 0.046, 0.046, 0.048, 0.045, 0.042, 
    0.033, 0.027, 0.015, 0.019,
  0.938, 0.264, 0.076, 0.062, 0.056, 0.055, 0.051, 0.049, 0.045, 0.044, 
    0.043, 0.036, 0.028, 0.017, 0.011,
  0.698, 0.203, 0.061, 0.048, 0.041, 0.038, 0.042, 0.042, 0.042, 0.042, 0.04, 
    0.039, 0.034, 0.041, 0.033,
  0.383, 0.108, 0.039, 0.031, 0.024, 0.021, 0.02, 0.018, 0.019, 0.025, 0.026, 
    0.033, 0.027, 0.028, 0.008,
  -0.004, -0.002, 0.007, 0.011, 0.006, 0.008, 0.009, 0.017, 0.02, 0.025, 
    0.036, 0.033, 0.03, 0.021, 0.027,
  -0.239, -0.054, -0.017, -0.011, -0.014, -0.013, -0.01, -0.009, -0.004, 
    0.003, -0.001, 0.006, 0.01, 0.038, 0.025,
  -0.555, -0.173, -0.05, -0.034, -0.026, -0.027, -0.021, -0.012, -0.018, 
    -0.02, 0.002, 0.016, 0.036, 0.021, -0.011,
  -0.452, -0.181, -0.049, -0.037, -0.032, -0.03, -0.028, -0.02, 0.137, 0.034, 
    -0.011, -0.025, -374.561, -499.512, -374.638,
  -561.938, -749.25, -749.25, -749.25, -561.965, -499.538, -499.539, 
    -499.538, -499.535, -499.535, -499.522, -499.528, -499.524, -749.25, 
    -561.938,
  -187.079, -249.686, -249.825, -249.783, -62.455, 0.009, 0.01, -0.023, 
    -0.047, -0.096, -0.165, -0.175, -0.119, -249.828, -187.39,
  0.627, 0.137, 0.079, 0.035, 0.036, 0.045, 0.059, 0.066, 0.082, 0.069, 
    0.054, 0.054, 0.033, 0.027, 0.057,
  0.95, 0.245, 0.109, 0.035, 0.034, 0.043, 0.048, 0.055, 0.059, 0.053, 0.045, 
    0.036, 0.028, 0.005, 0.02,
  0.815, 0.193, 0.071, 0.034, 0.028, 0.031, 0.032, 0.026, 0.038, 0.036, 
    0.046, 0.032, 0.017, 0.015, 0.014,
  0.294, 0.075, 0.018, 0.013, 0.016, 0.018, 0.022, 0.023, 0.009, 0.001, 
    -0.013, -0.005, 0.008, 0.015, 0.021,
  0.611, 0.137, 0.04, 0.025, 0.024, 0.024, 0.026, 0.03, 0.032, 0.03, 0.026, 
    0.024, 0.011, 0.007, 0.013,
  0.485, 0.091, 0.027, 0.02, 0.019, 0.022, 0.027, 0.023, 0.016, 0.017, 0.016, 
    0.018, 0.005, -0.011, 0.013,
  0.78, 0.138, 0.037, 0.029, 0.033, 0.031, 0.028, 0.027, 0.024, 0.011, 0.005, 
    -0, 0.007, -0.004, -0.008,
  1.018, 0.185, 0.063, 0.039, 0.032, 0.044, 0.049, 0.047, 0.042, 0.033, 
    0.027, 0.028, 0.022, 0.014, 0.011,
  1.697, 0.328, 0.101, 0.066, 0.06, 0.045, 0.046, 0.054, 0.049, 0.037, 0.021, 
    0.001, -0.008, -0.034, 0.007,
  1.785, 0.373, 0.144, 0.091, 0.093, 0.095, 0.092, 0.079, 0.08, 0.072, 0.06, 
    0.032, -0.002, -0.056, -0.028,
  1.377, 0.38, 0.15, 0.098, 0.085, 0.083, 0.095, 0.097, 0.085, 0.082, 0.067, 
    0.059, 0.041, 0.004, -0.01,
  0, -0.041, 0.016, 0.06, 0.064, 0.074, 0.072, 0.072, 0.074, 0.063, 0.071, 
    0.058, 0.024, -0.02, 0.002,
  -1.055, -0.303, -0.14, -0.047, -0.007, 0.021, 0.037, 0.046, 0.05, 0.048, 
    0.027, 0.026, 0.03, -0.012, 0.044,
  -0.995, -0.461, -0.288, -0.15, -0.074, -0.038, -0.022, -0.009, 0.007, 
    0.011, 0.022, 0.013, 0.013, 0.03, -0.003,
  -0.416, -0.263, -0.222, -0.144, -0.094, -0.061, -0.045, -0.037, -0.034, 
    -0.028, -0.026, -0.014, 0.006, 0.018, 0.042,
  -0.079, -0.022, 0.004, 0.01, -0.021, -0.042, -0.052, -0.051, -0.044, 
    -0.032, -0.014, -0.001, 0.017, 0.029, 0.075,
  0.069, 0.127, 0.158, 0.099, 0.031, -0.004, -0.013, -0.012, -0.012, -0.004, 
    0.009, 0.032, 0.069, 0.097, 0.065,
  0.045, 0.07, 0.122, 0.118, 0.04, -0.005, -0.019, -0.022, -0.012, -0.007, 
    0.012, 0.025, 0.053, 0.103, 0.07,
  -0.144, -0.097, -0.103, -0.09, -0.074, -0.062, -0.054, -0.05, -0.052, 
    -0.047, -0.035, -0.012, 0.024, 0.091, 0.09,
  -0.413, -0.315, -0.27, -0.195, -0.103, -0.064, -0.057, -0.057, -0.046, 
    -0.036, -0.024, -0.001, 0.044, 0.118, 0.094,
  -0.427, -0.253, -0.198, -0.11, -0.04, -0.015, -0.006, -0.009, -0.002, 
    0.011, 0.024, 0.039, 0.076, 0.151, 0.2,
  -0.096, 0.002, 0.032, 0.04, 0.058, 0.07, 0.086, 0.109, 0.113, 0.109, 0.111, 
    0.12, 0.102, 0.105, 0.086,
  0.855, 0.307, 0.198, 0.139, 0.131, 0.143, 0.146, 0.147, 0.149, 0.155, 
    0.149, 0.143, 0.128, 0.121, 0.11,
  1.621, 0.471, 0.241, 0.174, 0.162, 0.167, 0.173, 0.18, 0.183, 0.178, 0.165, 
    0.145, 0.129, 0.103, 0.085,
  2.212, 0.546, 0.202, 0.137, 0.134, 0.136, 0.141, 0.142, 0.139, 0.132, 
    0.121, 0.104, 0.089, 0.067, 0.027,
  2.218, 0.557, 0.165, 0.11, 0.096, 0.098, 0.099, 0.098, 0.095, 0.084, 0.072, 
    0.057, 0.051, 0.054, 0.043,
  1.761, 0.473, 0.127, 0.087, 0.077, 0.074, 0.07, 0.068, 0.065, 0.067, 0.06, 
    0.051, 0.046, 0.041, 0.041,
  1.266, 0.35, 0.094, 0.064, 0.054, 0.052, 0.051, 0.052, 0.05, 0.047, 0.043, 
    0.04, 0.038, 0.038, 0.046,
  0.915, 0.26, 0.071, 0.054, 0.048, 0.045, 0.043, 0.04, 0.038, 0.037, 0.035, 
    0.033, 0.031, 0.034, 0.046,
  0.605, 0.191, 0.061, 0.051, 0.045, 0.04, 0.04, 0.04, 0.041, 0.041, 0.041, 
    0.033, 0.029, 0.052, 0.076,
  0.363, 0.103, 0.033, 0.027, 0.021, 0.019, 0.022, 0.025, 0.028, 0.031, 
    0.025, 0.046, 0.05, 0.061, 0.05,
  0.024, 0.032, 0.016, 0.012, 0.005, 0.004, 0.003, 0.004, 0.004, 0.013, 
    0.016, 0.021, 0.016, 0.033, 0.034,
  -0.195, -0.06, -0.018, -0.008, -0.002, -0.004, -0, 0.004, 0.005, 0.015, 
    0.021, 0.018, 0.021, 0.06, 0.041,
  -0.62, -0.177, -0.045, -0.022, -0.015, -0.013, -0.021, -0.025, -0.022, 
    -0.015, -0.015, 0.018, 0.064, 0.132, -124.75,
  -0.744, -0.248, -0.055, -0.04, -0.033, -0.037, -0.039, -374.641, -499.515, 
    -499.511, -0.021, 0.027, -499.479, -499.455, -499.444,
  -0.261, 0.009, 0.096, 0.034, -499.485, -124.827, 0.067, 0.074, -499.495, 
    -499.499, -374.646, -0.073, -124.936, -499.526, -499.506,
  0.312, 0.066, 0.094, 0.053, 0.039, 0.042, 0.05, 0.059, 0.067, 0.06, 0.052, 
    0.031, 0.013, -0.032, -124.9,
  0.238, 0.091, 0.068, 0.028, 0.024, 0.032, 0.04, 0.048, 0.06, 0.065, 0.07, 
    0.067, 0.055, 0.021, 0.015,
  0.007, -0.005, -0.012, -0.004, 0.004, 0.009, 0.008, 0.008, 0.004, 0.005, 
    0.005, -0.001, 0.001, -0.022, -0.003,
  -0.559, -0.092, -0.036, -0.016, -0.009, -0.002, -0.004, 0.012, 0.016, 
    0.017, -0.001, -0.017, -0.034, -0.052, -0.009,
  0.06, -0.025, -0.006, 0.001, 0.006, 0.008, 0.017, 0.013, 0.013, 0.011, 
    0.016, 0.022, 0.019, 0.028, 0.024,
  0.394, 0.093, 0.025, 0.021, 0.024, 0.025, 0.026, 0.023, 0.015, 0.009, 
    0.004, 0.003, 0.005, 0.007, 0.031,
  0.608, 0.122, 0.029, 0.022, 0.016, 0.016, 0.015, 0.015, 0.009, 0.003, 0, 
    -0.011, -0.015, -0.039, -0.01,
  0.609, 0.138, 0.043, 0.03, 0.027, 0.029, 0.026, 0.024, 0.011, 0.001, 
    -0.005, -0.018, -0.017, -0.022, -0.017,
  1.393, 0.28, 0.09, 0.06, 0.06, 0.059, 0.056, 0.05, 0.043, 0.03, 0.005, 
    -0.018, -0.031, -0.055, -0.02,
  1.951, 0.401, 0.138, 0.086, 0.074, 0.073, 0.075, 0.07, 0.06, 0.05, 0.029, 
    0.012, -0.018, -0.063, -0.062,
  2.054, 0.46, 0.181, 0.113, 0.102, 0.101, 0.1, 0.099, 0.097, 0.074, 0.049, 
    0.009, -0.007, -0.071, -0.009,
  1.303, 0.337, 0.162, 0.106, 0.093, 0.097, 0.105, 0.113, 0.107, 0.107, 
    0.088, 0.057, 0.016, -0.052, 0.022,
  -0.265, -0.006, 0.038, 0.052, 0.066, 0.074, 0.077, 0.08, 0.088, 0.078, 
    0.073, 0.061, 0.052, -0.018, 0.015,
  -1.287, -0.394, -0.164, -0.062, -0.015, 0.003, 0.014, 0.018, 0.014, 0.004, 
    0.016, 0.025, 0.021, -0.002, 0.022,
  -1.121, -0.563, -0.404, -0.218, -0.117, -0.067, -0.044, -0.038, -0.028, 
    -0.022, -0.029, -0.028, -0.014, 0.007, 0.036,
  -0.556, -0.359, -0.28, -0.182, -0.133, -0.098, -0.076, -0.063, -0.053, 
    -0.047, -0.045, -0.033, -0.021, 0.022, 0.077,
  0.017, 0.057, 0.072, 0.036, 0.004, -0.028, -0.04, -0.043, -0.04, -0.039, 
    -0.033, -0.021, -0.002, 0.023, 0.053,
  0.156, 0.234, 0.278, 0.28, 0.156, 0.078, 0.049, 0.038, 0.041, 0.041, 0.049, 
    0.063, 0.066, 0.101, 0.05,
  0.104, 0.132, 0.172, 0.157, 0.091, 0.045, 0.037, 0.045, 0.047, 0.054, 
    0.061, 0.076, 0.112, 0.114, 0.082,
  -0.192, -0.125, -0.107, -0.103, -0.082, -0.065, -0.054, -0.061, -0.059, 
    -0.06, -0.048, -0.029, 0.001, 0.067, 0.076,
  -0.533, -0.454, -0.421, -0.267, -0.161, -0.125, -0.115, -0.105, -0.102, 
    -0.091, -0.074, -0.051, -0.011, 0.062, 0.115,
  -0.857, -0.482, -0.367, -0.207, -0.085, -0.058, -0.059, -0.062, -0.058, 
    -0.042, -0.023, -0.009, 0.02, 0.078, 0.203,
  -0.849, -0.33, -0.176, -0.068, -0.026, -0.011, 0.001, 0.009, 0.02, 0.021, 
    0.033, 0.044, 0.051, 0.077, 0.038,
  0.481, 0.149, 0.108, 0.086, 0.092, 0.105, 0.118, 0.128, 0.134, 0.139, 
    0.134, 0.129, 0.103, 0.065, 0.088,
  2.217, 0.606, 0.3, 0.182, 0.156, 0.163, 0.161, 0.172, 0.168, 0.169, 0.162, 
    0.14, 0.09, 0.03, 0.024,
  2.993, 0.758, 0.282, 0.178, 0.159, 0.157, 0.162, 0.16, 0.158, 0.141, 0.13, 
    0.108, 0.071, 0.036, -0.029,
  2.829, 0.7, 0.22, 0.146, 0.13, 0.131, 0.131, 0.129, 0.124, 0.119, 0.102, 
    0.082, 0.073, 0.034, 0.023,
  2.265, 0.615, 0.171, 0.112, 0.099, 0.094, 0.092, 0.089, 0.083, 0.072, 
    0.064, 0.055, 0.039, 0.036, 0.052,
  1.392, 0.378, 0.101, 0.069, 0.057, 0.053, 0.05, 0.044, 0.04, 0.035, 0.035, 
    0.035, 0.038, 0.04, 0.06,
  0.783, 0.226, 0.062, 0.04, 0.032, 0.029, 0.03, 0.029, 0.023, 0.022, 0.02, 
    0.023, 0.023, 0.029, 0.036,
  0.415, 0.112, 0.033, 0.025, 0.02, 0.017, 0.013, 0.01, 0.014, 0.014, 0.012, 
    0.013, 0.015, 0.029, 0.041,
  0.076, 0.026, 0.011, 0.009, 0.005, 0, -0.004, -0.003, -0.005, -0.002, 
    0.003, 0.015, 0.023, 0.029, 0.042,
  -0.061, -0.03, -0.011, -0.007, -0.01, -0.009, -0.007, -0.001, 0.002, 
    -0.005, -0, 0.002, 0.009, 0.026, 0.019,
  -0.239, -0.064, -0.011, -0.008, -0.007, -0.006, -0.009, -0.018, -0.012, 
    -0.002, 0.004, 0.01, 0.02, 0.065, 0.039,
  -0.351, -0.111, -0.008, 0.005, 0.02, 0.017, 0.028, 0.029, 0.049, 0.062, 
    0.062, 0.086, 0.09, 0.161, 0.095,
  -0.578, -0.115, -0.043, -0.02, -0.005, -374.613, -374.561, 0.167, -374.632, 
    -124.901, -499.458, -499.432, -124.713, -499.481, -374.622,
  -374.26, -499.41, -499.419, -499.481, -561.931, -749.25, -749.25, -749.25, 
    -749.25, -749.25, -749.25, -561.901, -499.457, -561.918, -561.938,
  0.251, 0.111, 0.103, 0.027, -62.424, -249.735, -249.72, -249.71, -249.7, 
    -249.692, -249.71, -62.365, 0.071, -62.401, -187.307,
  -0.386, -0.062, -0.026, -0.011, -0.004, 0.001, 0.009, 0.009, 0.01, 0.008, 
    0.021, 0.031, 0.033, 0.031, 0.026,
  -0.444, -0.029, -0, -0.01, -0.002, -0.009, -0.002, -0.001, 0.012, 0.014, 
    0.029, 0.017, 0.006, -0.01, 0.021,
  -0.586, -0.117, -0.041, -0.019, -0.012, -0.005, -0.011, -0.011, -0.012, 
    -0.005, -0.014, -0.033, -0.063, -0.08, -0.028,
  -0.116, -0.029, -0.012, -0, 0.005, 0.008, 0.011, 0.009, -0.002, -0.014, 
    -0.008, -0.009, -0.009, -0.024, -0.017,
  0.421, 0.078, 0.027, 0.017, 0.018, 0.018, 0.017, 0.017, 0.01, 0.003, 
    -0.002, -0.006, -0.015, -0.012, 0.001,
  0.773, 0.175, 0.045, 0.028, 0.026, 0.024, 0.026, 0.022, 0.026, 0.023, 0.02, 
    0.009, 0.003, -0.032, -0.006,
  1.137, 0.257, 0.076, 0.048, 0.04, 0.039, 0.034, 0.031, 0.026, 0.015, 0.006, 
    -0.008, -0.006, -0.008, -0.016,
  1.796, 0.36, 0.122, 0.075, 0.068, 0.07, 0.082, 0.078, 0.073, 0.056, 0.039, 
    0.016, 0.012, -0.014, 0.004,
  2.385, 0.484, 0.171, 0.099, 0.085, 0.087, 0.087, 0.079, 0.084, 0.082, 
    0.078, 0.054, 0.037, 0.016, 0.005,
  2.427, 0.545, 0.223, 0.138, 0.12, 0.12, 0.124, 0.131, 0.13, 0.097, 0.088, 
    0.087, 0.045, -0.015, 0.004,
  1.06, 0.366, 0.191, 0.128, 0.116, 0.125, 0.135, 0.142, 0.142, 0.139, 0.124, 
    0.089, 0.057, 0.004, 0.002,
  -0.551, -0.084, 0, 0.034, 0.056, 0.061, 0.071, 0.076, 0.075, 0.08, 0.079, 
    0.092, 0.057, -0.014, 0.027,
  -1.454, -0.47, -0.234, -0.081, -0.024, -0.006, -0.003, -0.001, 0.002, 
    -0.006, -0.004, -0.008, 0.006, 0.031, 0.05,
  -1.444, -0.743, -0.505, -0.259, -0.132, -0.087, -0.074, -0.068, -0.067, 
    -0.069, -0.071, -0.07, -0.067, -0.009, 0.057,
  -0.464, -0.314, -0.26, -0.209, -0.146, -0.107, -0.09, -0.085, -0.083, 
    -0.088, -0.084, -0.082, -0.064, -0.015, 0.057,
  0.069, 0.112, 0.111, 0.117, 0.044, -0.014, -0.023, -0.021, -0.022, -0.014, 
    -0.005, -0.012, -0.014, -0.025, 0.115,
  0.311, 0.393, 0.494, 0.406, 0.188, 0.102, 0.088, 0.085, 0.085, 0.092, 
    0.092, 0.087, 0.079, 0.02, 0.061,
  0.126, 0.23, 0.292, 0.233, 0.092, 0.057, 0.048, 0.044, 0.058, 0.07, 0.092, 
    0.099, 0.118, 0.064, 0.015,
  -0.339, -0.298, -0.243, -0.182, -0.129, -0.106, -0.105, -0.103, -0.097, 
    -0.095, -0.082, -0.055, -0.007, 0.07, -0.006,
  -0.837, -0.658, -0.555, -0.316, -0.173, -0.137, -0.134, -0.132, -0.13, 
    -0.12, -0.104, -0.077, -0.02, 0.072, 0.023,
  -1.051, -0.615, -0.462, -0.26, -0.138, -0.096, -0.079, -0.079, -0.071, 
    -0.059, -0.047, -0.037, 0.026, 0.109, 0.059,
  -0.938, -0.319, -0.185, -0.067, -0.033, -0.024, -0.019, -0.01, 0.007, 
    0.014, 0.03, 0.043, 0.061, 0.102, -0.016,
  0.156, 0.036, 0.08, 0.075, 0.085, 0.09, 0.092, 0.104, 0.11, 0.104, 0.106, 
    0.087, 0.087, 0.064, -0.063,
  1.884, 0.552, 0.287, 0.174, 0.15, 0.152, 0.166, 0.17, 0.171, 0.177, 0.167, 
    0.131, 0.09, 0.052, -0,
  3.09, 0.754, 0.309, 0.184, 0.162, 0.166, 0.168, 0.173, 0.177, 0.166, 0.143, 
    0.106, 0.071, 0.029, 0.022,
  2.912, 0.744, 0.237, 0.158, 0.141, 0.138, 0.133, 0.125, 0.121, 0.106, 
    0.089, 0.072, 0.027, -0.017, -0.002,
  2.443, 0.636, 0.178, 0.113, 0.094, 0.092, 0.093, 0.093, 0.082, 0.07, 0.049, 
    0.023, -0.001, -0.021, -0.005,
  1.565, 0.421, 0.114, 0.076, 0.067, 0.06, 0.056, 0.047, 0.033, 0.025, 0.02, 
    0.017, 0.01, 0.006, 0.004,
  0.798, 0.226, 0.057, 0.04, 0.032, 0.028, 0.026, 0.023, 0.024, 0.017, 0.008, 
    0.005, 0.003, 0.004, 0.035,
  0.132, 0.023, 0.007, 0.002, -0.001, -0.002, -0.005, -0.007, -0.009, -0.011, 
    -0.005, -0.003, 0.007, 0.025, 0.034,
  -0.162, -0.061, -0.022, -0.018, -0.021, -0.024, -0.023, -0.021, -0.022, 
    -0.021, -0.018, -0.01, -0.003, 0.007, 0.004,
  -0.422, -0.125, -0.038, -0.034, -0.032, -0.032, -0.035, -0.035, -0.036, 
    -0.033, -0.027, -0.019, -0.01, 0.003, 0.022,
  -0.638, -0.195, -0.059, -0.043, -0.038, -0.037, -0.032, -0.024, -0.012, 
    -0.006, 0.006, 0.012, 0.016, 0.018, -0.001,
  -0.736, -0.248, -0.082, -0.056, -0.043, -0.026, -0.018, -0.009, -0.009, 
    -0.004, -0.004, 0.11, -187.24, 0.166, -187.272,
  -374.851, -499.577, -499.525, -499.515, -499.511, -499.52, -499.52, 
    -499.519, -499.509, -499.502, 0.179, -499.386, -686.767, -499.442, 
    -561.938,
  -374.437, -499.455, -499.504, -499.504, -499.494, -499.493, -499.487, 
    -499.483, -499.478, -499.473, 0.059, -374.613, -0.072, -374.661, -374.651,
  -0.817, -0.222, -0.046, -0.015, -0.006, 0.01, 0.04, 0.049, 0.012, -0.036, 
    -0.045, -499.504, 0.096, 0.072, 0.002,
  -1.298, -0.356, -0.19, -0.105, -0.047, -0.041, -0.037, -0.036, -0.005, 
    0.011, 0.011, 0.009, -0.004, -0.006, -0.002,
  -0.763, -0.173, -0.101, -0.043, -0.028, -0.025, -0.026, -0.029, -0.03, 
    -0.027, -0.022, -0.013, -0.02, -0.013, 0.001,
  -0.786, -0.172, -0.082, -0.037, -0.019, -0.012, -0.004, -0.001, -0.008, 
    -0.011, -0.025, -0.024, -0.029, -0.031, -0.006,
  -0.503, -0.143, -0.049, -0.016, -0.011, -0.011, -0.013, -0.015, -0.015, 
    -0.009, -0.013, -0.015, -0.022, -0.03, -0.013,
  -0.242, -0.051, -0.019, -0.004, -0.001, -0, -0, -0.004, -0.008, -0.024, 
    -0.028, -0.02, -0.018, -0.02, -0.011,
  0.384, 0.06, 0.02, 0.013, 0.014, 0.011, 0.008, 0.001, -0.008, -0.013, 
    -0.008, -0.013, -0.02, -0.026, -0.012,
  1.159, 0.238, 0.077, 0.045, 0.042, 0.041, 0.041, 0.045, 0.042, 0.031, 
    0.007, -0.003, -0.002, -0.016, -0.033,
  2.145, 0.428, 0.155, 0.088, 0.078, 0.083, 0.09, 0.083, 0.08, 0.069, 0.064, 
    0.038, 0.012, -0.024, -0.017,
  2.908, 0.59, 0.218, 0.12, 0.105, 0.104, 0.107, 0.118, 0.11, 0.104, 0.097, 
    0.076, 0.065, 0.017, -0.028,
  3.018, 0.647, 0.237, 0.133, 0.12, 0.123, 0.133, 0.116, 0.128, 0.128, 0.135, 
    0.111, 0.07, 0.037, -0.038,
  1.397, 0.459, 0.229, 0.126, 0.104, 0.104, 0.107, 0.118, 0.113, 0.107, 
    0.113, 0.108, 0.09, -0.003, -0.001,
  -1.133, -0.215, -0.036, 0.034, 0.059, 0.066, 0.071, 0.064, 0.068, 0.078, 
    0.074, 0.061, 0.043, 0.018, 0.023,
  -2.177, -0.722, -0.304, -0.083, -0.024, -0.006, 0.002, 0.012, 0.007, 
    -0.013, -0.023, -0.02, -0.019, -0.004, 0.059,
  -1.796, -0.892, -0.559, -0.279, -0.147, -0.111, -0.097, -0.099, -0.1, 
    -0.091, -0.085, -0.087, -0.089, -0.034, 0.081,
  -0.684, -0.451, -0.385, -0.217, -0.138, -0.108, -0.102, -0.103, -0.103, 
    -0.101, -0.102, -0.1, -0.095, -0.036, 0.096,
  0.124, 0.153, 0.182, 0.068, -0.014, -0.025, -0.033, -0.029, -0.027, -0.022, 
    -0.02, -0.02, -0.028, -0.02, 0.062,
  0.387, 0.475, 0.552, 0.431, 0.175, 0.108, 0.101, 0.103, 0.113, 0.121, 
    0.121, 0.112, 0.119, 0.002, 0.039,
  0.14, 0.267, 0.349, 0.257, 0.14, 0.084, 0.073, 0.079, 0.087, 0.098, 0.109, 
    0.129, 0.132, 0.074, -0.001,
  -0.417, -0.342, -0.262, -0.16, -0.095, -0.074, -0.073, -0.073, -0.071, 
    -0.052, -0.031, -0.013, 0.017, 0.074, 0.127,
  -0.948, -0.72, -0.573, -0.303, -0.172, -0.141, -0.141, -0.138, -0.141, 
    -0.131, -0.111, -0.081, -0.02, 0.057, 0.091,
  -1.293, -0.746, -0.536, -0.265, -0.149, -0.121, -0.105, -0.1, -0.097, 
    -0.091, -0.082, -0.067, -0.007, 0.093, 0.051,
  -1.115, -0.416, -0.225, -0.1, -0.052, -0.045, -0.052, -0.046, -0.037, 
    -0.024, -0.023, -0.016, 0.011, 0.073, 0.109,
  -0.093, 0.009, 0.04, 0.053, 0.054, 0.067, 0.082, 0.087, 0.093, 0.089, 
    0.091, 0.088, 0.086, 0.052, 0.132,
  2.41, 0.637, 0.33, 0.203, 0.185, 0.184, 0.182, 0.191, 0.192, 0.18, 0.166, 
    0.128, 0.077, -0.021, 0.006,
  3.531, 0.849, 0.342, 0.224, 0.195, 0.193, 0.195, 0.195, 0.188, 0.171, 
    0.142, 0.069, 0.01, -0.073, -0.01,
  3.284, 0.789, 0.259, 0.167, 0.147, 0.143, 0.143, 0.141, 0.129, 0.107, 
    0.067, 0.041, 0.014, -0.029, -0.052,
  2.591, 0.648, 0.187, 0.123, 0.107, 0.101, 0.1, 0.089, 0.079, 0.065, 0.051, 
    0.03, 0.005, -0.01, -0.034,
  1.52, 0.387, 0.102, 0.072, 0.062, 0.062, 0.057, 0.053, 0.05, 0.039, 0.025, 
    0.014, 0.008, 0.018, 0.007,
  0.993, 0.264, 0.068, 0.045, 0.035, 0.031, 0.026, 0.024, 0.017, 0.011, 0.01, 
    0.012, 0.011, 0.021, 0.026,
  0.353, 0.068, 0.01, 0.006, 0, -0.004, -0.003, -0.005, -0.006, 0.002, 0.01, 
    0.01, 0.015, 0.034, 0.022,
  -0.227, -0.075, -0.021, -0.016, -0.014, -0.017, -0.016, -0.013, -0.003, 
    -0.003, 0, 0.005, 0.018, 0.032, 0.02,
  -0.395, -0.149, -0.042, -0.027, -0.023, -0.021, -0.027, -0.026, -0.029, 
    -0.02, -0.007, -0.007, 0.018, 0.037, 0.046,
  -0.642, -0.176, -0.057, -0.046, -0.038, -0.029, -0.018, -0.012, -0.005, 
    0.002, 0.009, 0.002, 0.016, 0.058, 0.009,
  -0.752, -0.268, -0.086, -0.069, -0.061, -0.052, -0.044, -0.029, -0.029, 
    -0.023, -0.028, -0.018, 0.028, 0.072, -124.807,
  -0.528, -0.232, -0.067, -0.053, -0.055, -0.052, -0.048, -0.046, -249.768, 
    -0.004, 0.006, 0.007, 0.068, -499.412, -499.496,
  -1.378, -0.337, -499.625, -0.081, -0.049, -499.514, -499.515, -499.516, 
    -499.501, -499.501, 0.017, -124.866, -499.501, -499.498, -374.627,
  -1.273, -0.12, -0.074, -0.034, -0.027, -0.027, -0.028, -0.017, -0.006, 
    0.006, 0.046, 0.07, 0.025, -124.859, -124.871,
  -1.323, -0.305, -0.161, -0.068, -0.033, -0.025, -0.012, 0.001, 0.01, 0.01, 
    0.005, 0.012, 0.013, 0.018, 0.022,
  -0.782, -0.151, -0.077, -0.037, -0.026, -0.017, -0.008, 0.005, 0.013, 
    0.019, 0.022, 0.018, 0.018, 0.03, 0.002,
  -0.776, -0.152, -0.061, -0.02, -0.009, 0.001, 0.01, 0.011, 0.015, 0.02, 
    0.021, 0.017, 0.013, 0.006, 0.009,
  -0.52, -0.092, -0.038, -0.012, -0.002, 0.002, 0.006, 0.014, 0.014, 0.015, 
    0.009, 0.007, -0.001, -0.007, -0,
  -0.154, -0.031, -0.017, -0.006, 0, 0.002, 0.007, 0.007, 0.012, 0.008, 0.01, 
    0.004, 0.005, -0.005, -0.02,
  0.341, 0.06, 0.025, 0.021, 0.023, 0.03, 0.035, 0.038, 0.035, 0.032, 0.029, 
    0.018, 0.007, -0.003, -0.012,
  1.322, 0.261, 0.084, 0.044, 0.044, 0.044, 0.047, 0.051, 0.054, 0.053, 
    0.048, 0.038, 0.025, 0.003, -0.01,
  1.782, 0.336, 0.126, 0.069, 0.065, 0.072, 0.077, 0.078, 0.072, 0.056, 
    0.035, 0.023, 0.004, -0.031, -0.003,
  3.29, 0.627, 0.213, 0.109, 0.092, 0.087, 0.086, 0.083, 0.076, 0.066, 0.052, 
    0.024, 0.004, -0.051, -0.059,
  3.939, 0.819, 0.272, 0.143, 0.126, 0.123, 0.118, 0.114, 0.112, 0.098, 
    0.089, 0.059, 0.024, -0.033, -0.054,
  2.48, 0.656, 0.268, 0.149, 0.14, 0.146, 0.153, 0.159, 0.143, 0.13, 0.106, 
    0.084, 0.044, -0.027, 0.002,
  0.095, 0.114, 0.124, 0.103, 0.101, 0.097, 0.099, 0.104, 0.111, 0.115, 
    0.114, 0.083, 0.059, -0.017, 0.02,
  -1.819, -0.511, -0.231, -0.057, -0.007, 0.019, 0.034, 0.023, 0.03, 0.026, 
    0.028, 0.031, -0.001, -0.012, 0.032,
  -2.029, -1, -0.542, -0.207, -0.098, -0.082, -0.079, -0.069, -0.074, -0.077, 
    -0.076, -0.075, -0.054, -0.041, 0.041,
  -0.927, -0.574, -0.432, -0.235, -0.148, -0.115, -0.104, -0.111, -0.117, 
    -0.117, -0.115, -0.098, -0.081, -0.04, 0.033,
  -0.114, -0.019, 0.026, -0.03, -0.052, -0.044, -0.041, -0.042, -0.047, 
    -0.033, -0.031, -0.033, -0.047, -0.024, -0.006,
  0.28, 0.389, 0.456, 0.311, 0.111, 0.054, 0.06, 0.077, 0.108, 0.108, 0.094, 
    0.099, 0.079, 0.005, -0.049,
  0.126, 0.215, 0.273, 0.211, 0.093, 0.064, 0.058, 0.061, 0.066, 0.075, 
    0.104, 0.107, 0.11, 0.053, 0.061,
  -0.544, -0.415, -0.289, -0.173, -0.097, -0.078, -0.074, -0.067, -0.057, 
    -0.043, -0.047, -0.038, -0.003, 0.054, 0.092,
  -1.163, -0.804, -0.647, -0.306, -0.174, -0.144, -0.143, -0.14, -0.134, 
    -0.118, -0.093, -0.073, -0.028, 0.053, 0.106,
  -1.435, -0.748, -0.439, -0.194, -0.118, -0.101, -0.088, -0.085, -0.086, 
    -0.084, -0.074, -0.051, -0.004, 0.079, 0.08,
  -0.868, -0.398, -0.196, -0.058, -0.01, -0.01, -0.014, -0.017, -0.014, 
    -0.001, -0.001, 0.005, 0.032, 0.051, 0.032,
  0.837, 0.313, 0.225, 0.127, 0.108, 0.119, 0.131, 0.137, 0.135, 0.13, 0.12, 
    0.102, 0.084, 0.053, 0.074,
  2.823, 0.714, 0.363, 0.215, 0.183, 0.182, 0.186, 0.192, 0.196, 0.187, 
    0.179, 0.146, 0.1, 0.026, 0.014,
  3.992, 0.947, 0.393, 0.231, 0.197, 0.196, 0.199, 0.202, 0.193, 0.18, 0.154, 
    0.114, 0.076, -0.01, -0.03,
  3.693, 0.873, 0.292, 0.181, 0.161, 0.159, 0.157, 0.152, 0.149, 0.123, 
    0.089, 0.044, 0.016, -0.037, -0.023,
  2.692, 0.643, 0.198, 0.129, 0.11, 0.105, 0.105, 0.098, 0.09, 0.082, 0.065, 
    0.046, 0.029, 0.019, -0.016,
  1.736, 0.436, 0.122, 0.078, 0.068, 0.065, 0.062, 0.055, 0.042, 0.027, 
    0.017, 0.018, 0.009, 0.022, -0.011,
  0.947, 0.223, 0.06, 0.04, 0.036, 0.031, 0.031, 0.03, 0.028, 0.024, 0.014, 
    0.009, -0, 0.015, 0.005,
  0.42, 0.115, 0.031, 0.022, 0.018, 0.015, 0.015, 0.013, 0.003, 0.004, 0.006, 
    0.007, 0.01, 0.022, -0.002,
  0.036, -0.009, -0.008, -0.008, -0.008, -0.007, -0.002, -0.003, 0.005, 
    0.003, -0.001, 0.003, 0.02, 0.028, 0.023,
  -0.37, -0.108, -0.03, -0.019, -0.014, -0.009, -0.006, -0.002, 0.01, 0.037, 
    0.042, 0.018, 0.025, 0.05, 0.069,
  -0.667, -0.207, -0.065, -0.049, -0.04, -0.035, -0.024, -0.002, 0.016, 
    0.041, 0.061, 0.08, 0.099, 0.121, 0.097,
  -0.571, -0.219, -0.082, -0.075, -0.068, -0.065, -0.057, -0.036, -0.023, 
    -0.021, 0.075, 0.21, -62.017, 0.648, 0.836,
  -374.673, -499.519, -499.511, -499.522, -499.524, -499.524, -499.524, 
    -374.646, -374.583, 0.286, -499.453, -499.372, -61.763, -499.227, -374.542,
  -1.728, -0.459, -0.233, -0.077, -0.034, -499.506, -499.503, -499.504, 
    -499.504, -499.503, -499.506, -499.522, -686.821, -749.25, -561.938,
  -1.02, -0.369, -0.199, -0.073, -0.038, -0.04, -0.033, -0.028, -0.018, 
    -0.019, -0.015, -0.038, -187.342, -249.774, -187.384,
  -1.627, -0.461, -0.288, -0.104, -0.061, -0.05, -0.045, -0.036, -0.03, 
    -0.019, -0.017, -0.002, 0.005, 0.013, 0.012,
  -1.608, -0.388, -0.224, -0.086, -0.056, -0.048, -0.045, -0.035, -0.027, 
    -0.022, -0.011, -0.007, -0.012, 0.008, 0.016,
  -1.128, -0.315, -0.161, -0.06, -0.04, -0.034, -0.031, -0.028, -0.025, 
    -0.022, -0.019, -0.017, -0.015, -0.005, -0.008,
  -0.615, -0.151, -0.068, -0.024, -0.013, -0.009, -0.007, 0, 0.006, 0.009, 
    0.007, 0.006, 0.007, 0, 0.005,
  0.009, 0.005, 0.003, -0.002, -0.002, -0, 0.004, 0.007, 0.009, 0.011, 0.016, 
    0.015, 0.016, 0.014, 0.005,
  0.543, 0.103, 0.031, 0.01, 0.01, 0.013, 0.018, 0.022, 0.024, 0.025, 0.027, 
    0.027, 0.023, 0.015, 0.002,
  0.866, 0.156, 0.053, 0.024, 0.024, 0.026, 0.03, 0.031, 0.032, 0.033, 0.027, 
    0.022, 0.004, -0.004, -0.009,
  1.797, 0.336, 0.111, 0.053, 0.047, 0.047, 0.045, 0.045, 0.039, 0.034, 
    0.028, 0.023, 0.017, 0, -0.012,
  3.254, 0.604, 0.207, 0.097, 0.086, 0.085, 0.087, 0.084, 0.081, 0.067, 
    0.052, 0.037, 0.01, -0.029, 0.01,
  4.018, 0.809, 0.289, 0.14, 0.117, 0.11, 0.11, 0.111, 0.109, 0.094, 0.068, 
    0.036, 0.019, -0.054, 0.021,
  3.567, 0.81, 0.322, 0.171, 0.154, 0.15, 0.147, 0.151, 0.149, 0.138, 0.122, 
    0.089, 0.044, -0.023, 0.012,
  1.449, 0.471, 0.235, 0.155, 0.15, 0.152, 0.162, 0.156, 0.148, 0.14, 0.137, 
    0.115, 0.065, 0.003, 0.052,
  -0.743, -0.311, -0.094, 0.008, 0.044, 0.059, 0.063, 0.063, 0.063, 0.073, 
    0.072, 0.062, 0.038, -0.008, 0.047,
  -1.778, -0.9, -0.494, -0.172, -0.074, -0.044, -0.039, -0.033, -0.031, 
    -0.03, -0.035, -0.052, -0.048, 0.001, 0.054,
  -0.999, -0.693, -0.468, -0.233, -0.141, -0.112, -0.103, -0.094, -0.097, 
    -0.102, -0.1, -0.081, -0.058, -0.002, 0.044,
  -0.308, -0.178, -0.085, -0.061, -0.061, -0.053, -0.04, -0.046, -0.046, 
    -0.038, -0.034, -0.027, -0.029, 0.016, 0.027,
  0.156, 0.291, 0.344, 0.198, 0.069, 0.042, 0.034, 0.044, 0.057, 0.066, 
    0.085, 0.099, 0.069, 0.014, 0.053,
  0.119, 0.262, 0.26, 0.136, 0.037, 0.019, 0.024, 0.025, 0.036, 0.057, 0.061, 
    0.072, 0.075, 0.057, 0.035,
  -0.622, -0.519, -0.372, -0.185, -0.102, -0.076, -0.07, -0.067, -0.059, 
    -0.04, -0.018, -0.004, 0.012, 0.048, 0.099,
  -1.357, -0.972, -0.634, -0.257, -0.143, -0.126, -0.12, -0.113, -0.102, 
    -0.096, -0.086, -0.07, -0.023, 0.029, 0.08,
  -1.645, -0.917, -0.516, -0.2, -0.121, -0.113, -0.104, -0.101, -0.096, 
    -0.088, -0.073, -0.046, -0.004, 0.061, 0.081,
  -1.158, -0.534, -0.293, -0.102, -0.053, -0.042, -0.036, -0.02, -0.017, 
    -0.003, 0.001, 0.008, 0.03, 0.057, 0.056,
  0.338, 0.132, 0.126, 0.079, 0.069, 0.07, 0.074, 0.075, 0.078, 0.089, 0.081, 
    0.074, 0.074, 0.067, 0.032,
  2.818, 0.76, 0.374, 0.201, 0.171, 0.167, 0.171, 0.178, 0.175, 0.172, 0.155, 
    0.122, 0.08, 0.026, 0.012,
  4.043, 0.915, 0.386, 0.218, 0.188, 0.175, 0.168, 0.163, 0.148, 0.141, 
    0.109, 0.076, 0.05, 0.02, -0.037,
  3.537, 0.8, 0.299, 0.182, 0.157, 0.156, 0.153, 0.144, 0.136, 0.101, 0.073, 
    0.049, -0.003, -0.028, -0.035,
  2.664, 0.602, 0.203, 0.127, 0.109, 0.097, 0.094, 0.085, 0.069, 0.058, 
    0.037, 0.012, -0.018, -0.076, -0.025,
  1.993, 0.466, 0.147, 0.097, 0.078, 0.072, 0.065, 0.059, 0.052, 0.042, 0.03, 
    0.012, 0.007, 0.015, 0.003,
  1.218, 0.314, 0.089, 0.055, 0.044, 0.044, 0.041, 0.038, 0.035, 0.028, 
    0.022, 0.017, 0.007, 0.007, 0.007,
  0.508, 0.143, 0.04, 0.026, 0.019, 0.017, 0.017, 0.015, 0.011, 0.012, 0.005, 
    0.007, 0.008, 0.019, 0.034,
  0.182, 0.036, 0.009, 0.01, 0.008, 0.01, 0.011, 0.02, 0.022, 0.022, 0.022, 
    0.028, 0.023, 0.026, 0.055,
  -0.145, -0.055, -0.017, -0.014, -0.009, -0.006, 0.001, 0.005, 0.012, 0.023, 
    0.048, 0.046, 0.046, 0.063, 0.049,
  -0.361, -0.125, -0.041, -0.027, -0.029, -0.027, -0.015, -0.009, 0.006, 
    0.016, 0.016, 0.038, 0.079, 0.075, 0.11,
  -0.514, -0.17, -0.065, -0.047, -0.042, -0.043, -0.037, -0.025, -0.032, 
    -0.029, -0.028, 0.018, 0.004, -0.05, -124.919,
  -0.245, -0.095, -0.035, -0.035, -0.029, -0.024, -0.016, -0.024, -374.621, 
    -499.488, -499.495, -0.02, -499.523, -499.531, -499.509,
  -0.299, -0.087, 0.024, 0.004, -124.852, -499.509, -499.508, -499.505, 
    -0.031, -0.036, -499.51, -499.516, -749.25, -749.25, -561.938,
  -1.641, -0.379, -0.293, -0.124, -0.054, -0.047, -0.048, -0.049, -0.04, 
    -0.033, -0.026, -0.03, -249.764, -249.743, -187.306,
  -1.972, -0.527, -0.383, -0.145, -0.085, -0.068, -0.066, -0.058, -0.055, 
    -0.049, -0.037, -0.026, -0.013, -0.001, 0.004,
  -0.956, -0.281, -0.218, -0.078, -0.049, -0.049, -0.051, -0.051, -0.044, 
    -0.04, -0.032, -0.021, -0.021, -0.012, 0,
  -0.226, -0.085, -0.087, -0.042, -0.034, -0.037, -0.037, -0.032, -0.035, 
    -0.028, -0.025, -0.026, -0.018, -0.011, 0,
  -0.206, -0.078, -0.043, -0.019, -0.014, -0.014, -0.012, -0.014, -0.013, 
    -0.011, -0.01, -0.012, -0.014, -0.018, 0.001,
  -0.05, -0.043, -0.026, -0.013, -0.009, -0.007, -0.008, -0.003, 0, -0.002, 
    -0.004, -0.005, -0.009, -0.021, -0.021,
  0.35, 0.021, -0.009, -0.003, -0.001, 0, 0.003, 0.002, 0.002, 0.001, -0, 0, 
    -0.008, -0.022, -0.027,
  0.941, 0.139, 0.032, 0.003, 0.001, -0.001, 0.002, 0.001, -0.001, -0.004, 
    -0.011, -0.016, -0.024, -0.034, -0.045,
  1.969, 0.375, 0.129, 0.045, 0.042, 0.041, 0.042, 0.035, 0.029, 0.017, 
    0.018, 0.006, -0.006, -0.019, -0.013,
  4.173, 0.814, 0.253, 0.084, 0.066, 0.064, 0.065, 0.065, 0.057, 0.043, 
    0.022, -0.001, -0.023, -0.065, -0.057,
  5.351, 1.093, 0.372, 0.14, 0.122, 0.113, 0.103, 0.097, 0.087, 0.063, 0.036, 
    0.016, -0.008, -0.032, -0.063,
  5.829, 1.42, 0.518, 0.215, 0.183, 0.17, 0.166, 0.16, 0.149, 0.138, 0.112, 
    0.074, 0.018, -0.037, -0.038,
  3.649, 1.161, 0.48, 0.238, 0.225, 0.225, 0.241, 0.244, 0.239, 0.217, 0.19, 
    0.149, 0.08, -0.029, 0.029,
  0.162, 0.125, 0.141, 0.116, 0.141, 0.158, 0.172, 0.176, 0.171, 0.162, 
    0.156, 0.13, 0.108, 0.067, 0.081,
  -1.092, -0.556, -0.242, -0.045, 0.017, 0.038, 0.036, 0.04, 0.044, 0.041, 
    0.034, 0.054, 0.066, 0.025, 0.104,
  -0.758, -0.621, -0.372, -0.137, -0.085, -0.053, -0.036, -0.032, -0.033, 
    -0.021, -0.006, -0.007, 0.017, 0.031, 0.078,
  -0.286, -0.28, -0.185, -0.089, -0.058, -0.048, -0.032, -0.019, -0.011, 
    -0.014, -0.016, -0.022, 0.014, 0.031, 0.063,
  -0.031, 0.103, 0.176, 0.082, 0.026, 0.015, 0.017, 0.024, 0.027, 0.041, 
    0.043, 0.057, 0.08, 0.061, 0.086,
  -0.127, 0.023, 0.116, 0.019, -0.022, -0.016, -0.006, 0.001, 0.014, 0.03, 
    0.052, 0.071, 0.082, 0.079, 0.108,
  -0.533, -0.457, -0.283, -0.127, -0.083, -0.074, -0.076, -0.075, -0.07, 
    -0.054, -0.034, -0.006, 0.028, 0.064, 0.101,
  -1.281, -0.896, -0.523, -0.18, -0.094, -0.08, -0.081, -0.086, -0.081, 
    -0.073, -0.057, -0.039, -0.016, 0.041, 0.1,
  -1.461, -0.807, -0.385, -0.127, -0.067, -0.059, -0.057, -0.052, -0.052, 
    -0.055, -0.051, -0.049, -0.018, 0.037, 0.091,
  -0.948, -0.37, -0.136, -0.027, -0.009, -0.006, 0.003, 0.002, 0.001, 0.007, 
    0.009, 0.015, 0.025, 0.019, 0.033,
  0.399, 0.208, 0.147, 0.096, 0.081, 0.08, 0.08, 0.09, 0.087, 0.078, 0.076, 
    0.075, 0.064, 0.069, 0.022,
  2.094, 0.617, 0.38, 0.175, 0.14, 0.14, 0.142, 0.139, 0.134, 0.125, 0.118, 
    0.103, 0.072, 0.013, -0.007,
  2.942, 0.692, 0.338, 0.166, 0.134, 0.126, 0.12, 0.121, 0.128, 0.128, 0.117, 
    0.088, 0.046, 0.005, -0.011,
  2.742, 0.613, 0.281, 0.154, 0.13, 0.117, 0.113, 0.103, 0.092, 0.081, 0.064, 
    0.049, 0.025, 0.021, -0.004,
  2.423, 0.516, 0.198, 0.124, 0.105, 0.097, 0.094, 0.089, 0.083, 0.067, 
    0.055, 0.036, 0.023, -0.001, -0.004,
  1.799, 0.386, 0.136, 0.092, 0.076, 0.069, 0.066, 0.063, 0.059, 0.057, 
    0.048, 0.048, 0.027, 0.019, -0.001,
  1.215, 0.294, 0.09, 0.067, 0.06, 0.055, 0.054, 0.051, 0.044, 0.037, 0.025, 
    0.019, 0.01, -0.002, -0.007,
  0.75, 0.195, 0.057, 0.042, 0.034, 0.029, 0.024, 0.024, 0.024, 0.023, 0.025, 
    0.024, 0.016, 0.018, 0.022,
  0.512, 0.15, 0.044, 0.031, 0.028, 0.026, 0.024, 0.022, 0.017, 0.012, 0.011, 
    0.01, 0.01, 0.022, 0.062,
  0.328, 0.096, 0.032, 0.018, 0.013, 0.009, 0.004, 0.004, 0.002, 0.014, 
    0.009, -0.003, -0.013, -0.019, 0.034,
  0.175, 0.064, 0.012, 0.016, 0.014, 0.006, 0.003, 0, 0.005, -0.011, -0.007, 
    0.003, -0.005, 0.008, -0.02,
  -187.021, -187.236, 0.02, 0.009, 0.011, 0.016, 0.017, 0.016, -0.001, 
    -0.022, -0.039, -0.05, -0.053, -0.08, -0.069,
  -187.269, -187.312, -0.006, -0.014, -0.013, -499.506, -499.507, -0.056, 
    -374.648, -499.51, -499.513, -499.522, -499.526, -499.53, -374.643,
  -374.761, -124.716, 0.171, 0.015, -374.67, -0.107, -0.112, -124.97, 
    -499.527, -0.127, -0.148, -499.538, -499.526, -749.25, -561.938,
  -1.82, -0.3, -0.355, -0.153, -0.08, -0.074, -0.082, -0.095, -0.112, -0.108, 
    -0.106, -0.1, -0.092, -249.797, -187.349,
  -1.315, -0.303, -0.357, -0.158, -0.085, -0.083, -0.081, -0.075, -0.066, 
    -0.061, -0.055, -0.055, -0.053, -0.051, -0.016,
  -1.02, -0.151, -0.221, -0.078, -0.054, -0.064, -0.073, -0.074, -0.077, 
    -0.083, -0.078, -0.079, -0.062, -0.042, -0.023,
  -0.221, 0.088, -0.065, -0.051, -0.043, -0.047, -0.052, -0.056, -0.054, 
    -0.048, -0.037, -0.035, -0.027, -0.027, 0.011,
  0.746, 0.185, 0.023, -0.028, -0.028, -0.034, -0.04, -0.045, -0.044, -0.041, 
    -0.043, -0.042, -0.039, -0.039, -0.009,
  0.418, 0.112, -0.012, -0.026, -0.023, -0.027, -0.031, -0.033, -0.033, 
    -0.035, -0.034, -0.032, -0.03, -0.046, -0.003,
  0.366, 0.058, -0.036, -0.026, -0.023, -0.026, -0.029, -0.029, -0.03, 
    -0.028, -0.024, -0.015, -0.005, -0.011, 0,
  1.424, 0.287, 0.049, -0.004, -0.003, -0.002, -0.002, -0.001, 0, 0.002, 
    0.003, -0.011, -0.012, -0.019, 0.012,
  3.491, 0.728, 0.195, 0.035, 0.026, 0.023, 0.022, 0.017, 0.013, 0.007, 
    0.006, 0.009, 0.004, -0.007, 0.014,
  7.5, 1.571, 0.43, 0.095, 0.071, 0.063, 0.056, 0.05, 0.039, 0.027, 0.014, 
    -0.001, -0.012, -0.031, -0.007,
  13.084, 2.858, 0.732, 0.162, 0.121, 0.108, 0.102, 0.091, 0.073, 0.054, 
    0.03, 0.011, -0.012, -0.028, -0.021,
  15.538, 3.826, 0.99, 0.257, 0.199, 0.18, 0.162, 0.145, 0.132, 0.114, 0.089, 
    0.05, 0.004, -0.044, -0.044,
  13.733, 3.697, 0.932, 0.277, 0.219, 0.2, 0.185, 0.176, 0.154, 0.137, 0.118, 
    0.091, 0.052, 0.011, -0.036,
  6.567, 2.072, 0.586, 0.212, 0.201, 0.206, 0.2, 0.198, 0.182, 0.162, 0.142, 
    0.106, 0.067, 0.007, -0.012,
  -2.908, -0.907, -0.19, -0.016, 0.039, 0.055, 0.066, 0.071, 0.073, 0.077, 
    0.075, 0.058, 0.045, 0.01, 0.033,
  -4.035, -1.885, -0.553, -0.155, -0.079, -0.053, -0.037, -0.031, -0.033, 
    -0.036, -0.036, -0.03, 0.01, -0.001, 0.005,
  -2.622, -1.308, -0.421, -0.115, -0.076, -0.063, -0.059, -0.054, -0.042, 
    -0.028, -0.001, 0.024, 0.064, 0.03, 0.09,
  -0.748, -0.244, 0.004, -0.002, -0.018, -0.022, -0.022, -0.018, -0.022, 
    -0.016, -0.015, 0.028, 0.083, 0.094, 0.074,
  -1.031, -0.562, -0.162, -0.07, -0.066, -0.057, -0.049, -0.042, -0.031, 
    -0.018, -0, 0.01, 0.042, 0.008, 0.038,
  -2.468, -1.45, -0.632, -0.199, -0.099, -0.083, -0.073, -0.066, -0.057, 
    -0.042, -0.029, -0.003, 0.04, 0.043, 0.081,
  -2.442, -1.759, -0.658, -0.18, -0.09, -0.068, -0.064, -0.06, -0.052, 
    -0.044, -0.026, -0.001, 0.033, 0.083, 0.11,
  -2.056, -1.038, -0.414, -0.103, -0.057, -0.05, -0.04, -0.033, -0.026, 
    -0.016, -0.008, -0, 0.019, 0.083, 0.076,
  -0.991, -0.341, -0.077, -0.007, -0, 0.005, 0.008, 0.008, 0.006, 0.011, 
    0.011, 0.012, 0.019, 0.055, 0.086,
  0.583, 0.246, 0.124, 0.054, 0.05, 0.051, 0.053, 0.059, 0.062, 0.067, 0.075, 
    0.058, 0.055, 0.056, 0.091,
  1.144, 0.448, 0.281, 0.109, 0.081, 0.079, 0.079, 0.089, 0.083, 0.07, 0.07, 
    0.068, 0.06, 0.058, 0.062,
  1.983, 0.505, 0.284, 0.103, 0.08, 0.078, 0.081, 0.077, 0.081, 0.08, 0.077, 
    0.059, 0.044, 0.028, 0.014,
  1.675, 0.361, 0.216, 0.107, 0.082, 0.076, 0.078, 0.079, 0.072, 0.06, 0.037, 
    0.021, 0.006, 0, -0.01,
  1.608, 0.354, 0.191, 0.087, 0.069, 0.064, 0.058, 0.056, 0.047, 0.039, 
    0.031, 0.006, -0.009, -0.028, -0.017,
  1.418, 0.299, 0.134, 0.076, 0.066, 0.06, 0.055, 0.046, 0.034, 0.025, 0.01, 
    0.002, -0.006, -0.017, -0.012,
  1.223, 0.267, 0.105, 0.065, 0.054, 0.049, 0.044, 0.037, 0.032, 0.019, 0.01, 
    0.004, -0.001, -0.023, -0.015,
  0.932, 0.23, 0.072, 0.055, 0.048, 0.041, 0.033, 0.023, 0.015, 0.012, 0.01, 
    -0.001, -0.014, -0.025, -0.024,
  0.709, 0.192, 0.051, 0.047, 0.039, 0.031, 0.026, 0.02, 0.02, 0.011, 0.003, 
    0.002, -0.017, -0.015, 0.002,
  0.45, 0.152, 0.053, 0.048, 0.042, 0.034, 0.02, 0.011, 0.002, -0.009, 
    -0.011, -0.02, -0.019, -0.036, -0.065,
  0.214, 0.092, 0.027, 0.026, 0.023, 0.02, 0.028, 0.014, 0.002, -0.002, 0, 
    -0.005, -0.018, -0.008, 0.032,
  -0.011, -187.278, -249.743, -249.749, -0.01, -0.027, -0.042, -0.047, 
    -0.047, -0.05, -0.074, -0.017, -0.001, 0.334, 0.066,
  -374.789, -187.415, -249.771, -249.76, -499.504, -499.507, -499.509, 
    -124.906, -0.06, -374.656, -374.629, -249.736, -0.138, -0.103, -374.646,
  -375.353, -1.85, -1.358, -0.275, -0.118, -499.528, -124.956, -0.103, -0.1, 
    -0.104, -0.117, -0.1, -124.956, -499.497, -374.621,
  -0.607, -0.292, -0.42, -0.134, -0.079, -0.085, -0.089, -0.078, -0.062, 
    -0.053, -0.026, -0.008, 0.025, 0.016, 0.046,
  -0.78, -0.354, -0.461, -0.132, -0.071, -0.072, -0.076, -0.073, -0.072, 
    -0.061, -0.05, -0.045, -0.042, -0.007, 0.017,
  0.306, -0.11, -0.199, -0.082, -0.052, -0.055, -0.056, -0.058, -0.05, 
    -0.049, -0.039, -0.024, -0.012, -0.011, 0.016,
  0.314, 0.016, -0.103, -0.038, -0.028, -0.033, -0.038, -0.039, -0.044, 
    -0.038, -0.03, -0.014, -0, 0.026, 0.04,
  1.116, 0.236, 0.082, -0.004, -0.015, -0.022, -0.025, -0.024, -0.022, -0.02, 
    -0.016, -0.013, -0.007, 0, 0.014,
  1.527, 0.321, 0.109, 0.005, -0.005, -0.01, -0.014, -0.018, -0.022, -0.019, 
    -0.016, -0.013, -0.005, 0.001, 0.025,
  1.666, 0.327, 0.091, 0.001, -0.006, -0.012, -0.017, -0.017, -0.015, -0.011, 
    -0.001, 0.006, 0.019, 0.019, 0.025,
  2.084, 0.523, 0.189, 0.025, 0.01, 0.006, 0.007, 0.007, 0.007, 0.007, 0.003, 
    0.011, 0.014, 0.018, 0.032,
  3.538, 0.87, 0.25, 0.029, 0.015, 0.011, 0.005, 0.005, 0.002, 0.002, 0, 
    -0.004, -0.005, -0.006, -0,
  8.154, 2.038, 0.563, 0.089, 0.05, 0.041, 0.036, 0.022, 0.013, 0.005, 
    -0.002, -0.008, -0.013, -0.011, -0.002,
  15.272, 4.048, 1.086, 0.187, 0.111, 0.089, 0.073, 0.06, 0.044, 0.025, 
    0.009, -0.007, -0.018, -0.035, -0.008,
  21.165, 5.972, 1.524, 0.298, 0.182, 0.154, 0.127, 0.108, 0.091, 0.065, 
    0.045, 0.016, -0.012, -0.038, -0.046,
  21.415, 6.575, 1.589, 0.347, 0.237, 0.204, 0.18, 0.149, 0.121, 0.092, 
    0.061, 0.026, 0.01, -0.033, -0.033,
  13.372, 4.384, 1.165, 0.273, 0.193, 0.174, 0.169, 0.165, 0.157, 0.135, 
    0.104, 0.068, 0.008, -0.066, -0.06,
  -0.626, -0.167, -0.006, 0.035, 0.051, 0.072, 0.071, 0.077, 0.065, 0.053, 
    0.038, 0.026, 0.023, -0.015, -0.015,
  -7.262, -2.727, -0.576, -0.129, -0.076, -0.058, -0.049, -0.049, -0.052, 
    -0.043, -0.038, -0.027, -0.018, -0.039, -0.02,
  -7.66, -2.41, -0.559, -0.157, -0.089, -0.072, -0.071, -0.066, -0.052, 
    -0.046, -0.039, -0.025, -0.01, -0.005, -0.01,
  -4.938, -1.347, -0.28, -0.069, -0.048, -0.048, -0.04, -0.029, -0.025, 
    -0.019, -0.004, 0.003, 0.023, 0.013, 0.013,
  -8.493, -2.72, -0.542, -0.149, -0.08, -0.061, -0.053, -0.055, -0.054, 
    -0.043, -0.035, -0.012, 0.005, -0, 0.006,
  -9.22, -3.043, -0.696, -0.165, -0.079, -0.065, -0.058, -0.05, -0.034, 
    -0.024, -0.018, -0.01, 0.02, 0.025, 0.038,
  -9.01, -2.813, -0.626, -0.139, -0.065, -0.051, -0.047, -0.04, -0.037, 
    -0.033, -0.019, -0.014, -0.005, 0.001, 0.028,
  -7.216, -1.804, -0.371, -0.064, -0.024, -0.012, -0.005, -0.004, -0.002, 
    0.008, 0.01, -0.007, -0.002, 0.012, 0.009,
  -3.544, -0.967, -0.192, -0.018, 0.008, 0.015, 0.023, 0.03, 0.036, 0.032, 
    0.029, 0.034, 0.024, 0.034, 0.024,
  1.621, 0.663, 0.232, 0.062, 0.044, 0.049, 0.05, 0.052, 0.055, 0.062, 0.061, 
    0.052, 0.026, 0.049, 0.026,
  4.256, 1.218, 0.434, 0.098, 0.061, 0.057, 0.061, 0.067, 0.066, 0.062, 
    0.047, 0.03, 0.024, 0.02, 0.004,
  3.211, 0.876, 0.34, 0.076, 0.05, 0.046, 0.041, 0.037, 0.03, 0.024, 0.02, 
    0.015, 0.008, 0.017, 0.005,
  2.23, 0.554, 0.269, 0.067, 0.039, 0.033, 0.034, 0.03, 0.029, 0.019, 0.012, 
    -0.001, -0.011, -0.011, 0.031,
  1.281, 0.285, 0.165, 0.06, 0.044, 0.041, 0.039, 0.036, 0.032, 0.028, 0.017, 
    0.006, 0.011, 0.007, 0.011,
  1.042, 0.241, 0.144, 0.063, 0.05, 0.046, 0.045, 0.042, 0.031, 0.023, 0.021, 
    0.024, 0.021, 0.007, 0.004,
  0.985, 0.225, 0.128, 0.064, 0.052, 0.049, 0.048, 0.046, 0.044, 0.042, 
    0.033, 0.018, 0.004, -0.026, -0.035,
  0.992, 0.218, 0.103, 0.06, 0.049, 0.049, 0.047, 0.047, 0.046, 0.04, 0.022, 
    0.016, -0.009, -0.03, -0.017,
  0.915, 0.283, 0.111, 0.072, 0.06, 0.054, 0.053, 0.052, 0.04, 0.024, 0.022, 
    0.017, 0.003, 0.007, -0.02,
  1.165, 0.391, 0.124, 0.095, 0.086, 0.08, 0.068, 0.054, 0.048, 0.032, 0.023, 
    0.037, 0.011, -0.016, -0.055,
  0.664, 0.222, 0.073, 0.053, 0.042, 0.032, 0.024, 0.019, 0.037, 0.05, 0.038, 
    0.021, -0.009, -0.045, -0.042,
  -0.699, -62.444, 0.011, -249.709, -62.396, 0.033, 0.022, 0.002, -0.014, 
    -0.031, -0.037, -0.037, -0.045, -0.018, -187.325,
  0.001, -62.33, 0.028, -249.72, -437.045, -499.487, -499.488, -499.489, 
    -499.491, -499.493, -499.495, -499.495, -499.512, -499.519, -561.938,
  -0.366, -0.393, -0.588, -0.177, -0.095, -0.104, -0.126, -499.542, -0.063, 
    -0.06, -0.061, -124.914, -499.54, -499.554, -374.458,
  -0.198, -0.308, -0.54, -0.162, -0.096, -0.115, -0.123, -0.125, -0.111, 
    -0.098, -0.067, -0.053, -0.038, -0.048, 0.182,
  -0.523, -0.229, -0.37, -0.131, -0.084, -0.067, -0.061, -0.059, -0.081, 
    -0.09, -0.079, -0.063, -0.005, 0.013, 0.053,
  0.958, 0.171, 0.014, -0.021, -0.025, -0.03, -0.037, -0.038, -0.035, -0.029, 
    -0.012, 0.005, 0.011, 0.028, 0.046,
  1.92, 0.493, 0.302, 0.052, 0.015, 0.001, -0.006, -0.012, -0.012, -0.009, 
    -0.013, -0.006, 0.013, 0.031, 0.04,
  2.835, 0.795, 0.455, 0.075, 0.021, 0.008, -0.001, -0.007, -0.011, -0.01, 
    -0.008, -0.002, 0.007, 0.019, 0.043,
  2.666, 0.738, 0.364, 0.063, 0.021, 0.012, 0.006, 0.003, -0.001, -0.005, 
    -0.003, 0.003, 0.007, 0.024, 0.036,
  3.11, 0.898, 0.49, 0.076, 0.027, 0.017, 0.011, 0.009, 0.007, 0.01, 0.01, 
    0.015, 0.026, 0.041, 0.044,
  3.643, 1.008, 0.414, 0.06, 0.023, 0.019, 0.013, 0.007, 0.006, 0.007, 0.014, 
    0.023, 0.024, 0.025, 0.027,
  4.113, 1.215, 0.497, 0.068, 0.027, 0.018, 0.015, 0.016, 0.017, 0.016, 
    0.018, 0.014, 0.016, 0.022, 0.031,
  6.796, 1.889, 0.732, 0.101, 0.043, 0.035, 0.034, 0.035, 0.03, 0.022, 0.02, 
    0.018, 0.017, 0.022, 0.031,
  12.695, 3.898, 1.38, 0.221, 0.117, 0.099, 0.085, 0.073, 0.059, 0.052, 
    0.037, 0.028, 0.025, 0.009, 0.023,
  21.464, 6.808, 2.193, 0.357, 0.192, 0.165, 0.149, 0.127, 0.106, 0.092, 
    0.074, 0.045, 0.019, -0.025, -0.019,
  25.838, 8.642, 2.679, 0.487, 0.264, 0.227, 0.205, 0.187, 0.177, 0.146, 
    0.127, 0.083, 0.041, -0.013, -0.016,
  21.015, 7.86, 2.216, 0.417, 0.27, 0.246, 0.215, 0.184, 0.164, 0.157, 0.134, 
    0.087, 0.06, 0, -0.065,
  7.822, 2.709, 0.657, 0.171, 0.127, 0.119, 0.12, 0.123, 0.116, 0.092, 0.07, 
    0.06, 0.042, 0.011, -0.04,
  -3.3, -1.05, -0.153, -0.033, -0.023, -0.017, -0.022, -0.023, -0.018, 
    -0.018, -0.026, -0.016, 0.011, -0.013, -0.074,
  -6.332, -2.552, -0.552, -0.109, -0.055, -0.049, -0.041, -0.035, -0.032, 
    -0.026, -0.011, 0.007, 0.017, -0.005, -0.008,
  -8.749, -2.517, -0.421, -0.075, -0.038, -0.024, -0.023, -0.019, -0.007, 0, 
    -0.006, 0.003, 0.016, 0.007, -0.014,
  -6.871, -2.06, -0.445, -0.117, -0.074, -0.071, -0.064, -0.059, -0.059, 
    -0.048, -0.034, -0.021, -0.009, -0.004, -0.008,
  -6.704, -2.595, -0.666, -0.154, -0.065, -0.052, -0.041, -0.042, -0.035, 
    -0.034, -0.023, -0.009, -0.016, -0.011, -0.01,
  -6.659, -1.995, -0.364, -0.069, -0.027, -0.022, -0.023, -0.02, -0.026, 
    -0.027, -0.024, -0.028, -0.037, 0.007, -0.01,
  -4.35, -1.184, -0.22, -0.017, 0.002, 0.004, 0.01, 0.007, -0.004, -0.005, 
    -0.015, -0.03, -0.026, -0.02, -0.002,
  1.289, 0.287, 0.062, 0.029, 0.026, 0.02, 0.012, 0.008, 0.006, 0.004, 0.002, 
    -0.004, -0.016, -0.002, -0.018,
  3.724, 1.142, 0.325, 0.073, 0.033, 0.032, 0.032, 0.028, 0.022, 0.011, 
    0.001, -0.015, -0.032, -0.013, -0.014,
  5.652, 1.518, 0.457, 0.075, 0.034, 0.031, 0.029, 0.024, 0.015, 0.002, 
    -0.01, -0.028, -0.045, -0.02, -0.023,
  3.456, 0.729, 0.152, 0.017, 0.006, 0.002, -0.002, -0.012, -0.018, -0.026, 
    -0.032, -0.037, -0.051, -0.052, -0.024,
  0.693, 0.137, 0.026, -0.005, -0.007, -0.009, -0.011, -0.012, -0.018, 
    -0.026, -0.031, -0.029, -0.019, -0.022, -0.028,
  1.773, 0.382, 0.14, 0.029, 0.016, 0.012, 0.01, 0.011, 0.006, -0, -0.007, 
    -0.015, -0.015, -0.03, -0.014,
  1.827, 0.397, 0.194, 0.045, 0.028, 0.028, 0.033, 0.031, 0.026, 0.023, 
    0.022, 0.011, 0.004, -0.021, -0.028,
  2.021, 0.457, 0.22, 0.065, 0.046, 0.045, 0.048, 0.05, 0.052, 0.051, 0.039, 
    0.03, 0.01, -0.012, -0.027,
  1.58, 0.353, 0.166, 0.061, 0.049, 0.049, 0.048, 0.051, 0.051, 0.048, 0.041, 
    0.042, 0.017, -0.025, -0.059,
  1.328, 0.323, 0.149, 0.098, 0.079, 0.077, 0.074, 0.064, 0.052, 0.03, 0.015, 
    -0.01, -0.057, -0.075, -0.108,
  0.759, 0.255, 0.103, 0.075, 0.063, 0.06, 0.061, 0.059, 0.054, 0.038, 0.021, 
    0.013, 0.01, -0.019, -0.108,
  0.748, 0.459, 0.288, 0.106, 0.082, 0.054, 0.032, 0.009, -0.01, 0.048, 
    0.024, 0.017, -0.017, -0.109, -0.131,
  0.532, 0.183, 0.051, 0.063, 0.061, 0.041, 0.059, 0.035, 0.045, 0.031, 
    0.005, -0.025, -0.046, -187.384, -187.438,
  -374.422, -499.439, -499.467, -499.46, -499.477, 0.123, 0.138, 0.161, 
    -499.473, -499.471, -0.08, -0.09, -499.529, -686.82, -561.938,
  -375.153, -374.908, -0.576, -0.163, -374.664, -499.519, -499.527, -499.533, 
    -499.533, -0.121, -0.123, -0.108, -0.109, -499.532, -374.635,
  0.121, -0.123, -0.305, -0.103, -0.063, -0.067, -0.079, -0.094, -0.107, 
    -0.112, -0.117, -0.116, -0.124, -0.1, -0.058,
  -0.488, -0.293, -0.257, -0.073, -0.069, -0.087, -0.104, -0.096, -0.085, 
    -0.09, -0.081, -0.08, -0.064, -0.058, -0.021,
  1.174, 0.26, 0.061, -0.017, -0.016, -0.023, -0.025, -0.037, -0.041, -0.044, 
    -0.036, -0.033, -0.032, -0.022, -0.001,
  2.258, 0.616, 0.452, 0.085, 0.029, 0.014, 0.003, -0.009, -0.019, -0.024, 
    -0.03, -0.027, -0.012, 0.016, 0.031,
  4.256, 1.343, 0.935, 0.178, 0.063, 0.043, 0.027, 0.018, 0.008, 0.005, 
    0.001, -0.004, -0.006, -0.008, 0.003,
  3.827, 1.225, 0.825, 0.164, 0.062, 0.047, 0.04, 0.033, 0.028, 0.026, 0.019, 
    0.017, 0.016, 0.02, 0.013,
  3.695, 1.172, 0.742, 0.133, 0.05, 0.039, 0.033, 0.024, 0.019, 0.018, 0.019, 
    0.019, 0.013, 0.014, 0.014,
  3.275, 0.891, 0.476, 0.073, 0.022, 0.016, 0.01, 0.01, 0.01, 0.007, 0.004, 
    0.005, 0.005, 0.009, 0.007,
  2.827, 0.848, 0.417, 0.064, 0.024, 0.017, 0.015, 0.008, 0.007, 0.004, 
    0.006, 0.003, -0.003, -0.004, 0.005,
  4.915, 1.405, 0.715, 0.101, 0.037, 0.033, 0.026, 0.024, 0.02, 0.018, 0.003, 
    -0.006, -0.009, 0.001, 0.002,
  9.402, 2.796, 1.321, 0.188, 0.086, 0.082, 0.081, 0.073, 0.057, 0.041, 
    0.036, 0.026, 0.017, -0.013, 0.004,
  15.594, 5.263, 2.298, 0.366, 0.179, 0.156, 0.142, 0.131, 0.115, 0.106, 
    0.075, 0.04, 0.011, 0.006, -0.006,
  20.877, 7.599, 3.364, 0.532, 0.269, 0.23, 0.205, 0.184, 0.166, 0.131, 
    0.094, 0.083, 0.056, -0.009, -0.037,
  19.812, 7.47, 2.946, 0.535, 0.285, 0.236, 0.228, 0.201, 0.175, 0.146, 
    0.122, 0.105, 0.072, -0.045, -0.089,
  11.002, 4.727, 1.512, 0.284, 0.159, 0.155, 0.139, 0.114, 0.113, 0.13, 
    0.124, 0.114, 0.1, 0.068, -0.004,
  1.311, 0.471, -0.058, -0.036, -0.041, -0.028, -0.014, 0.007, 0.013, 0.008, 
    0.006, -0.001, -0.009, -0.018, -0.029,
  -8.711, -3.416, -0.699, -0.116, -0.036, -0.019, -0.009, 0, 0.013, 0.007, 
    0.015, 0.023, 0.027, 0.04, -0.009,
  -12.718, -4.094, -0.829, -0.154, -0.062, -0.039, -0.028, -0.022, -0.016, 
    -0.012, -0.018, -0.018, -0.007, 0.094, -0.004,
  -5.904, -2.341, -0.556, -0.132, -0.084, -0.082, -0.078, -0.072, -0.074, 
    -0.069, -0.053, -0.038, -0.002, 0.014, -0.032,
  -0.536, -0.249, -0.343, -0.113, -0.052, -0.037, -0.032, -0.027, -0.025, 
    -0.017, -0.014, -0.014, -0.009, -0.025, -0.045,
  -1.545, -0.508, 0.025, 0.008, 0.004, 0.002, -0.009, -0.012, -0.02, -0.033, 
    -0.041, -0.049, -0.048, -0.063, -0.047,
  0.681, 0.69, 0.341, 0.085, 0.032, 0.015, 0.003, -0.007, -0.017, -0.03, 
    -0.038, -0.044, -0.068, -0.055, -0.042,
  2.29, 0.759, 0.198, 0.029, 0.017, 0.016, 0.015, 0.01, 0.002, 0.003, 0, 
    -0.021, -0.047, -0.057, -0.046,
  1.788, 0.724, 0.254, 0.051, 0.014, 0.01, 0.004, -0.001, -0.008, -0.022, 
    -0.033, -0.044, -0.06, -0.029, -0.015,
  -1.046, -0.589, -0.295, -0.079, -0.035, -0.034, -0.038, -0.045, -0.059, 
    -0.067, -0.072, -0.072, -0.055, -0.024, -0.011,
  -1.896, -0.953, -0.4, -0.087, -0.04, -0.039, -0.04, -0.039, -0.039, -0.039, 
    -0.04, -0.042, -0.048, -0.023, -0.014,
  -0.536, -0.211, -0.13, -0.031, -0.012, -0.009, -0.008, -0.011, -0.015, 
    -0.019, -0.023, -0.024, -0.031, -0.014, 0.002,
  1.813, 0.57, 0.189, 0.021, 0.006, 0.005, 0.004, 0.002, 0, -0.003, -0.001, 
    -0.006, -0.013, -0.006, -0.006,
  2.408, 0.512, 0.226, 0.052, 0.027, 0.023, 0.021, 0.016, 0.013, 0.013, 
    0.009, -0.005, -0.009, -0.023, -0.021,
  3.14, 0.805, 0.343, 0.083, 0.053, 0.051, 0.054, 0.047, 0.045, 0.036, 0.011, 
    0.007, 0.004, -0.016, -0.037,
  2.414, 0.508, 0.261, 0.101, 0.065, 0.059, 0.061, 0.064, 0.062, 0.057, 
    0.049, 0.035, 0.013, -0.033, -0.08,
  1.679, 0.391, 0.191, 0.105, 0.086, 0.076, 0.07, 0.066, 0.056, 0.048, 0.038, 
    0.003, -0.034, -0.093, -0.144,
  0.577, 0.124, 0.107, 0.078, 0.07, 0.078, 0.08, 0.075, 0.048, 0.025, -0.026, 
    -0.043, -0.058, -0.111, -0.21,
  0.604, 0.14, 0.071, 0.076, 0.054, 0.036, 0.028, 0.003, -0.017, -0.036, 
    -0.042, -0.046, -0.042, -0.093, -0.165,
  -0.251, 0.002, 0.035, 0.043, 0.03, 0.017, 0.008, -0.01, 0.006, -0.036, 
    -0.029, -0.035, -0.087, 0.06, -437.02,
  0.106, 0.127, 0.042, 0.056, -124.828, -124.83, -499.484, -499.504, 
    -499.518, -374.674, -0.105, -499.507, -499.465, -499.421, -561.938,
  -1.912, -0.745, -375.082, -499.545, -499.521, -499.52, -0.074, -0.078, 
    -0.094, -499.527, -499.527, -499.521, -499.512, -499.529, -561.938,
  -0.838, -0.556, -0.566, -0.166, -0.106, -0.109, -0.096, -0.091, -0.072, 
    -0.07, -0.092, -0.09, -0.098, -0.076, -187.34,
  0.361, 0.169, 0.109, 0.003, -0.006, -0.02, -0.037, -0.042, -0.057, -0.057, 
    -0.044, -0.042, -0.033, -0.023, 0.003,
  1.354, 0.234, 0.078, -0.007, -0.007, -0.004, 0.002, -0.004, -0.011, -0.021, 
    -0.027, -0.02, -0.013, 0.004, 0.018,
  4.133, 1.239, 0.958, 0.197, 0.055, 0.036, 0.018, 0.006, 0.004, 0.001, 
    0.001, -0.004, -0.01, -0.008, 0.002,
  4.337, 1.344, 1.006, 0.208, 0.082, 0.063, 0.051, 0.039, 0.024, 0.012, 
    0.002, -0.003, -0.005, -0.007, -0.012,
  4.328, 1.36, 1.061, 0.212, 0.086, 0.066, 0.058, 0.05, 0.042, 0.036, 0.028, 
    0.02, 0.009, -0.003, -0.015,
  3.927, 1.301, 0.95, 0.174, 0.067, 0.056, 0.05, 0.041, 0.04, 0.034, 0.032, 
    0.02, 0.004, -0.01, -0.005,
  2.251, 0.592, 0.385, 0.055, 0.017, 0.011, 0.01, 0.007, 0.002, -0.002, 
    -0.004, -0.004, -0.007, -0.016, -0.021,
  2.13, 0.659, 0.437, 0.07, 0.019, 0.014, 0.009, 0.003, -0.001, -0.009, 
    -0.012, -0.02, -0.026, -0.028, -0.026,
  3.637, 1.017, 0.471, 0.071, 0.016, 0.009, 0.006, -0.002, -0.007, -0.009, 
    -0.013, -0.021, -0.018, -0.012, -0.003,
  7.422, 2.09, 1.076, 0.176, 0.07, 0.058, 0.05, 0.045, 0.036, 0.021, 0.004, 
    -0.005, -0.014, -0.01, -0.019,
  10.835, 3.628, 1.82, 0.258, 0.102, 0.088, 0.078, 0.066, 0.055, 0.04, 0.025, 
    0.01, -0.003, -0.025, -0.013,
  17.863, 6.618, 3.304, 0.556, 0.209, 0.168, 0.143, 0.123, 0.103, 0.082, 
    0.06, 0.033, 0.014, -0.016, -0.014,
  16.709, 6.632, 2.882, 0.506, 0.203, 0.171, 0.156, 0.142, 0.125, 0.113, 0.1, 
    0.085, 0.047, 0.022, 0.012,
  5.948, 2.89, 1.167, 0.245, 0.121, 0.096, 0.088, 0.084, 0.084, 0.08, 0.063, 
    0.054, 0.048, 0.048, 0.045,
  -3.866, -1.6, -0.376, -0.066, -0.026, -0.019, -0.006, -0.008, -0.011, 
    -0.012, -0.003, 0.001, 0.008, 0.031, 0.059,
  -8.382, -3.074, -0.595, -0.095, -0.038, -0.025, -0.019, -0.019, -0.02, 
    -0.014, -0.024, -0.022, 0.006, 0.101, 0.004,
  -9.449, -3.053, -0.811, -0.136, -0.041, -0.036, -0.041, -0.049, -0.038, 
    -0.041, -0.033, -0.005, 0.038, 0.058, -0.034,
  -5.398, -2.377, -0.723, -0.214, -0.117, -0.095, -0.075, -0.075, -0.068, 
    -0.053, -0.034, -0.033, -0.027, 0.006, -0.041,
  -1.644, -1.077, -0.474, -0.121, -0.036, -0.028, -0.034, -0.039, -0.034, 
    -0.026, -0.021, -0.013, -0.007, -0.001, -0.038,
  -0.277, 0.204, 0.232, 0.097, 0.018, 0.006, 0.012, 0.018, 0.011, 0.013, 0, 
    -0.008, -0.025, -0.055, -0.034,
  3.227, 1.059, 0.354, -0.006, -0.012, -0.004, -0.008, -0.012, -0.016, 
    -0.022, -0.023, -0.021, -0.031, -0.044, -0.032,
  3.54, 1.378, 0.604, 0.142, 0.04, 0.01, 0, -0.004, -0, 0.002, -0.002, 
    -0.019, -0.014, -0.018, -0.02,
  1.218, 0.209, -0.008, -0.004, -0.006, -0.007, -0.01, -0.012, -0.017, 
    -0.022, -0.02, -0.016, -0.02, -0.006, -0.01,
  -1.336, -0.832, -0.312, -0.077, -0.032, -0.031, -0.034, -0.038, -0.036, 
    -0.036, -0.032, -0.024, -0.005, 0.016, 0.008,
  -1.244, -0.339, -0.212, -0.045, -0.028, -0.024, -0.026, -0.029, -0.031, 
    -0.03, -0.022, -0.01, -0.009, 0.006, 0.03,
  -0.106, -0.176, -0.114, -0.025, -0.007, -0.006, -0.001, -0, 0.001, 0.002, 
    0.005, 0.002, -0.008, 0.01, 0.012,
  2.104, 0.643, 0.297, 0.06, 0.026, 0.019, 0.017, 0.013, 0.007, 0.003, 
    -0.013, -0.02, -0.008, 0.008, 0.016,
  3.544, 0.997, 0.552, 0.1, 0.048, 0.042, 0.04, 0.031, 0.012, 0.01, 0.013, 
    0.011, 0.008, -0.005, -0.014,
  3.324, 0.797, 0.49, 0.106, 0.055, 0.049, 0.051, 0.051, 0.06, 0.054, 0.05, 
    0.036, 0.013, -0.011, -0.037,
  3.534, 0.775, 0.433, 0.137, 0.081, 0.075, 0.074, 0.073, 0.066, 0.056, 
    0.045, 0.024, 0.005, -0.029, -0.028,
  2.778, 0.698, 0.359, 0.147, 0.095, 0.087, 0.083, 0.079, 0.074, 0.055, 
    0.039, 0.018, 0.003, -0.037, -0.043,
  1.518, 0.366, 0.218, 0.103, 0.08, 0.081, 0.048, 0.04, 0.029, 0.026, 0.029, 
    0.012, -0.015, -0.082, -0.079,
  0.663, 0.129, 0.059, 0.022, 0.024, 0.014, 0.023, 0.04, 0.04, 0.029, 0.001, 
    -0.056, -0.066, -0.106, -0.261,
  0.095, -249.794, -249.761, 0.08, 0.028, 0.041, 0.027, 0.004, 0.001, 0.007, 
    0.006, -0.017, -0.051, -0.135, -437.177,
  -375.348, -749.25, -749.25, -499.468, -499.475, -499.472, -499.487, 
    -499.503, -499.511, -0.043, -0.056, -374.648, -499.503, -499.601, -561.938,
  -375.026, -499.704, -499.713, -499.543, -499.517, -499.522, -499.515, 
    -499.513, -0.133, -0.123, -124.96, -499.514, -499.515, -686.811, -561.938,
  -0.224, -0.176, -0.283, -0.076, -0.035, -0.039, -0.048, -0.06, -0.064, 
    -0.084, -0.101, -0.091, -0.08, -187.329, -187.321,
  1.296, 0.332, 0.1, -0.007, -0.02, -0.022, -0.033, -0.05, -0.062, -0.063, 
    -0.029, -0.057, -0.048, -0.043, -0.008,
  1.091, 0.221, 0.199, 0.007, -0.017, -0.024, -0.027, -0.023, -0.038, -0.042, 
    -0.044, -0.041, -0.055, -0.043, -0.019,
  2.969, 0.876, 0.735, 0.158, 0.067, 0.05, 0.042, 0.029, 0.03, 0.017, 0.005, 
    -0.013, -0.022, -0.012, -0.008,
  4.443, 1.451, 1.216, 0.254, 0.114, 0.099, 0.085, 0.071, 0.045, 0.031, 
    0.014, 0, -0.013, -0.015, -0.035,
  4.684, 1.545, 1.274, 0.247, 0.102, 0.081, 0.073, 0.068, 0.058, 0.039, 
    0.025, 0.015, 0.004, -0.024, -0.034,
  3.59, 1.128, 0.844, 0.166, 0.069, 0.058, 0.052, 0.041, 0.032, 0.021, 0.007, 
    -0.002, -0.016, -0.041, -0.055,
  2.724, 0.828, 0.556, 0.109, 0.04, 0.034, 0.027, 0.02, 0.014, 0.009, 0.006, 
    -0.002, -0.024, -0.036, -0.045,
  2.51, 0.894, 0.602, 0.089, 0.021, 0.01, 0.01, 0.005, -0.001, -0.005, 
    -0.018, -0.027, -0.038, -0.048, -0.049,
  3.631, 0.967, 0.506, 0.071, 0.018, 0.013, 0.006, 0.005, -0.002, -0.011, 
    -0.017, -0.026, -0.03, -0.025, -0.026,
  6.562, 1.918, 1.132, 0.172, 0.047, 0.031, 0.024, 0.017, 0.014, 0.013, 
    0.009, 0.01, 0.002, 0, 0,
  10.122, 3.529, 1.832, 0.306, 0.099, 0.073, 0.066, 0.055, 0.046, 0.032, 
    0.028, 0.016, 0.012, 0.01, 0.013,
  14.121, 5.179, 2.712, 0.463, 0.162, 0.124, 0.103, 0.084, 0.071, 0.062, 
    0.049, 0.042, 0.026, 0.029, 0.02,
  10.54, 4.33, 2.205, 0.399, 0.145, 0.111, 0.103, 0.097, 0.088, 0.078, 0.074, 
    0.061, 0.05, 0.046, 0.031,
  5.227, 2.373, 0.962, 0.17, 0.061, 0.048, 0.038, 0.033, 0.035, 0.037, 0.036, 
    0.037, 0.031, 0.034, 0.026,
  -3.642, -1.662, -0.497, -0.132, -0.058, -0.052, -0.037, -0.034, -0.025, 
    -0.021, -0.016, -0.008, 0.01, 0.038, 0.031,
  -9.107, -3.135, -0.675, -0.122, -0.054, -0.023, -0.027, -0.026, -0.019, 
    -0.016, -0.01, -0.002, 0.01, 0.024, 0.025,
  -9.451, -3.25, -0.627, -0.096, -0.037, -0.042, -0.028, -0.028, -0.026, 
    -0.032, -0.022, -0.018, -0.002, 0.024, 0.042,
  -6.722, -2.316, -0.77, -0.211, -0.102, -0.088, -0.084, -0.085, -0.077, 
    -0.06, -0.059, -0.045, -0.027, 0.001, 0.004,
  -3.09, -1.195, -0.452, -0.098, -0.031, -0.028, -0.027, -0.027, -0.021, 
    -0.011, -0.011, -0.009, -0.007, -0.024, -0.015,
  2.799, 0.995, 0.658, 0.158, 0.033, 0.014, 0.021, 0.017, 0.015, 0.007, 
    0.006, 0.013, -0.011, -0.016, -0.049,
  3.807, 1.436, 0.381, 0.035, 0.008, 0.016, 0.021, 0.012, 0.003, 0.004, 
    0.015, -0.002, -0.016, -0.038, -0.024,
  -0.02, -0.194, 0.147, 0.073, 0.019, 0.007, 0.002, 0.005, 0.015, 0.013, 0, 
    -0.004, -0.003, -0.034, -0.01,
  1.105, 0.234, 0.146, 0.018, -0.006, -0.01, -0.008, -0.006, -0.007, -0.005, 
    -0.008, -0.013, -0.017, -0.01, 0.016,
  0.923, 0.077, -0.121, -0.04, -0.022, -0.023, -0.024, -0.028, -0.029, 
    -0.029, -0.026, -0.02, -0.018, -0.033, 0.01,
  -0.447, -0.157, -0.148, -0.034, -0.016, -0.011, -0.011, -0.013, -0.014, 
    -0.014, -0.014, -0.018, -0.002, -0.048, 0.034,
  0.383, -0.021, -0.018, -0.001, 0.008, 0.007, 0.01, 0.009, 0.011, 0.007, 
    -0.004, 0.002, -0.044, -0.017, 0.013,
  2.539, 0.841, 0.477, 0.096, 0.041, 0.031, 0.032, 0.026, 0.02, 0.026, 0.014, 
    -0.022, -0.004, 0.004, -0.034,
  4.179, 1.241, 0.705, 0.123, 0.057, 0.051, 0.047, 0.045, 0.029, 0.016, 
    0.004, 0.015, -0.004, -0.004, -0.066,
  4.341, 1.099, 0.689, 0.129, 0.065, 0.053, 0.047, 0.039, 0.03, 0.03, 0.022, 
    -0.001, -0.005, -0.011, -0.067,
  2.953, 0.674, 0.37, 0.119, 0.064, 0.062, 0.062, 0.056, 0.044, 0.027, 0.024, 
    0.011, 0.002, -0.047, -0.069,
  3.334, 0.868, 0.499, 0.14, 0.099, 0.083, 0.082, 0.074, 0.071, 0.066, 0.043, 
    0.007, -0.032, -0.049, -0.044,
  2.079, 0.567, 0.278, 0.123, 0.07, 0.063, 0.051, 0.048, 0.039, 0.023, 0.017, 
    0.004, -0.01, -0.064, -0.005,
  1.133, 0.08, 0.034, 0.024, 0.028, 0.027, 0.03, 0.021, 0.01, 0.002, -0.001, 
    -0.002, -0.023, -0.032, -124.844,
  0.36, -62.392, -187.301, 0.002, 0.005, 0.008, 0.002, 0.002, 0.011, 0.031, 
    0.056, 0.046, 0.037, -249.652, -561.859,
  -374.62, -561.948, -686.805, -499.508, -499.505, -499.502, -499.499, 
    -499.496, -499.492, -499.486, -499.483, -499.47, -499.455, -749.25, 
    -561.938,
  -1.623, -0.746, -250.428, -0.254, -0.119, -0.106, -124.964, -499.53, 
    -499.529, -499.528, -499.537, -499.538, -499.544, -499.535, -374.645,
  -0.563, -0.255, -249.949, -0.141, -0.069, -0.06, -0.056, -0.106, -0.107, 
    -0.14, -0.149, -0.135, -0.073, -0.048, -374.666,
  2.931, 0.643, 0.289, 0.021, -0.02, -0.029, -0.053, -0.022, -0.026, -0.032, 
    -0.031, -0.054, -0.054, -0.054, -0.048,
  2.402, 0.716, 0.631, 0.129, 0.072, 0.048, 0.036, 0.02, 0.034, 0.029, 0.041, 
    0.043, 0.026, 0.01, -0.014,
  3.597, 0.849, 0.753, 0.169, 0.052, 0.058, 0.054, 0.063, 0.036, 0.037, 
    0.013, 0.032, 0.013, -0.021, -0.066,
  4.359, 1.432, 1.169, 0.226, 0.095, 0.081, 0.076, 0.061, 0.053, 0.035, 
    0.007, -0.019, -0.046, -0.096, -0.102,
  3.344, 1.013, 0.872, 0.177, 0.078, 0.067, 0.067, 0.059, 0.053, 0.042, 
    0.031, 0.006, -0.018, -0.029, -0.042,
  3.494, 1.166, 0.923, 0.184, 0.072, 0.063, 0.05, 0.042, 0.037, 0.028, 0.03, 
    0.009, -0.007, -0.033, -0.043,
  2.666, 0.842, 0.562, 0.099, 0.029, 0.027, 0.026, 0.028, 0.023, 0.017, 
    0.003, -0.005, -0.02, -0.036, -0.037,
  2.371, 0.671, 0.561, 0.111, 0.043, 0.032, 0.03, 0.022, 0.013, 0.007, 
    -0.002, -0.008, -0.019, -0.028, -0.029,
  3.973, 1.28, 0.824, 0.122, 0.024, 0.014, 0.006, 0.004, -0.001, -0.009, 
    -0.011, -0.015, -0.019, -0.019, -0.01,
  6.651, 2.047, 1.159, 0.187, 0.047, 0.032, 0.025, 0.018, 0.017, 0.008, 
    0.014, 0.008, -0.001, -0.009, 0.004,
  10.481, 3.333, 1.871, 0.329, 0.108, 0.082, 0.083, 0.073, 0.064, 0.07, 
    0.056, 0.052, 0.037, 0.029, 0.03,
  13.649, 5.054, 2.995, 0.485, 0.162, 0.124, 0.11, 0.099, 0.089, 0.075, 
    0.067, 0.068, 0.049, 0.052, 0.057,
  9.792, 4.492, 2.302, 0.419, 0.154, 0.12, 0.125, 0.105, 0.099, 0.104, 0.086, 
    0.084, 0.063, 0.077, 0.02,
  6.899, 2.848, 1.255, 0.169, 0.07, 0.065, 0.063, 0.055, 0.052, 0.043, 0.038, 
    0.031, 0.032, 0.036, 0.03,
  1.733, 0.124, -0.115, -0.022, -0.019, -0.018, -0.01, -0.01, -0.019, -0.022, 
    -0.01, -0.004, -0.003, 0.039, 0.01,
  -8.022, -3.172, -0.783, -0.118, -0.057, -0.037, -0.037, -0.023, -0.023, 
    -0.025, -0.026, -0.016, -0.008, 0.01, 0.003,
  -11.657, -3.532, -0.807, -0.158, -0.056, -0.036, -0.028, -0.037, -0.039, 
    -0.039, -0.029, -0.032, -0.05, -0.038, -0.001,
  -6.321, -2.167, -0.52, -0.103, -0.027, -0.026, -0.031, -0.043, -0.041, 
    -0.04, -0.043, -0.026, -0.045, -0.036, -0.035,
  -0.895, -1.09, -0.299, 0.014, 0.009, 0.007, -0.003, -0.003, -0.006, -0.02, 
    -0.027, -0.025, -0.014, -0.012, -0.013,
  -3.264, 0.056, 0.447, 0.156, 0.071, 0.06, 0.046, 0.036, 0.031, 0.039, 
    0.048, 0.047, 0.038, -0.002, -0.053,
  4.51, 1.877, 0.824, 0.194, 0.062, 0.046, 0.045, 0.05, 0.06, 0.061, 0.046, 
    0.03, 0.033, -0.021, -0.035,
  5.3, 1.911, 0.988, 0.156, 0.036, 0.028, 0.03, 0.029, 0.026, 0.018, 0.004, 
    -0.002, -0.017, -0.04, -0.016,
  3.338, 0.945, 0.308, 0.041, -0.003, -0.012, -0.013, -0.023, -0.029, -0.024, 
    -0.013, -0.024, -0.035, -0.072, 0.001,
  1.151, 0.809, 0.583, 0.099, 0.016, -0.002, -0.014, -0.019, -0.022, -0.028, 
    -0.041, -0.039, -0.053, -0.082, -0.006,
  -1.404, -0.63, -0.378, -0.082, -0.038, -0.04, -0.042, -0.042, -0.044, 
    -0.04, -0.039, -0.056, -0.066, -0.036, -0.025,
  0.906, 0.182, 0.109, 0.006, 0.016, 0.016, 0.007, -0.003, -0.008, -0.032, 
    -0.038, -0.028, -0.026, -0.033, -0.015,
  2.603, 0.68, 0.4, 0.079, 0.025, 0.016, 0.006, -0.006, -0.006, -0.003, 
    0.004, 0.019, 0.007, 0.025, -0.076,
  3.55, 0.95, 0.717, 0.139, 0.055, 0.041, 0.046, 0.048, 0.039, 0.02, 0.023, 
    0.032, -0.013, -0.041, -0.142,
  5.392, 1.398, 0.952, 0.197, 0.086, 0.079, 0.074, 0.068, 0.065, 0.054, 
    0.035, 0.01, -0.032, -0.052, -0.154,
  3.668, 0.903, 0.621, 0.19, 0.108, 0.108, 0.105, 0.118, 0.116, 0.118, 0.095, 
    0.084, 0.041, -0.04, -0.118,
  4.019, 0.879, 0.44, 0.198, 0.132, 0.132, 0.145, 0.175, 0.141, 0.116, 0.11, 
    0.051, 0.007, 0.062, -0.057,
  3.287, 0.731, 0.305, 0.098, 0.064, 0.057, 0.046, 0.032, 0.027, 0.008, 
    0.014, 0.037, 0.02, -0.005, -124.941,
  1.338, 0.414, 0.204, 0.074, 0.045, 0.042, 0.05, 0.067, 0.068, 0.054, -0.02, 
    -0.067, -0.025, -0.054, -499.561,
  -374.24, -499.406, -499.442, -499.497, -499.505, -499.49, -499.489, 0.004, 
    0.004, -0.008, 0.007, -0.005, -124.929, -249.889, -562.028,
  -374.438, 0.043, 0.016, 0.026, 0.029, -499.493, -499.494, -499.481, 
    -499.481, -499.483, -499.515, -499.523, -499.53, -749.25, -561.938 ;
}
