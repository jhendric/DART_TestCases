netcdf cam_phis {
dimensions:
	time = UNLIMITED ; // (1 currently)
	lat = 96 ;
	lon = 144 ;
variables:
	float PHIS(time, lat, lon) ;
		PHIS:units = "m2/s2" ;
		PHIS:long_name = "Surface geopotential" ;
	double lat(lat) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
	double lon(lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
	double time(time) ;
		time:long_name = "time" ;
		time:units = "days since 1986-01-01 00:00:00" ;
		time:calendar = "noleap" ;
		time:bounds = "time_bnds" ;

// global attributes:
		:Conventions = "CF-1.0" ;
		:source = "CAM" ;
		:case = "FV1.9x2.5_no_leap-ICs-1" ;
		:title = "" ;
		:logname = "raeder" ;
		:host = "bl0312en.ucar.ed" ;
		:Version = "$Name$" ;
		:revision_Id = "$Id$" ;
		:initial_file = "caminput.nc" ;
		:topography_file = "/fis/cgd/cseg/csm/inputdata/atm/cam/topo/USGS-gtopo30_1.9x2.5_remap_c050602.nc" ;
		:landfrac_file = "/fis/cgd/cseg/csm/inputdata/atm/cam/landfrac/landfrac_1.9x2.5_gx1v4_c060922.nc" ;
		:sst_file = "/blhome/raeder/Cam3/cam3.5/models/atm/cam/bld/FV1.9x2.5-O3/sst_HadOIBl_bc_1.9x2.5_1986.nc" ;
		:history = "Wed Nov  7 12:27:34 2007: ncks -v PHIS topog_file.nc cam_phis.nc" ;
data:

 PHIS =
  27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 
    27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 
    27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 
    27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 
    27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 
    27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 
    27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 
    27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 
    27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 
    27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 
    27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 
    27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 
    27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 
    27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 
    27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 
    27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 
    27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 
    27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 
    27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 
    27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 27964.65, 
    27964.65, 27964.65, 27964.65, 27964.65,
  27186.26, 27245.15, 27303.67, 27363.11, 27424.91, 27490.52, 27561.3, 
    27638.38, 27722.55, 27814.14, 27912.97, 28018.34, 28129, 28243.3, 
    28359.21, 28474.54, 28587.04, 28694.58, 28795.25, 28887.53, 28970.3, 
    29042.91, 29105.18, 29157.33, 29199.91, 29233.77, 29259.9, 29279.37, 
    29293.22, 29302.43, 29307.8, 29309.99, 29309.46, 29306.47, 29301.13, 
    29293.38, 29283.07, 29269.93, 29253.63, 29233.83, 29210.12, 29182.15, 
    29149.53, 29111.94, 29069.13, 29020.94, 28967.35, 28908.49, 28844.69, 
    28776.46, 28704.53, 28629.78, 28553.19, 28475.81, 28398.69, 28322.74, 
    28248.71, 28177.09, 28108.07, 28041.49, 27976.82, 27913.16, 27849.26, 
    27783.51, 27714.05, 27638.77, 27555.43, 27461.75, 27355.57, 27234.98, 
    27098.55, 26945.46, 26775.71, 26590.25, 26391.09, 26181.24, 25964.7, 
    25746.23, 25531.17, 25325.07, 25133.4, 24961.22, 24812.89, 24691.81, 
    24600.3, 24539.48, 24509.25, 24508.33, 24534.39, 24584.1, 24653.36, 
    24737.44, 24831.17, 24929.18, 25026.13, 25116.95, 25197.1, 25262.82, 
    25311.27, 25340.75, 25350.71, 25341.77, 25315.62, 25274.9, 25222.89, 
    25163.36, 25100.26, 25037.48, 24978.66, 24927.01, 24885.21, 24855.34, 
    24838.82, 24836.51, 24848.63, 24874.91, 24914.6, 24966.61, 25029.51, 
    25101.73, 25181.58, 25267.36, 25357.46, 25450.41, 25544.96, 25640.09, 
    25735.02, 25829.23, 25922.41, 26014.39, 26105.15, 26194.71, 26283.09, 
    26370.27, 26456.14, 26540.53, 26623.14, 26703.63, 26781.63, 26856.79, 
    26928.82, 26997.61, 27063.19, 27125.89,
  25620.17, 25793.49, 25953.01, 26104.97, 26256.56, 26415.38, 26588.98, 
    26784.11, 27005.92, 27257.23, 27537.95, 27844.96, 28172.43, 28512.48, 
    28856.07, 29193.83, 29516.95, 29817.81, 30090.61, 30331.67, 30539.58, 
    30714.92, 30859.74, 30976.91, 31069.51, 31140.38, 31191.92, 31226.07, 
    31244.44, 31248.43, 31239.37, 31218.59, 31187.44, 31147.24, 31099.17, 
    31044.15, 30982.76, 30915.21, 30841.45, 30761.24, 30674.26, 30580.09, 
    30478.13, 30367.57, 30247.46, 30116.89, 29975.31, 29822.77, 29660.12, 
    29488.96, 29311.51, 29130.35, 28948.14, 28767.4, 28590.32, 28418.57, 
    28253.02, 28093.56, 27938.91, 27786.57, 27633, 27473.95, 27304.89, 
    27121.4, 26919.54, 26695.85, 26447.12, 26169.77, 25858.88, 25507.03, 
    25103.61, 24634.9, 24085.96, 23444.12, 22703.8, 21871.14, 20966.71, 
    20025.22, 19091.72, 18215.35, 17442.24, 16809.41, 16340.88, 16046.59, 
    15923.8, 15960.12, 16137.19, 16434.21, 16830.47, 17306.72, 17845.31, 
    18429.29, 19041.07, 19661.19, 20267.71, 20836.72, 21343.97, 21767.39, 
    22089.64, 22300.14, 22395.84, 22380.51, 22263.16, 22056.07, 21773.28, 
    21429.98, 21042.47, 20628.51, 20207.31, 19798.94, 19423.05, 19097.22, 
    18835.42, 18646.83, 18535.49, 18500.45, 18536.54, 18635.41, 18786.6, 
    18978.76, 19200.61, 19441.77, 19693.31, 19948.06, 20200.85, 20448.69, 
    20691.01, 20929.68, 21168.68, 21413.2, 21668.42, 21938.26, 22224.49, 
    22526.42, 22841.17, 23164.26, 23490.35, 23813.74, 24128.81, 24430.31, 
    24713.69, 24975.48, 25213.68, 25428.03,
  23224.47, 23717.37, 24186.37, 24630.65, 25054.25, 25464.61, 25869.36, 
    26274.06, 26683.63, 27106.53, 27557.1, 28052, 28602.28, 29206.92, 
    29852.81, 30520.95, 31193.53, 31856.21, 32494.94, 33092.34, 33629.87, 
    34095.25, 34488.6, 34820.87, 35105.77, 35351.64, 35558.45, 35720.11, 
    35828.23, 35874.65, 35852.18, 35754.41, 35576.12, 35314.75, 34973.2, 
    34563.16, 34106.54, 33632.43, 33169.26, 32735.91, 32337.26, 31966.38, 
    31611.13, 31260.24, 30906.37, 30546.27, 30179.53, 29806.99, 29429.42, 
    29046.67, 28657.53, 28260.19, 27852.96, 27434.68, 27003.94, 26556.7, 
    26082.95, 25564.11, 24973.01, 24278.3, 23453.96, 22492.31, 21413.24, 
    20259.65, 19076.85, 17889.58, 16697.04, 15490.38, 14275.01, 13076.12, 
    11925.55, 10845.76, 9844.748, 8921.265, 8071.467, 7292.27, 6583.354, 
    5950.438, 5408.041, 4978.049, 4683.716, 4542.633, 4562.133, 4737.79, 
    5054.342, 5489.032, 6017.175, 6618.163, 7279.115, 7994.639, 8763.503, 
    9584.766, 10455.85, 11373.51, 12336.34, 13346.03, 14404.31, 15504.57, 
    16620.84, 17701.66, 18675.77, 19469.08, 20022.62, 20300.92, 20289.7, 
    19991.34, 19425.47, 18632.14, 17669.94, 16605.53, 15499.53, 14397.09, 
    13326.85, 12307.1, 11355.11, 10496.39, 9770.248, 9227.747, 8919.911, 
    8878.892, 9100.168, 9536.284, 10109.38, 10739.48, 11373.25, 11995.68, 
    12619.51, 13263.33, 13934.6, 14625.81, 15320.74, 16003.1, 16661.97, 
    17293.02, 17897.37, 18478.97, 19041.61, 19587.2, 20117.22, 20635.96, 
    21150.94, 21669.04, 22191.54, 22713.02,
  22417.5, 23051.69, 23657.84, 24224.45, 24749.53, 25245.5, 25733.78, 
    26234.79, 26762.36, 27325.96, 27935.55, 28601.93, 29332.13, 30124.06, 
    30963.92, 31826.04, 32673.79, 33463.82, 34157.7, 34737.94, 35215.55, 
    35620.92, 35986.31, 36333.22, 36668.48, 36985.38, 37267.64, 37496.04, 
    37654.39, 37730.79, 37714.95, 37598.14, 37378.92, 37067.87, 36683.85, 
    36244.66, 35761.64, 35241.92, 34693.32, 34126.38, 33552.3, 32979.91, 
    32414.67, 31859.73, 31316.13, 30781.3, 30248.68, 29710.77, 29162.9, 
    28603.58, 28031.34, 27441.95, 26829.42, 26190.56, 25528.11, 24847.67, 
    24147.64, 23407.36, 22580.64, 21597.01, 20368.77, 18807.66, 16860.49, 
    14556.18, 12030.81, 9501.132, 7194.498, 5274.433, 3801.305, 2741.315, 
    2006.385, 1497.051, 1131.365, 856.2452, 644.0604, 481.7646, 362.1895, 
    282.1283, 244.6253, 261.9262, 356.0871, 552.3108, 865.1786, 1288.869, 
    1800.997, 2375.265, 2991.462, 3638.965, 4317.204, 5034.471, 5802.548, 
    6628.329, 7510.292, 8444.884, 9436.913, 10502.75, 11661.27, 12917.83, 
    14251.9, 15614.01, 16929.15, 18102.96, 19034.18, 19634.42, 19844.94, 
    19639.96, 19020.91, 18014.47, 16676.79, 15092.66, 13358.42, 11557.51, 
    9755.001, 8017.002, 6424.147, 5056.713, 3970.976, 3192.482, 2724.203, 
    2557.852, 2678.048, 3046.786, 3581.377, 4170.693, 4740.897, 5310.691, 
    5971.424, 6804.241, 7811.792, 8921.145, 10039.51, 11105.42, 12103.54, 
    13051.69, 13981.17, 14921.08, 15885.93, 16866.94, 17834.3, 18752.77, 
    19599.86, 20373.56, 21088.14, 21764.12,
  22900.21, 23649.86, 24372.21, 25051.78, 25695.37, 26345.51, 27067.86, 
    27909.95, 28866.01, 29880.32, 30880.1, 31810.36, 32647.22, 33383.53, 
    34010.47, 34516.41, 34892.64, 35135.9, 35259.56, 35310.66, 35363.2, 
    35478.56, 35672.8, 35928.18, 36221.98, 36525.68, 36792.78, 36977.77, 
    37066.95, 37078.52, 37036.94, 36954.85, 36835.46, 36685.65, 36523.71, 
    36372.84, 36241.98, 36102.16, 35883.79, 35520.01, 35003.7, 34389.06, 
    33738.59, 33082.79, 32421.09, 31740.8, 31035.08, 30315, 29606.35, 
    28928.8, 28278.85, 27635.21, 26977.06, 26296.91, 25603.24, 24913.5, 
    24237.96, 23559.23, 22821.93, 21940.28, 20806.82, 19290.23, 17242.61, 
    14551.02, 11267.03, 7758.481, 4647.438, 2433.174, 1172.14, 574.6496, 
    317.1083, 203.3765, 145.4849, 109.2428, 84.71848, 72.68057, 77.64095, 
    104.5364, 160.9121, 267.1834, 461.226, 780.9632, 1243.98, 1852.956, 
    2609.165, 3503.982, 4508.043, 5585.703, 6712.549, 7867.815, 9017.383, 
    10112.52, 11103.67, 11958, 12674.25, 13288.54, 13860.62, 14443.19, 
    15067.99, 15764.48, 16558.77, 17418.56, 18217.65, 18793.62, 19038.17, 
    18916.56, 18416.62, 17501.4, 16104.43, 14164.92, 11711.29, 8965.97, 
    6330.557, 4181.153, 2666.665, 1706.244, 1122.213, 759.0228, 531.2693, 
    412.9299, 415.9275, 578.4724, 920.5079, 1375.048, 1801.02, 2096.488, 
    2285.003, 2515.514, 3012.255, 3951.976, 5315.381, 6903.256, 8518.902, 
    10082.66, 11594.28, 13062.57, 14483.36, 15852.89, 17170.98, 18416.17, 
    19539.5, 20510.48, 21356.51, 22138.43,
  24375.65, 25461.65, 26512.56, 27520.4, 28502.48, 29464.02, 30370.13, 
    31190.95, 31944.56, 32662.08, 33343.23, 33970.46, 34534.53, 35024.33, 
    35410.25, 35655.2, 35740.34, 35679.59, 35512.07, 35268.89, 34952.03, 
    34575.61, 34211.07, 33952.5, 33842.38, 33838.41, 33851.28, 33827.71, 
    33790.04, 33796.19, 33902.33, 34152.98, 34547.62, 35024.86, 35501.45, 
    35905.61, 36186.51, 36316.96, 36268.8, 36001.98, 35520.82, 34905.21, 
    34249.77, 33605.51, 32981.43, 32368.58, 31756.07, 31132.86, 30486.59, 
    29809.34, 29101.01, 28360.47, 27582.01, 26774.54, 25976.24, 25237.66, 
    24590.59, 24019.72, 23450.85, 22770.47, 21835.97, 20433.75, 18290.58, 
    15241.83, 11429.57, 7403.327, 3983.118, 1746.911, 634.7671, 197.2689, 
    51.85196, 10.93079, 1.828578, 0.3839194, 1.204691, 6.253378, 23.55615, 
    65.73219, 149.3034, 308.0591, 598.4453, 1059.647, 1684.734, 2474.722, 
    3482.187, 4740.067, 6194.331, 7764.123, 9409.945, 11089.67, 12703.96, 
    14130.52, 15267.54, 16036.32, 16418.12, 16490.57, 16379.4, 16204.43, 
    16064.26, 16023.73, 16136.92, 16443.7, 16875.73, 17256.1, 17457.6, 
    17471.63, 17292.62, 16783.13, 15675.36, 13744.65, 11023.08, 7900.057, 
    5010.912, 2878.776, 1609.572, 961.2789, 619.5726, 385.8229, 205.1509, 
    89.77342, 52.93753, 116.1101, 315.1409, 628.2042, 930.9473, 1085.413, 
    1042.746, 888.2654, 868.71, 1307.2, 2391.373, 4041.021, 5988.839, 
    7983.176, 9907.196, 11736.23, 13464.98, 15103.35, 16681.68, 18208.38, 
    19643.18, 20948.27, 22140.88, 23270.95,
  25695.79, 27081.99, 28434.04, 29654.77, 30699.72, 31520.71, 32053.69, 
    32346.78, 32585.97, 32924.98, 33370.14, 33855.83, 34338.55, 34791.46, 
    35174.71, 35435.45, 35530.78, 35446.46, 35184.82, 34706.57, 33890.93, 
    32621.44, 30888.28, 28830.39, 26777.08, 25232.08, 24685.71, 25263.88, 
    26529.28, 27883.79, 29140.31, 30400.24, 31694.61, 32982.4, 34200.29, 
    35209.36, 35851.65, 36122.49, 36116.58, 35849.95, 35326.01, 34641.87, 
    33911.73, 33208.11, 32582.09, 32055.82, 31610.05, 31228.32, 30932.38, 
    30705.57, 30421.66, 29935.6, 29200.01, 28279.03, 27311.04, 26418.78, 
    25638.17, 24951.8, 24328.03, 23703.37, 22958.99, 21848.85, 19970.93, 
    17066.17, 13302.97, 9183.135, 5392.329, 2574.933, 958.8969, 269.6212, 
    56.44107, 9.036517, 1.17475, 0.1047391, 0.08433444, 0.7304005, 4.708305, 
    19.98744, 62.04337, 158.7266, 347.18, 636.0524, 986.334, 1413.601, 
    2070.024, 3103.514, 4512.625, 6181.769, 7943.577, 9638.643, 11166.79, 
    12470.75, 13499.92, 14183.89, 14482.26, 14461.05, 14234.91, 13838.52, 
    13197.76, 12294.03, 11317.6, 10582.96, 10361.99, 10745.95, 11534, 
    12391.6, 13146.99, 13667.44, 13550.1, 12313.25, 10040.14, 7462.203, 
    5304.062, 3958.116, 3485.002, 3573.707, 3696.702, 3428.001, 2677.082, 
    1679.085, 800.1777, 283.815, 114.918, 132.8278, 195.9278, 230.4856, 
    214.6023, 160.8648, 125.1436, 210.8089, 574.463, 1375.375, 2618.324, 
    4141.682, 5796.549, 7554.833, 9498.054, 11715.59, 14207.88, 16828.67, 
    19270.85, 21291.06, 22919.11, 24333.01,
  26185.52, 27651.14, 29120.7, 30412.91, 31437.23, 32127.64, 32465.89, 
    32588.89, 32717.69, 32937.75, 33088.46, 33037.62, 32941.87, 33024.74, 
    33322.29, 33676.79, 33866.96, 33781.04, 33428.95, 32812.12, 31838.75, 
    30403.08, 28483.4, 26040.81, 22942.09, 19761.75, 17854.79, 17750.71, 
    19026.7, 21204.26, 23747.83, 26205.99, 28461.32, 30515.07, 32282.28, 
    33645.14, 34531.73, 34967.52, 35037.45, 34761.95, 34141.4, 33271.23, 
    32280.02, 31391.42, 30876.96, 30724.14, 30731.66, 30810.19, 30935.32, 
    31038.42, 31004.07, 30680.52, 30000.06, 29072.72, 28063.38, 27082.6, 
    26182.58, 25382.43, 24689.1, 24056.15, 23344.13, 22345.94, 20812.45, 
    18533.59, 15416.45, 11616.49, 7670.764, 4249.194, 1840.859, 571.071, 
    117.8327, 16.32637, 1.791123, 0.1364987, 0, 0.001181933, 0.01550921, 
    0.424223, 3.621308, 15.08246, 37.97477, 63.84698, 78.08475, 84.70919, 
    149.7283, 443.6675, 1147.309, 2252.98, 3553.398, 4822.203, 5910.796, 
    6748.62, 7347.12, 7723.121, 7842.925, 7646.05, 7071.206, 6152.107, 
    5048.549, 3973.927, 3151.208, 2718.489, 2720.075, 3275.79, 4465.581, 
    6054.079, 7590.766, 8663.942, 9098.691, 8914.203, 8099.083, 6923.543, 
    6029.688, 5731.014, 6039.444, 6890.127, 7763.997, 8068.308, 7372.962, 
    5282.832, 2561.166, 751.8923, 130.2302, 13.46113, 0.8698198, 0.07036915, 
    0.05355769, 0.4829412, 3.47977, 19.94032, 88.40761, 288.9372, 696.6401, 
    1291.898, 1948.775, 2684.935, 3906.83, 6081.432, 9330.554, 13340.6, 
    17348.65, 20646.26, 23054.75, 24764.87,
  19172.72, 21443.09, 23994.53, 25610.28, 26418.5, 26798.1, 26777.76, 
    26235.83, 25536.28, 25224.1, 25092.02, 24929.08, 24895.7, 25242.55, 
    26055.85, 27047.21, 28137.1, 29233.13, 29908.51, 30138.54, 30075.12, 
    29402.96, 27877.7, 25922.09, 23207.86, 19396.56, 15359.48, 12231.72, 
    11318.33, 13435.39, 17997.38, 22406.66, 26002.41, 28661.9, 30574.93, 
    31999.9, 32949.11, 33460.78, 33572.46, 33259.48, 32488.85, 31517.29, 
    30520.88, 29687.08, 29314, 29273.68, 29420.7, 29862.39, 30423.46, 
    30711.77, 30735.39, 30469.81, 29804.86, 28892.29, 27881.74, 26880.95, 
    25926.21, 25037.46, 24207.38, 23412.45, 22631.31, 21805.54, 20494.58, 
    18282.35, 15186.39, 11336.48, 7519.791, 4521.761, 2282.648, 747.7747, 
    120.3773, 8.225907, 0.7941887, 0, 0, 0, 0.0007971468, 0.008256547, 
    0.2628858, 1.710443, 5.302103, 9.76335, 11.88603, 11.37717, 13.62868, 
    43.33743, 164.1795, 438.7764, 834.2753, 1249.177, 1612.015, 1868.544, 
    2042.367, 2158.712, 2192.61, 2111.001, 1849.512, 1425.859, 970.9859, 
    623.862, 454.9272, 405.9891, 420.3945, 581.6924, 1034.803, 1729.825, 
    2414.245, 2840.406, 2976.147, 2963.666, 2964.323, 3115.261, 3363.127, 
    3532.117, 3910.705, 5172.766, 7268.119, 8994.217, 9123.664, 6542.087, 
    2589.216, 519.0128, 55.0522, 1.635361, 0.1578896, 0, 0.002752773, 
    0.02851219, 0.2455015, 1.650202, 8.925238, 35.28441, 93.27203, 180.3756, 
    286.096, 408.29, 663.449, 1354.246, 3002.688, 5879.507, 9566.156, 
    13483.03, 16461.07, 17928.2,
  4313.024, 5816.496, 7901.469, 9034.239, 9318.464, 9258.712, 8874.063, 
    8038.409, 7103.399, 6592.029, 6507.513, 6949.442, 8439.663, 10964.22, 
    13637.15, 15552.31, 17741.74, 21257.65, 24662.39, 26533.11, 27165.58, 
    27326.95, 27229.59, 26220.49, 23381.56, 19273.82, 14033.77, 7838.789, 
    5190.861, 7239.552, 12747.53, 18228.61, 22831.84, 25771.91, 27599.08, 
    28849.56, 29677.69, 30259.88, 30422.1, 30074.89, 29247, 28414.46, 
    27694.52, 27194.85, 26843.95, 26575.12, 26492.11, 26647.41, 27143.28, 
    27856.96, 28219.34, 28224.57, 28004.39, 27485.4, 26641.34, 25552.45, 
    24210.3, 22599.98, 20937.7, 19434.86, 18370.57, 17859.99, 17232.6, 
    15517.73, 12701.54, 9793.259, 7024.802, 4619.617, 2560.33, 855.9818, 
    129.4445, 7.812388, 0.6848783, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.5919593, 4.488182, 12.87185, 20.50311, 21.87522, 13.37326, 
    3.296993, 0.3604679, 0.05395666, 0.02458276, 0.4456268, 4.824979, 
    37.49536, 137.891, 222.3743, 237.945, 228.8067, 195.3754, 136.8071, 
    87.71975, 63.35634, 56.18608, 64.63151, 165.9963, 617.352, 1831.066, 
    4332.24, 7937.484, 9311.427, 6820.944, 2497.599, 475.4007, 44.91589, 
    0.9601032, 0.08416811, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.06531837, 0.7450849, 
    5.638033, 35.63519, 185.484, 679.3601, 1599.286, 2617.844, 3400.24, 
    3783.76,
  644.2036, 889.1565, 1278.208, 1559.896, 1651.242, 1599.407, 1433.637, 
    1232.369, 1064.5, 986.5582, 974.1686, 1035.731, 1362.222, 2341.133, 
    3781.271, 4669.477, 5990.6, 8742.049, 11978.9, 14827.62, 17678.97, 
    20997.9, 22380.4, 21595.88, 18729.55, 14670.96, 9805.814, 4260.419, 
    1850.601, 2181.675, 4254.269, 7512.767, 11144.87, 14374.17, 16960.16, 
    18513.09, 19511.98, 20430.92, 20780.17, 20690.73, 20511.6, 20447.7, 
    20350.16, 19863.21, 18846.99, 17877.49, 17238.94, 16982.42, 17079.19, 
    18135.14, 19946.57, 20775.32, 21144.03, 21449.11, 21474.66, 20700.49, 
    18315.52, 14760.22, 11188.17, 8768.12, 7636.176, 7259.302, 6870.397, 
    5839.05, 4672.041, 4157.707, 3699.902, 2740.814, 1557.44, 508.6417, 
    71.08331, 4.343347, 0.3460977, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.0740389, 0.6459464, 1.938928, 3.104336, 3.343138, 2.016799, 
    0.4454522, 0.04990899, 0.007363489, 0.003690658, 0.05635976, 0.6642428, 
    5.154191, 20.8287, 33.82635, 35.76065, 34.75151, 31.43798, 24.42945, 
    14.94588, 9.82199, 8.680184, 10.97821, 39.22594, 173.9137, 656.759, 
    2413.631, 6239.508, 8021.936, 5696.852, 1818.486, 311.4715, 26.22496, 
    0.3794534, 0.03023658, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00816965, 0.1025249, 
    0.7771776, 4.987491, 26.26073, 99.64046, 239.8762, 394.1499, 513.128, 
    568.0305,
  0, 0, 0.0005078155, 0.006997778, 0.1163272, 0.7367138, 1.252682, 0.8104286, 
    0.1806187, 0.02244175, 0.3135114, 3.804642, 16.88047, 44.5103, 104.5338, 
    210.6332, 500.6873, 1331.913, 2812.702, 4571.016, 6497.979, 8630.35, 
    9341.724, 7968.512, 5442.454, 4377.802, 3544.312, 1856.888, 615.2691, 
    205.2272, 174.7061, 617.7067, 1873.289, 3436.563, 5122.625, 6701.429, 
    8080.928, 9118.433, 9873.976, 10331.67, 10797.7, 11703.75, 12027.35, 
    10924.5, 8509.828, 7136.96, 6315.416, 5832.227, 5803.43, 6602.431, 
    7870.045, 8372.047, 8918.041, 10337.66, 11189.47, 10673.26, 8709.469, 
    5829.629, 3078.336, 1622.868, 970.9292, 702.5196, 545.8555, 310.4319, 
    114.0817, 27.76163, 5.467812, 0.858987, 0.06233507, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.0003313541, 0.004566112, 0.1956071, 1.446218, 2.503947, 
    1.465766, 0.2558022, 0.1053435, 0.904193, 10.15138, 57.36354, 241.581, 
    956.5835, 2644.975, 3446.669, 2395.922, 700.6553, 114.4011, 9.138411, 
    0.2086599, 0.01514206, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  0, 0, 6.77799e-05, 0.001023044, 0.01621336, 0.1144704, 0.1977729, 
    0.1261899, 0.02631027, 0.003280883, 0.04184546, 0.5624956, 2.588432, 
    6.811506, 16.13963, 32.30251, 76.06861, 204.4936, 436.1432, 692.5161, 
    1089.581, 1877.08, 2177.605, 1620.103, 887.5189, 711.1821, 605.5343, 
    338.9854, 106.8159, 33.10867, 26.39963, 95.98602, 291.6489, 508.6147, 
    790.9503, 1179.764, 1604.813, 2009.515, 2372.291, 2631.253, 2914.435, 
    3431.634, 3616.469, 3114.135, 1983.219, 1378.036, 1057.467, 915.5228, 
    908.9252, 1130.728, 1525.676, 1695.996, 1954.588, 2687.721, 3125.379, 
    2923.202, 2179.797, 1187.995, 488.3473, 238.2528, 149.9181, 109.7114, 
    85.17854, 48.05018, 17.384, 4.172407, 0.8313661, 0.1291341, 0.008555546, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4.422698e-05, 0.0006675451, 0.02655648, 
    0.2245476, 0.3961303, 0.2274994, 0.03593997, 0.01614599, 0.1247067, 
    1.48698, 8.900066, 40.31473, 200.7085, 789.3536, 1223.602, 1144.888, 
    782.3504, 332.6047, 79.92854, 12.68148, 1.097704, 0.1113666, 0.03898836, 
    0.008531528, 0.001070376, 0.0001130616, 7.490692e-06, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001135151, 0.001871196, 
    0.2933303, 3.77181, 14.11033, 28.31798, 32.80766, 17.90432, 2.005178, 
    0.08103865, 0.004916167, 0, 0, 0, 0, 0, 0, 0, 0.002293951, 0.03261531, 
    0.135428, 0.2686073, 1.172866, 8.215911, 19.7438, 24.00299, 24.71234, 
    23.8788, 22.27837, 21.61855, 19.8869, 9.83814, 0.9403888, 0.04486308, 
    0.3881319, 3.702516, 7.009894, 7.338465, 6.962504, 3.66244, 0.3749718, 
    0.008415032, 0.0005104935, 0, 0, 0, 0.0006699499, 0.007215244, 
    0.01376054, 0.01443049, 0.01376054, 0.007215244, 0.0006699499, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01135449, 
    0.1871687, 6.717066, 82.56052, 353.3378, 838.8438, 1025.743, 711.491, 
    198.2725, 32.1896, 2.707453, 0.543451, 0.3767251, 0.1229696, 0.01393998, 
    0.0009847098, 5.97369e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.599066e-05, 0.0002870158, 
    0.04150159, 0.5902486, 2.249106, 4.549339, 5.290384, 2.866273, 0.2902914, 
    0.01243022, 0.0006925311, 0, 0, 0, 0, 0, 0, 0, 0.0003231445, 0.005067816, 
    0.02165641, 0.04269382, 0.1754849, 1.304499, 3.17598, 3.84675, 3.957216, 
    3.82293, 3.562867, 3.460082, 3.200881, 1.571724, 0.1333093, 0.007172065, 
    0.05561999, 0.5925216, 1.128279, 1.174432, 1.120581, 0.5860649, 
    0.05363419, 0.00129075, 7.191224e-05, 0, 0, 0, 9.437455e-05, 0.001154643, 
    0.002214911, 0.002309285, 0.002214911, 0.001154643, 9.437455e-05, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001599486, 
    0.02870912, 0.6675689, 9.522529, 75.06126, 406.6666, 662.3284, 468.7576, 
    127.9132, 20.46117, 1.973706, 2.526686, 4.004407, 2.186197, 0.1963685, 
    0.003923194, 0.01339374, 0.1806512, 0.5394768, 0.6934713, 0.695494, 
    0.3657747, 0.03166351, 0.0003920928, 2.184487e-05, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9.283473e-05, 
    0.001828027, 0.06207564, 0.8030464, 2.198592, 2.718675, 2.719725, 
    1.514571, 0.6683925, 5.29901, 9.658494, 5.285271, 0.4488438, 0.01477729, 
    0.03395966, 0.5132058, 1.560962, 2.00036, 2.013977, 1.053347, 0.0805508, 
    0.001084236, 5.506198e-05, 0, 0, 0, 0, 0,
  0.04792644, 0.04944829, 0.04792644, 0.02472415, 0.001521856, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.00203538, 0.04469763, 
    0.295601, 1.112031, 1.556278, 0.8188768, 0.05046803, 1.24695e-05, 
    5.678191e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7.986405e-05, 0.001753842, 0.01495718, 0.09819482, 
    0.1634836, 0.08689179, 0.00550568, 3.093187e-05, 1.408534e-06, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.230079e-05, 0.0002701295, 
    0.02813597, 0.5866554, 6.455871, 56.65936, 101.8061, 90.10284, 51.06049, 
    14.45378, 1.235231, 0.4683793, 0.4517413, 0.2471059, 0.1793826, 2.362316, 
    7.180734, 9.09159, 11.2123, 16.91186, 19.10843, 10.63887, 2.016544, 
    1.671056, 1.833801, 0.9595191, 0.06389478, 0.000951031, 4.330676e-05, 0, 
    0, 0, 0.001521856, 0.02472415,
  0.1482812, 0.1522212, 0.1482812, 0.07611061, 0.003939966, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.04385795, 0.922843, 
    3.11191, 4.57322, 4.889295, 2.520827, 0.1306927, 3.679783e-05, 
    1.47004e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.0002067619, 0.005175635, 0.04362213, 0.3027289, 
    0.5081891, 0.2689387, 0.0155401, 0.0002996282, 1.196987e-05, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001045335, 0.002616667, 
    0.2415794, 5.684264, 50.17545, 379.0208, 655.1815, 494.604, 146.3282, 
    22.55096, 1.008638, 0.01944646, 0.0007768684, 0, 2.877954e-07, 
    7.204055e-06, 0.4781821, 10.10358, 34.90278, 54.33404, 59.2133, 31.01679, 
    2.509005, 0.972548, 0.966929, 0.5001705, 0.0285402, 0.0004903651, 
    1.958964e-05, 0, 0, 0, 0.003939966, 0.07611061,
  0.1361185, 0.1390523, 0.1361185, 0.06952613, 0.002933725, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002215103, 0.006515329, 
    0.322533, 6.757172, 13.03208, 10.73655, 4.41509, 0.9557945, 0.03590861, 
    3.219573e-05, 1.094601e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001539562, 0.004528347, 0.03772542, 
    0.2778987, 0.4746493, 0.344362, 0.1278027, 0.07374797, 0.05096208, 
    0.02574415, 0.01890281, 0.03261318, 0.045626, 0.0237575, 0.001112949, 
    1.924223e-05, 6.542036e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002444531, 
    0.07190151, 1.577956, 34.0541, 222.501, 744.5187, 976.5635, 623.3536, 
    128.4989, 29.13472, 8.040648, 2.931512, 1.184197, 0.2164492, 0.007728054, 
    3.978266e-06, 0.3560505, 9.083056, 31.93711, 49.75407, 54.39948, 
    28.16852, 1.600645, 0.3707701, 0.3142673, 0.1202021, 0.005773611, 
    0.0001501696, 5.105514e-06, 0, 0, 0, 0.002933725, 0.06952613,
  0.06823246, 0.069372, 0.06823246, 0.034686, 0.001139536, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001074524, 0.03884725, 
    0.8476766, 18.58176, 35.4615, 20.92489, 2.772711, 0.3416718, 0.00954563, 
    1.537124e-05, 4.251719e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.980066e-05, 0.002161973, 0.01496307, 
    0.05835358, 0.235656, 0.9119001, 1.315496, 1.099961, 0.5176945, 
    0.1631588, 0.0641709, 0.1077679, 0.1519436, 0.07851037, 0.002950856, 
    6.084931e-05, 1.683106e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.005818404, 
    0.2103527, 11.16079, 315.8098, 1044.664, 1337.024, 1372.026, 741.9431, 
    78.5648, 38.18816, 28.42251, 13.21813, 3.732393, 0.5421274, 0.01499545, 
    2.876616e-06, 0.1383084, 4.460155, 15.95938, 24.88061, 27.29289, 
    14.02054, 0.541092, 0.01317933, 0.0003645433, 0, 0, 0, 0, 0, 0, 0, 
    0.001139536, 0.034686,
  0.02101068, 0.02126315, 0.02101068, 0.01063157, 0.0002524708, 0, 0, 0, 0, 
    0, 0, 0, 0.00844903, 0.3557896, 0.7031302, 0.7115793, 0.7031302, 
    0.3557896, 0.01707058, 0.3630546, 0.7165817, 0.6847982, 0.512033, 
    0.1488378, 0.00457988, 0.05620059, 1.054281, 29.02113, 55.80347, 
    29.66103, 1.57717, 0.1344037, 0.002839801, 4.505025e-06, 9.419929e-08, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.324918e-05, 0.0006336341, 0.00452559, 0.01837974, 0.2388466, 7.130684, 
    13.92852, 13.96372, 13.04031, 5.983763, 0.1893657, 0.08814278, 0.1256073, 
    0.06442416, 0.001840049, 4.774116e-05, 9.982595e-07, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.004166299, 0.1992508, 18.24148, 734.2082, 2264.723, 2788.599, 
    2840.083, 1493.061, 95.05952, 33.17323, 19.87603, 8.112919, 2.783719, 
    0.4632005, 0.009941556, 1.028544e-06, 0.03064586, 1.345777, 4.899528, 
    7.643676, 8.411407, 4.28409, 0.1159704, 0.002191166, 4.581691e-05, 0, 0, 
    0, 0, 0, 0, 0, 0.0002524708, 0.01063157,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01357099, 0.9256372, 2.746326, 
    2.774058, 2.746326, 0.9256371, 0.02878217, 1.032453, 2.740266, 2.535823, 
    1.832779, 0.5232378, 0.008443364, 0.06082897, 0.930916, 34.27751, 
    66.50745, 33.98212, 0.6632777, 0.01811019, 0.0002409436, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4.999232e-06, 0.0003757602, 0.3415694, 23.29524, 83.61237, 122.2198, 
    133.3142, 59.05472, 0.8948763, 0.03781823, 0.05554514, 0.02830629, 
    0.0005496274, 1.47553e-05, 1.963091e-07, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.00168429, 0.1265973, 12.6156, 794.9864, 2985.171, 4849.62, 5416.181, 
    2892.07, 152.0495, 12.62461, 0.2050776, 0.004345741, 9.995815e-05, 
    4.833648e-06, 6.430838e-08, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.8350303, 2.541396, 2.541396, 
    2.541396, 0.8350302, 0, 0.9359525, 2.537376, 2.329607, 1.687663, 
    0.4681671, 0, 0.04156165, 0.3206185, 25.41992, 50.04424, 25.06427, 
    0.0288688, 0.002886881, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 61.31417, 122.6283, 110.2689, 69.99321, 
    18.29769, 0, 8.385805e-05, 0.000646905, 14.95389, 149.5271, 813.4948, 
    1190.372, 658.1776, 43.12158, 4.367698, 0.07345625, 0.1769785, 0.2276383, 
    0.1138191, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.06191495, 0.6191495, 
    552.5746, 2510.801, 5559.89, 6678.021, 3809.328, 322.1697, 32.30903, 
    0.04383782, 0.004399965, 7.705145e-06, 7.705149e-07, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3549694, 1.080342, 1.080342, 
    1.080342, 0.3549694, 0, 0.3978712, 1.078632, 0.9903104, 0.7174214, 
    0.1990167, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 258.4443, 516.8886, 455.0822, 
    266.6425, 67.41572, 0, 0, 0, 21.01506, 210.1506, 2011.937, 3410.235, 
    2225.024, 356.1162, 35.91751, 0.3780788, 0.7149077, 0.8797389, 0.4398694, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 115.3018, 1153.018, 5304.901, 
    7242.988, 4790.614, 800.8521, 80.31123, 0.1076154, 0.01076155, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0926432, 0.2819576, 0.2819576, 
    0.2819576, 0.09264319, 0, 0.1038401, 0.2815115, 0.2584604, 0.1872393, 
    0.05194123, 0, 0, 0, 0, 0, 0.009834385, 0.02993074, 0.02993074, 
    0.02993074, 0.009834385, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.08482186, 0.8482186, 277.3235, 552.1702, 470.2016, 
    238.2391, 56.07396, 0, 0, 0, 16.03948, 160.3948, 1609.068, 2749.782, 
    2288.183, 1038.106, 297.6017, 37.36808, 4.838406, 0.52457, 0.05245703, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 97.04083, 970.4084, 5297.848, 
    7762.104, 5560.417, 1155.333, 128.9432, 6.456263, 0.866859, 0.1053488, 
    0.01053488, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.05965352, 
    0.119307, 0.05965352, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.05568269, 0.1694691, 0.1694691, 0.1694691, 0.05568269, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.087032, 
    10.87032, 300.5141, 569.2869, 454.0257, 155.7347, 27.06052, 0, 0, 0, 0, 
    0, 25.93337, 259.3337, 1164.493, 1571.732, 1011.037, 154.2265, 15.42266, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 89.78883, 897.8884, 
    5418.049, 8214.264, 6166.393, 1473.196, 312.7854, 79.6984, 10.80504, 
    1.350094, 0.1350095, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.4797766, 0.9595532, 0.4797766, 0, 0,
  0, 0, 0, 0, 0, 0.0003308039, 0.003308039, 1.003899, 1.998138, 1.055043, 
    0.03833825, 0.003833827, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.06815077, 0.2074154, 0.2074154, 0.2074154, 0.06815077, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.8867506, 2.698806, 2.602208, 2.290953, 0.7043344, 
    2.765588e-05, 3.585023e-06, 0, 0.07132614, 0.7132983, 7.920724, 64.22765, 
    584.1025, 982.3037, 829.3174, 402.8799, 92.58968, 0, 0, 0, 0, 0, 
    6.206638, 62.06639, 805.578, 1429.922, 923.5585, 142.8749, 14.2875, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 64.93711, 649.3712, 5611.286, 
    9326.408, 6734.803, 1695.047, 768.028, 437.1914, 90.94247, 6.027653, 
    0.6035296, 0.0003637868, 3.637869e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.03398576, 0.2980051, 1.145763, 1.483293, 0.7416465, 0, 0,
  0, 0, 0, 0, 0, 0.004564434, 0.04564435, 13.8518, 27.57033, 14.55749, 
    0.5289915, 0.05289917, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.07102577, 0.2161654, 0.2161654, 0.2161654, 0.07102577, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 12.23539, 37.23814, 35.90528, 31.61059, 9.71841, 
    0.0003815961, 4.946617e-05, 0, 0.9841585, 9.842094, 54.0905, 334.2164, 
    1408.636, 2471.152, 2496.967, 2507.191, 820.2721, 0, 0, 0, 0, 0, 
    1.330092, 13.30092, 263.1144, 487.3901, 323.5926, 54.72433, 5.472435, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24.57593, 245.7593, 5789.094, 
    10860.57, 7420.854, 1890.907, 1167.288, 866, 258.0073, 27.13439, 
    2.723981, 0.005019533, 0.0005019535, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.6152425, 1.872477, 1.872477, 1.872477, 0.6152424, 0, 0,
  0, 0, 0, 0, 0, 0.1283997, 1.283997, 245.9631, 761.6099, 798.4694, 805.9808, 
    371.1477, 58.23775, 5.823777, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.05729815, 0.1743857, 0.1743857, 0.1743857, 0.05729815, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 43.49913, 174.6985, 308.405, 353.2078, 231.8634, 
    50.84431, 15.4279, 3.881383, 26.02835, 131.2251, 571.3605, 1189.86, 
    1715.097, 2242.421, 3019.589, 3283.998, 1656.792, 10.13308, 1.016045, 
    0.001492281, 0.0001934439, 0, 0.5633195, 5.635185, 60.37441, 104.2911, 
    69.33343, 11.77251, 1.177251, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.02072012, 0.2072012, 9.135916, 87.00794, 5968.845, 11684.1, 8583.214, 
    2356.971, 1175.486, 744.048, 361.1835, 180.532, 38.27143, 2.443168, 
    0.2443169, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.4963304, 1.510571, 
    1.510571, 1.510571, 0.4963304, 0, 0,
  0, 0, 0, 0, 0, 1.711431, 17.11431, 1664.908, 5766.028, 7421.696, 7892.278, 
    4186.731, 872.8389, 87.28393, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 91.77586, 624.8071, 
    2078.208, 2648.577, 2057.986, 605.1616, 170.9187, 94.72673, 511.7992, 
    1139.142, 1678.019, 1840.485, 1833.359, 1826.232, 2720.288, 3614.343, 
    1991.329, 126.1406, 12.62822, 0.007720958, 0.001000865, 0, 0.8579454, 
    3.93457, 8.806867, 10.59856, 5.299281, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.1072044, 1.072044, 6.437263, 41.8597, 6182.193, 12244.63, 
    10026.11, 4174.647, 1174.806, 429.4693, 744.8412, 899.1722, 502.705, 
    36.3828, 3.638282, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 10.98548, 109.8548, 2337.88, 7764.558, 10856.66, 11778.21, 
    9115.008, 5030.763, 1201.502, 2.206624, 0.2206625, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0007992755, 
    0.007992755, 169.7217, 1032.166, 3156.549, 3982.457, 3394.681, 1826.19, 
    926.024, 672.563, 1036.512, 1513.166, 1675.918, 1697.789, 1641.187, 
    1613.488, 2592.993, 3572.499, 2440.581, 448.178, 44.82587, 0.008221637, 
    0.007612157, 0.007521384, 0.4045719, 1.44726, 2.022471, 2.206553, 
    0.8655198, 0.02647949, 0.02647949, 0.02647949, 0.01323975, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.02310508, 0.04621016, 0.02310508, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.06289042, 0.1257808, 0.06289042, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.08880578, 0.8880579, 4.062661, 21.97739, 7360.334, 14658.54, 12017.8, 
    5029.871, 1332.535, 380.7867, 1102.881, 1456.247, 1137.227, 327.7094, 
    45.18504, 0.07382406, 0.007382409, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0,
  0, 0, 0, 0, 0, 80.3664, 803.664, 3784.258, 8435.926, 11688.1, 13431.32, 
    13136.49, 11766.06, 3633.436, 38.84134, 3.884136, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01315869, 
    0.1315869, 262.8175, 1408.721, 3834.983, 4763.228, 4353.915, 3287.951, 
    2929.32, 2624.792, 2127.319, 1642.202, 1175.525, 912.8866, 1038.762, 
    1458.96, 2695.156, 3182.863, 2536.204, 864.1663, 149.0583, 0.002448812, 
    0.01516862, 0.04653164, 0.05798198, 0.0616147, 0.02024483, 0, 0.05544777, 
    0.1687541, 0.1687541, 0.1687541, 0.05544777, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1346276, 0.2692552, 0.1346276, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.3664469, 0.7328939, 0.3664469, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.580448, 15.80448, 9039.223, 18032.3, 14561.9, 5531.103, 1382.211, 
    427.3053, 1061.44, 1976.815, 2642.521, 2849.429, 1274.538, 1.215386, 
    0.1215386, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 409.0002, 2403.878, 6002.959, 9703.585, 12104.51, 13212.61, 
    12958.42, 11628.83, 3667.239, 94.93795, 12.48615, 0.2060911, 42.2706, 
    84.3351, 49.71484, 5.169377, 0.5169379, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0599484, 0.599484, 328.5462, 1670.151, 
    4300.141, 5297.01, 4812.155, 4327.3, 4466.051, 4604.802, 3963.276, 
    2240.267, 1324.843, 863.774, 1122.358, 1635.59, 2631.75, 3007.15, 
    2381.761, 774.28, 126.3984, 0.0004918285, 0.01943007, 0.03836832, 
    0.03279382, 0.01690868, 0.004017588, 0, 0.04712962, 0.143438, 0.143438, 
    0.143438, 0.04712961, 0, 0, 0, 0, 0, 0, 0, 0.002943106, 0.02943106, 
    0.1671345, 0.2483303, 0.1241651, 0, 0.005292299, 0.0105846, 0.008485228, 
    0.003152673, 0.001541, 0.0007570874, 0.0001308866, 0, 0, 0, 0.3348258, 
    0.6696516, 0.3348258, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0003395319, 
    0.003395319, 0.6898205, 6.826903, 9016.851, 18013.78, 15690.57, 8888.089, 
    2682.515, 669.7019, 1093.885, 2464.908, 4187.626, 4794.69, 2434.072, 
    25.188, 2.606315, 0.04167336, 0.004167338, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0,
  0, 0, 0, 0, 0, 1113.582, 4692.732, 8423.42, 11168.21, 11600.92, 11664.81, 
    11413.59, 10099.92, 3336.544, 202.5337, 28.27975, 2.327028, 577.5411, 
    1152.755, 714.869, 94.85712, 9.485716, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1311426, 1.311426, 356.9771, 1774.877, 
    4469.311, 5486.503, 5096.334, 4706.165, 5414.053, 6121.942, 5416.627, 
    3373.814, 1592.175, 1022.672, 1671.231, 3015.525, 3086.993, 3130.839, 
    1330.364, 165.2247, 16.52164, 0, 0.002677361, 0.00814849, 0.00814849, 
    0.00814849, 0.002677361, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.1255576, 0.2511151, 0.1981523, 0.06249677, 0.009815964, 0, 0.03527779, 
    0.07055558, 0.05656145, 0.02101532, 0.01027211, 0.005046648, 
    0.0008724733, 0, 0, 0, 0.08615055, 0.1723011, 0.08615055, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0.01448497, 0.02896993, 0.01547536, 0.001980784, 6359.022, 
    19353.54, 18865.88, 17390.88, 6262.19, 824.934, 1311.758, 2901.291, 
    5258.717, 6120.86, 3625.754, 387.8117, 40.38705, 0.7646985, 0.07646988, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0.07207831, 0.7207831, 1671.867, 6468.716, 10476.02, 11798.39, 
    11436.25, 10372.34, 9970.814, 9041.456, 3576.532, 361.6147, 49.70304, 
    3.248103, 1319.525, 2635.802, 1894.614, 403.0852, 60.89, 10.34525, 
    2.720905, 0.813978, 0.1156648, 0.01631759, 0.00163176, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1260166, 1.260166, 340.8816, 1705.791, 
    4328.974, 5320.716, 4966.01, 4611.304, 5327.546, 6043.788, 5441.552, 
    3649.521, 1909.913, 1334.936, 2017.494, 3412.285, 3225.934, 2521.503, 
    773.2611, 36.80882, 4.775006, 0.004011612, 15.80082, 31.59763, 17.88423, 
    1.435843, 0.158043, 0.01191227, 0.01312833, 0.01566495, 0.02172979, 
    0.02647408, 0.02569876, 0.02131886, 0.00619116, 0, 0.03606902, 
    0.07213805, 0.03705403, 0.001970011, 0.1169505, 0.2319311, 0.1325428, 
    0.01355373, 0.002038257, 0.0003231864, 0.03266844, 0.06501369, 
    0.05165879, 0.01801698, 0.008827461, 0.004734324, 0.0008519955, 0, 0, 0, 
    0.01769033, 0.03538066, 0.01769033, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.01262423, 0.02524847, 0.0128276, 0.0004067382, 5111.094, 17676.06, 
    22096.62, 23430.28, 8650.817, 1077.241, 1524.544, 2981.02, 5170.587, 
    5973.787, 5072.782, 2547.534, 700.1508, 55.51641, 5.550865, 0, 
    0.003463103, 0.006926205, 0.003463103, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 1.503165, 15.03165, 2139.101, 7822.355, 11400.98, 12447.22, 
    11229.59, 9500.495, 9160.496, 8573.722, 3866.707, 580.3088, 78.53415, 
    3.80173, 2004.922, 4006.043, 3283.891, 1372.212, 426.692, 80.53307, 
    21.18099, 6.336446, 0.9003974, 0.127025, 0.01270251, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0.05426566, 0.5426567, 129.477, 763.0168, 
    2064.251, 3071.403, 3156.496, 3241.59, 4342.653, 4860.217, 4586.532, 
    3734.051, 2769.331, 2437.281, 2885.591, 3333.9, 2597.936, 733.8609, 
    97.80436, 0.1915518, 0.05201121, 0.03122856, 122.9769, 245.9225, 
    154.2318, 21.57413, 2.421838, 0.2720145, 0.2930991, 0.3348363, 0.4183033, 
    0.4501407, 0.365643, 0.1425516, 0.02803748, 0, 0.2807808, 0.5615616, 
    0.3013227, 0.0410838, 0.07142995, 0.1017761, 0.05159655, 0.001416998, 
    0.001719869, 0.004273215, 0.01303107, 0.01656029, 0.008408367, 
    0.0002564475, 0.0006627321, 0.001069017, 0.0005345084, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4238.484, 15714.18, 23113.13, 
    25400.16, 12021.16, 1449.781, 1885.86, 3163.033, 3889.953, 4802.137, 
    7202.479, 8113.299, 5286.531, 842.3539, 84.22935, 0, 0.02695867, 
    0.05391733, 0.02695867, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 12.31137, 123.1137, 2871.398, 9353.699, 11812.82, 12295.94, 
    11150.76, 9516.146, 9184.122, 8599.535, 5021.76, 1158.312, 109.0841, 
    16.47654, 1992.565, 3968.653, 3579.226, 2310.689, 734.1765, 71.9956, 
    19.34044, 5.860137, 0.8327124, 0.1174754, 0.01174755, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01440574, 0.1440574, 35.6647, 232.3137, 
    616.6503, 1181.513, 1938.509, 2727.409, 3540.538, 4012.076, 3968.042, 
    3736.12, 2747.671, 2327.124, 2815.709, 3304.294, 1866.056, 146.5428, 
    14.70799, 0.04368644, 0.03027677, 0.02827959, 114.0034, 227.9785, 
    162.3127, 33.9598, 7.917964, 5.472927, 9.425361, 11.35953, 6.42819, 
    0.602105, 0.2582868, 0.140134, 0.02470286, 0, 0.2532881, 0.5065762, 
    0.376871, 0.2471659, 1.186429, 2.125692, 1.065098, 0.004503669, 
    0.007216135, 0.00995928, 0.009010181, 0.005856137, 0.001583, 
    5.381528e-05, 0.0001390738, 0.0002243322, 0.0001121661, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.371262, 33.71262, 4859.703, 17296.72, 
    23886.94, 26018.91, 10707.22, 1860.285, 2198.991, 3216.599, 4011.693, 
    5010.784, 7230.129, 8056.579, 6174.497, 1509.609, 158.7748, 7.459694e-07, 
    0.02493232, 0.0498639, 0.02493195, 0, 0, 0, 0, 0, 0, 0, 0.07724743, 
    0.1544949, 0.07724743,
  0, 0, 0, 67.72261, 677.2261, 5004.446, 10628.76, 11095.31, 11034.27, 
    10489.85, 9688.527, 9495.352, 9123.093, 6583.314, 2843.716, 753.333, 
    258.1969, 1335.112, 3535.766, 3411.818, 2985.559, 912.8926, 0.2369497, 
    0.8028175, 1.368685, 0.7157555, 0.02151565, 0.002151566, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003310521, 0.03310522, 7.838697, 
    77.69176, 912.3942, 2637.025, 3105.755, 3234.748, 2902.19, 2283.529, 
    1250.858, 874.0872, 1809.048, 2744.008, 1375.61, 2.468189, 0.2465518, 
    0.0001420851, 0.0005261838, 0.003105132, 26.51439, 54.39213, 53.74761, 
    51.70517, 48.22124, 46.90939, 71.20369, 95.49799, 48.83603, 0.7804139, 
    0.1680526, 0.04909702, 0.00636443, 0, 0.002959677, 0.0228318, 0.121636, 
    0.7977769, 10.6537, 19.0266, 9.538581, 0.02631116, 0.01810201, 0.0145201, 
    0.007311139, 0.002239376, 0.0002958344, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 82.09389, 820.939, 13907.36, 28097.25, 
    25787.46, 18303.41, 7655.936, 1948.218, 2312.226, 3213.627, 5045.565, 
    6795.439, 7430.12, 7629.989, 5506.786, 2470.066, 508.4637, 1.816516e-05, 
    0.004575375, 0.009132585, 0.004566292, 0, 0, 0, 0, 0, 0, 0, 0.7223098, 
    1.44462, 0.7223098,
  0, 0, 0, 66.08292, 660.8293, 5913.607, 11211.82, 11231.62, 11145.14, 
    10697.85, 10066.66, 9947.589, 9747.59, 8039.352, 5008.458, 2030.369, 
    1071.43, 1268.756, 1872.1, 2516.031, 2734.463, 1367.257, 0.05083049, 
    0.1721252, 0.29342, 0.1534438, 0.004612221, 0.0004612223, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 1.505038e-05, 4.58055e-05, 4.58055e-05, 4.58055e-05, 
    1.505038e-05, 0, 0, 0, 0.0007096628, 0.007096628, 1.680946, 16.66043, 
    498.1435, 1659.696, 2120.408, 2238.921, 1948.524, 1425.206, 615.375, 
    324.6988, 948.0128, 1571.327, 787.0386, 0.9635047, 0.1450839, 0.03019465, 
    0.01009072, 0.007096521, 7.938109, 29.97642, 45.88233, 50.68905, 
    46.26095, 42.90881, 65.469, 88.02921, 46.73733, 3.17178, 2.52306, 
    2.187362, 0.5993734, 9.600552e-06, 0.0006474314, 0.00493001, 0.08328172, 
    0.7425233, 9.781483, 17.40531, 8.727777, 0.025501, 0.01725241, 
    0.01365307, 0.004612495, 0.0006102445, 6.102447e-05, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.1836735, 1.836735, 439.136, 
    4352.789, 19949.68, 27193.45, 22052.49, 8920.01, 4352.97, 2800.102, 
    2983.538, 3442.551, 5093.219, 6717.39, 7153.562, 7278.383, 5621.601, 
    3086.687, 732.6945, 0.136214, 0.01683328, 0.001529464, 0.0001529465, 0, 
    0, 0, 0, 0, 0, 0, 0.6750964, 1.350193, 0.6750964,
  0, 0, 0, 30.36419, 303.6419, 4992.846, 11697.53, 12385.61, 12484.25, 
    12204.81, 11663.17, 11160.52, 10374.14, 9150.112, 7459.201, 4687.038, 
    2044.629, 552.8563, 241.2604, 1076.005, 1910.75, 955.3751, 4.136906e-05, 
    3.249723e-05, 2.799451e-05, 7.634227e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0.000176085, 0.0005359109, 0.0005359109, 0.0005359109, 0.000176085, 0, 
    0, 0, 0, 0, 0.0007601002, 0.007601003, 18.41974, 184.0378, 739.8884, 
    1229.256, 1180.844, 1001.692, 413.9426, 170.2719, 177.8063, 185.3407, 
    93.01933, 0.6979322, 0.9717527, 1.245573, 0.6755413, 0.1055093, 6.9332, 
    23.03252, 27.56659, 28.97515, 9.561351, 0.06097843, 0.3644165, 3.565483, 
    14.35878, 23.39712, 24.78287, 25.46469, 8.367282, 0.0002282386, 
    7.442775e-05, 5.151975e-05, 0.06898512, 0.1379187, 0.09818599, 
    0.02879044, 0.01855201, 0.01423064, 0.006178587, 0.001450879, 
    0.0002178425, 3.4645e-05, 3.464501e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 5.434189, 54.34189, 7888.495, 23719.22, 23648.46, 
    23559.2, 9216.556, 2197.815, 2602.103, 3585.305, 3747.348, 3858.869, 
    4048.121, 4470.917, 6195.183, 6885.095, 5993.554, 3353.053, 837.5305, 
    4.01944, 0.4019442, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.09833256, 0.1966651, 
    0.09833256,
  0, 0, 0, 9.472984, 94.72985, 4516.695, 11549.5, 12401.73, 12428.21, 
    12089.82, 11604.74, 11475.69, 11266.99, 10623.65, 9075.3, 5431.97, 
    1871.257, 308.7734, 57.20512, 505.2044, 953.2036, 476.6019, 0.0001367601, 
    0.000106123, 9.084192e-05, 2.465404e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.0002320404, 0.0004640808, 0.0004628713, 0.0004603998, 0.005017656, 
    0.04603549, 0.7303674, 6.342423, 27.6378, 36.86161, 36.13512, 35.40864, 
    97.7336, 269.9872, 375.2892, 434.3886, 450.472, 463.3162, 209.7334, 
    85.63971, 138.8353, 192.0309, 159.7993, 72.38734, 17.64039, 2.16099, 
    8.463503, 15.7628, 17.02695, 17.29432, 14.79291, 10.1878, 2.720242, 
    0.01518856, 0.1261912, 0.8714947, 8.581206, 22.4222, 23.45742, 23.83382, 
    7.83244, 0.000923419, 0.0002435896, 0.0001423384, 0.015385, 0.03062766, 
    0.02286101, 0.005609354, 0.003930971, 0.004262418, 0.3295383, 0.6548142, 
    0.334991, 0.005194465, 0.0005194467, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 33.88317, 338.8318, 11215.82, 21442.25, 19539.92, 
    13234.2, 4790.29, 1776.088, 2304.148, 3561.246, 3853.606, 3886.826, 
    3664.127, 3555.147, 4755.882, 6483.91, 5895.738, 3985.09, 1202.062, 
    70.25812, 7.025815, 0, 0, 0, 0, 0, 0.01580007, 0.03160014, 0.01580007, 0, 
    0.02152425, 0.0430485, 0.02152425,
  0, 0, 0, 1.161202, 11.61202, 2060.896, 7475.961, 10487.62, 11270.52, 
    11156.29, 11100.4, 11450.01, 12164.44, 11876.53, 10023.27, 4834.873, 
    1041.42, 110.0326, 5.411008, 5.179039, 4.94707, 1.682338, 0.003409128, 
    0.001600005, 0.0009329494, 0.0001710839, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.513629e-05, 5.027259e-05, 4.409142e-05, 3.146034e-05, 0.1759722, 
    1.759452, 60.39362, 244.41, 488.6774, 575.5962, 564.181, 552.7657, 
    612.2043, 671.6429, 372.0819, 33.64098, 11.50811, 4.927188, 11.09012, 
    41.21917, 164.8446, 405.3693, 967.9014, 1182.253, 594.0665, 5.880546, 
    115.9169, 225.9533, 129.9892, 11.77356, 1.497679, 0.1538868, 0.01752254, 
    0.002371602, 0.002377336, 0.002380142, 0.002032127, 0.001102619, 
    0.0005415835, 0.0003656891, 0.001456566, 0.002222702, 0.002036332, 
    0.001463721, 0.0009755949, 0.0005310506, 0.000295551, 0.0001540272, 
    3.009161e-05, 0, 5.098974, 10.19795, 5.216659, 0.08060553, 0.008060556, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 706.9301, 
    3924.714, 11060.33, 13804.53, 9150.005, 2285.323, 1686.736, 1598.032, 
    1792.606, 2209.976, 3102.02, 3441.118, 3244.567, 3048.016, 3747.704, 
    5177.501, 5094.348, 4700.992, 2964.582, 923.1309, 115.8131, 0, 0, 0, 0, 
    0, 0.246719, 0.4934381, 0.246719, 0, 0, 0, 0,
  0, 0, 0, 1.248457, 12.48457, 1623.141, 5934.384, 8540.462, 9403.34, 
    9429.018, 9454.695, 10475.89, 12236.68, 12099.37, 10891.95, 5238.875, 
    1042.449, 105.6806, 1.319386, 1.26298, 1.206573, 0.4955856, 0.05927191, 
    0.007506582, 0.0007050447, 5.952726e-05, 0, 3.506618e-05, 0.0001067232, 
    0.0001058979, 0.0001032386, 3.350732e-05, 0, 0, 0, 0, 0, 8.775258e-07, 
    8.775259e-06, 0.08576591, 0.8574749, 5.706918, 39.06234, 256.409, 
    507.3945, 550.2444, 554.0464, 545.5942, 541.4581, 594.1406, 646.8231, 
    331.8285, 16.83394, 15.3173, 19.73895, 58.80688, 212.9159, 870.5289, 
    1556.485, 1496.583, 1262.311, 395.2635, 29.582, 123.4484, 217.3147, 
    120.6063, 8.211332, 0.8919386, 0.03459873, 0.004959708, 0.001518488, 
    0.001459836, 0.001420882, 0.001346887, 0.001202703, 0.0006670093, 
    0.0004542583, 0.00129108, 0.002127902, 0.001936289, 0.001385043, 
    0.001045007, 0.0007123183, 0.000230237, 2.954654e-05, 3.830107e-06, 0, 
    4.894164, 9.788328, 5.006829, 0.07716764, 0.007716767, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001111064, 0.01111064, 1935.019, 
    6636.153, 8136.715, 8549.833, 3970.888, 1471.349, 1372.866, 1354.094, 
    1341.839, 1354.135, 2214.356, 2821.573, 2732.512, 2643.451, 2944.271, 
    3771.265, 4342.072, 4516.075, 3422.217, 889.4426, 99.89934, 0.0001035901, 
    1.035901e-05, 0, 0, 0, 0.237411, 0.474822, 0.237411, 0, 0, 0, 0,
  0, 0, 0, 6.023789, 60.23789, 1739.932, 5642.067, 6667.79, 6934.281, 
    6964.165, 6994.048, 8338.429, 10830.93, 11313.28, 11614.13, 5910.865, 
    1147.477, 114.8951, 0.1467319, 0.1325049, 0.130386, 0.7638891, 1.397392, 
    0.6993124, 0.0004966999, 6.438704e-05, 0, 0.0008221695, 0.002502255, 
    0.002482905, 0.002420556, 0.0007856201, 0, 0, 0, 0, 0, 0, 0, 4.778419, 
    47.78419, 429.8328, 1042.673, 971.6058, 748.7113, 243.5371, 45.03667, 
    166.3409, 287.6451, 228.8783, 78.57059, 21.09451, 10.60009, 69.2571, 
    675.9595, 2772.986, 5160.851, 6688.924, 7204.053, 3642.017, 911.0739, 
    521.6149, 364.0405, 102.0092, 10.89353, 1.095856, 0.002460042, 
    9.748816e-05, 0, 0.0006600723, 0.001320145, 0.001234693, 0.001149241, 
    0.001179363, 0.001240917, 0.001157486, 0.0008346804, 0.0002287629, 0, 
    1.106997e-06, 8.539688e-06, 0.001880983, 0.003740775, 0.001870387, 0, 0, 
    0, 0.1768553, 0.3537107, 0.1768553, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.02605026, 0.2605027, 3370.67, 6740.579, 6000.279, 
    3840.464, 2109.495, 1121.218, 895.3005, 841.9442, 805.2676, 770.867, 
    1352.691, 2123.948, 2340.076, 2431.492, 2478.649, 2535.088, 3393.956, 
    4023.987, 3088.425, 764.0002, 81.67622, 0.002428797, 0.0002428798, 0, 0, 
    0, 0.01696275, 0.03392551, 0.01696275, 0, 0, 0, 0,
  0, 1.039572e-06, 1.039572e-05, 22.28661, 222.8659, 2679.783, 4943.816, 
    4983.789, 5023.762, 5272.995, 6044.885, 8358.192, 10796.25, 12222.5, 
    12737.24, 7207.227, 1496.156, 149.8456, 0.1405272, 0.04408801, 
    0.02972473, 0.6995277, 1.369331, 0.6849535, 0.0002322409, 3.01053e-05, 0, 
    0.0008102039, 0.002465838, 0.002446901, 0.00238588, 0.0007744331, 0, 0, 
    0, 0, 0, 0.0002938204, 0.002938204, 31.66541, 221.6443, 675.4391, 
    1009.356, 953.8544, 747.7804, 245.8073, 48.51712, 194.4846, 340.4522, 
    265.7552, 82.77396, 33.37426, 28.13963, 332.4996, 1547.121, 3298.981, 
    5052.399, 6442.534, 6916.958, 3449.372, 670.5591, 461.1085, 368.3316, 
    99.12075, 2.484059, 0.2547401, 0.002522659, 0.0002958827, 0.0002071174, 
    0.0008417356, 0.001476354, 0.001117038, 0.0007577221, 0.0008942509, 
    0.001253623, 0.001454463, 0.00151854, 0.0006760532, 0, 1.27721e-06, 
    9.852764e-06, 0.001843624, 0.003662799, 0.0018314, 0, 0, 0, 0.0403183, 
    0.0806366, 0.0403183, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.02324555, 0.2324555, 1.28949, 1.90021, 1.113478, 0.3267456, 3369.819, 
    6739.312, 5977.694, 3757.882, 2080.636, 910.0921, 648.5076, 598.488, 
    616.9998, 699.8896, 1098.348, 1563.568, 1778.039, 1825.777, 1573.817, 
    1450.517, 2016.183, 2581.849, 1951.958, 452.7647, 45.28157, 0.00241942, 
    0.0002419421, 0, 0, 0, 0.003867056, 0.007734111, 0.003867056, 0, 0, 0, 0,
  0, 0.0001122792, 0.001122792, 150.0965, 1061.219, 3618.209, 4624.152, 
    4392.118, 3917.961, 4099.748, 5583.665, 10234.49, 14042.09, 14519.8, 
    14749.41, 9068.712, 2313.584, 233.6246, 1.055787, 0.1001325, 
    2.496587e-07, 0.02420647, 0.0484127, 0.02420635, 0, 0, 0, 0.0002604925, 
    0.0007928032, 0.0007928032, 0.0007928032, 0.0002604925, 0, 0, 0, 0, 0, 
    0.03173414, 0.3173414, 511.1442, 1021.362, 882.6575, 666.2275, 654.8926, 
    643.5576, 493.3875, 420.9432, 1593.704, 2766.464, 1957.906, 305.6334, 
    432.9385, 758.5954, 1509.482, 2329.285, 2778.57, 2943.356, 1178.309, 
    151.762, 79.99258, 56.52216, 44.58367, 37.33905, 10.2973, 0.0002115027, 
    0.001108008, 0.004066994, 0.007668766, 0.0100912, 0.01004725, 
    0.009334846, 0.003213911, 0.0002470525, 0.0004428438, 0.001076091, 
    0.002059528, 0.002422856, 0.001211428, 0, 8.910154e-05, 0.0001782031, 
    0.0001524435, 7.891689e-05, 1.879116e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.091171, 10.91171, 60.53003, 89.19787, 
    44.60469, 0.01151132, 3301.861, 6603.71, 5880.415, 3746.525, 2062.146, 
    857.5699, 581.14, 526.6676, 557.4343, 670.9172, 1120.427, 1305.641, 
    874.8467, 444.0523, 454.883, 477.0153, 455.8772, 352.8219, 99.97276, 
    0.5942796, 0.06269126, 0.001553941, 0.0001553942, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0,
  1.098693e-16, 0.0004779609, 0.004779609, 357.1668, 1666.482, 3825.272, 
    4624.152, 4392.118, 3917.961, 3987.533, 5097.925, 9898.258, 14107.42, 
    14512.33, 14669.13, 9614.183, 2823.646, 333.8418, 4.168117, 0.4155457, 
    2.496587e-07, 0.005628719, 0.01125719, 0.005628594, 0, 0, 0, 
    0.0002604925, 0.0007928032, 0.0007928032, 0.0007928032, 0.0002604925, 0, 
    0, 0, 0, 0, 0.135089, 1.35089, 745.8241, 1487.704, 1095.895, 295.2415, 
    353.5132, 519.5518, 980.6733, 1630.155, 2477.184, 2766.464, 1957.906, 
    305.6334, 418.7136, 730.1456, 1800.938, 2258.263, 1950.088, 1059.88, 
    309.0423, 35.28854, 18.60032, 13.14285, 10.36682, 8.682262, 2.394507, 
    0.0002875969, 0.00151004, 0.005130948, 0.008158744, 0.0100072, 
    0.01000526, 0.009334846, 0.003122899, 0.0003077274, 0.0003916338, 
    0.000837721, 0.00197798, 0.002422856, 0.001211428, 0, 0.0003628144, 
    0.0007256287, 0.0004546632, 6.291015e-05, 6.291018e-06, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.091171, 10.91171, 
    60.53003, 89.19787, 44.60028, 0.002693755, 3078.973, 6157.943, 5580.915, 
    3788.315, 2107.419, 850.6048, 577.6575, 526.6676, 557.4343, 670.9172, 
    1120.427, 1305.641, 1025.927, 333.4483, 155.1828, 102.7072, 92.15623, 
    84.06805, 24.2598, 0.1382636, 0.01540903, 0.0007536496, 7.536499e-05, 0, 
    0, 0, 0, 0, 1.152623e-16, 4.180794e-16, 5.855295e-16, 6.390876e-16, 
    3.866083e-16,
  0.05682618, 0.2754517, 2.417938, 454.9314, 1939.702, 3923.815, 4631.608, 
    4407.889, 3950.725, 3966.716, 4577.531, 7898.516, 11299.98, 12110.85, 
    12362.41, 8508.242, 3226.696, 1089.518, 284.5408, 33.58276, 2.442224, 
    0.2442225, 0, 0, 0, 0, 0, 0.0004599103, 0.001399727, 0.001323895, 
    0.001079548, 0.0003166726, 0, 0, 0, 0, 0, 26.91273, 269.1274, 1222.167, 
    1658.482, 880.9385, 103.3953, 150.2549, 464.8838, 2540.981, 4081.541, 
    2541.092, 663.7968, 571.466, 517.3333, 310.9243, 116.3975, 18.36589, 
    8.024241e-06, 8.024244e-07, 1.705142e-15, 4.215774e-16, 2.304081e-16, 
    2.117133e-07, 9.368882e-07, 1.334104e-06, 2.311174e-06, 8.121775e-05, 
    0.0007738663, 0.004258594, 0.006262574, 0.006073905, 0.005885235, 
    0.00708227, 0.008279306, 0.004389601, 0.0004998961, 0.0005782279, 
    0.0006565595, 0.0003282798, 0, 0, 0, 0.007565229, 0.01785835, 0.01629091, 
    0.01127916, 0.003067643, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1.250649, 4.791867, 7.580484, 8.43978, 4.219902, 
    2.225373e-05, 958.5879, 3720.193, 6074.091, 6820.671, 4061.626, 1302.581, 
    1625.553, 1948.525, 1757.375, 1566.226, 2055.224, 2544.223, 1702.908, 
    295.0663, 29.50664, 1.054233e-14, 1.054234e-15, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.05961554, 0.2162374, 0.3028453, 0.3305465, 0.1999601,
  0.2443869, 1.183256, 10.38507, 823.4487, 2975.459, 4320.497, 4707.417, 
    4383.14, 4058.863, 4157.164, 4787.176, 6612.297, 8642.739, 9955.06, 
    10388.85, 7829.682, 4193.498, 2519.233, 1362.418, 300.1956, 10.50304, 
    1.050304, 0, 0, 0, 0, 0, 0.0005682491, 0.001837062, 0.002064198, 
    0.002134688, 0.0007013976, 0, 0, 0, 0, 0, 97.07401, 507.012, 1340.935, 
    1658.482, 880.9385, 103.3953, 134.6479, 344.4873, 2391.601, 4081.541, 
    2391.92, 563.9221, 543.7419, 523.5618, 241.4428, 33.45951, 3.345969, 
    8.024241e-06, 8.024244e-07, 1.705142e-15, 4.215774e-16, 2.304081e-16, 
    2.117133e-07, 9.368882e-07, 1.334104e-06, 2.311174e-06, 0.0005493574, 
    0.002970647, 0.008204003, 0.01021081, 0.008048023, 0.005885235, 
    0.006465943, 0.00704665, 0.00386533, 0.0004593176, 0.0004125743, 
    0.0003782416, 0.0001078552, 0, 0, 0, 0.007565229, 0.01785835, 0.01629091, 
    0.01127916, 0.003067643, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.2937936, 1.125671, 1.780754, 1.982613, 0.9913178, 
    2.225373e-05, 132.2052, 1324.283, 6542.783, 9215.358, 5638.895, 2062.431, 
    3256.312, 4450.192, 3596.948, 2608.844, 2589.177, 2569.51, 1591.359, 
    256.188, 25.61881, 2.47653e-15, 2.476531e-16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.2563829, 0.9299515, 1.302418, 1.421549, 0.859949,
  433.5799, 287.5729, 242.8749, 1798.959, 5762.982, 7323.586, 7683.497, 
    5933.87, 5077.669, 5356.498, 6060.82, 6158.597, 6303.648, 7312.701, 
    8593.473, 9701.489, 10049.72, 7830.657, 2647.897, 680.7717, 125.6614, 
    12.56614, 0, 0, 0, 0, 0, 0.0001556969, 0.001556969, 0.02254836, 
    0.1927873, 167.8751, 335.1908, 174.8411, 6.531004, 1.854278, 1.157745, 
    152.9732, 631.6837, 1193.479, 1388.5, 1085.411, 316.5646, 49.2141, 
    6.903552, 993.9738, 1981.044, 1266.82, 552.5959, 570.2963, 587.9966, 
    313.5601, 13.68165, 2.121825, 0.3588678, 0.03588376, 1.480518e-06, 
    5.730036e-06, 3.426252e-05, 0.005026196, 0.04964763, 0.4542696, 1.242618, 
    1.505156, 1.570019, 1.029173, 0.3047601, 0.04544552, 0.00668003, 
    0.004026433, 0.002930236, 0.0007008254, 8.939771e-06, 5.227228e-06, 
    3.710989e-06, 8.487354e-07, 0, 2.05403e-05, 0.0002094468, 0.00407194, 
    0.00752631, 0.004026904, 0.0001806499, 1.8065e-05, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002974264, 0.01093055, 
    0.01272551, 0.01629124, 0.1947804, 1.723811, 23.62141, 200.2262, 
    5784.859, 10989.02, 7110.499, 3231.975, 5687.476, 8142.976, 6997.478, 
    3813.484, 1898.418, 585.3557, 166.7096, 48.21508, 4.82151, 2.292973e-17, 
    2.292974e-18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.09116257, 0.9116257, 96.83486, 
    370.8208, 611.7827, 688.9551, 622.1331,
  1092.358, 956.3947, 892.7322, 2532.357, 5731.584, 7321.451, 7747.953, 
    5967.929, 5096.854, 5554.03, 6011.207, 5606.674, 4780.019, 5614.333, 
    8380.578, 12411.32, 13877.85, 11278.29, 4519.609, 1864.108, 527.9578, 
    56.28817, 0, 0, 0, 0, 0, 0.0001559423, 0.001559423, 0.08725146, 
    0.8397668, 250.3151, 498.1816, 256.4548, 6.684432, 1.958864, 1.255056, 
    188.2258, 674.5204, 913.22, 980.5113, 732.075, 365.9533, 82.65025, 
    1.236456, 294.5695, 587.9026, 525.605, 463.3073, 628.5063, 793.7054, 
    407.5139, 7.591561, 1.529272, 0.3666435, 0.03665103, 6.494258e-06, 
    2.513468e-05, 0.0001502918, 0.005344455, 0.05074981, 0.4640736, 1.269685, 
    1.537849, 1.604106, 1.05126, 0.3109345, 0.0478405, 0.006323615, 
    0.001720604, 0.0005182105, 5.182107e-05, 0, 0, 0, 0, 0, 2.150387e-05, 
    0.0002150387, 0.001219289, 0.001810665, 0.0009053326, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.7546014, 
    7.546014, 34.79845, 189.5182, 5772.07, 11008.13, 7503.61, 3999.087, 
    6091.099, 8183.111, 7089.135, 3909.914, 1187.039, 129.0111, 35.34014, 
    10.68525, 1.068526, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.3998826, 3.998827, 
    557.7264, 1741.612, 1825.131, 1811.988, 1481.094,
  2052.988, 2264.309, 2991.278, 4066.584, 4899.867, 5024.401, 5034.279, 
    4602.175, 4390.721, 5123.589, 5856.458, 4997.251, 4138.045, 5971.476, 
    11084.1, 14826.67, 15954.62, 13263.24, 6657.731, 4879.024, 3741.198, 
    978.3235, 0.7253442, 0.07253445, 0, 0, 0, 3.984437e-05, 0.0003984437, 
    36.23237, 181.7545, 458.8062, 563.4329, 283.5041, 2.204198, 1.398648, 
    1.278672, 5.517494, 44.90092, 218.133, 305.7841, 267.7436, 157.1257, 
    70.9397, 19.54088, 28.08874, 55.52504, 85.80258, 181.2357, 774.6373, 
    1127.24, 571.9708, 5.994349, 1.293652, 0.3524861, 0.1024577, 0.03290403, 
    0.004716088, 0.00158576, 0.001715183, 0.002584164, 0.0185087, 0.05424368, 
    0.06567563, 0.06844267, 0.045229, 0.01444663, 0.005176244, 0.002239603, 
    0.0003630118, 9.29886e-06, 9.298865e-07, 0, 0, 0, 0, 0, 2.102817e-06, 
    1.074111e-05, 2.770026e-05, 3.412992e-05, 1.706496e-05, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002467534, 0.0004935067, 
    0.0002467534, 0, 0, 0, 0, 0, 0.01466242, 0.1466242, 414.4285, 828.429, 
    808.7675, 789.106, 1818.981, 4106.504, 4386.21, 4399.53, 3635.737, 
    2412.091, 1400.482, 547.1523, 88.60174, 2.32561, 0.635211, 0.1917381, 
    0.01917381, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0007440313, 0.007440314, 
    49.1109, 490.9528, 2821.446, 4209.326, 3981.679, 3263.404, 2527.968,
  2461.868, 2615.271, 3125.942, 3954.849, 4262.95, 3986.384, 3421.226, 
    3624.99, 4300.723, 5428.206, 5849.563, 4987.592, 4125.621, 6002.895, 
    11207.18, 14927.67, 16054.05, 13216.33, 6699.755, 4968.846, 3864.852, 
    1022.964, 3.246426, 0.3246428, 0, 0, 0, 3.46721e-05, 0.000346721, 
    316.4676, 963.1602, 941.0663, 869.9305, 275.1244, 0.5354841, 0.6241555, 
    1.21952, 4.217129, 24.81127, 180.8378, 291.7141, 238.4115, 140.2301, 
    133.6852, 127.1404, 46.87969, 11.49771, 14.91398, 142.9143, 836.8972, 
    1134.624, 572.2703, 3.613558, 0.902364, 0.280737, 0.09148554, 0.03701646, 
    0.01387003, 0.005972529, 0.0009493274, 0, 0, 0, 6.978983e-06, 
    6.978984e-05, 0.0003252165, 0.0006903397, 0.0009001797, 0.0009717774, 
    0.0003380678, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0002577465, 0.0005154929, 0.0002577465, 0, 
    0, 0, 0, 0, 0.06562467, 0.6562467, 835.3454, 1668.775, 1361.425, 
    733.3619, 658.5173, 626.3414, 2990.298, 4289.711, 2673.341, 444.7771, 
    221.0151, 134.159, 25.10958, 0.002673772, 0.0002673773, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0.003330064, 0.03330065, 51.32304, 512.5311, 2886.618, 
    4276.722, 4010.524, 3260.345, 2750.486,
  2594.078, 2726.095, 3161.236, 3776.569, 3999.115, 3660.263, 2967.825, 
    3311.389, 4577.306, 6954.816, 7855.193, 6565.634, 5126.263, 5789.71, 
    7985.026, 11027.42, 12122.37, 10432.76, 5796.287, 3294.123, 1378.205, 
    245.9346, 12.56301, 1.256301, 0, 0, 0, 0.001984232, 0.01984232, 967.8972, 
    2702.708, 2484.529, 1815.439, 505.4523, 0.02480829, 0.151334, 2.73372, 
    11.3533, 43.42969, 288.2057, 846.2703, 1401.405, 1751.174, 1701.072, 
    1422.215, 415.8674, 0.3002812, 98.23308, 308.3573, 329.4708, 336.0264, 
    110.5801, 0.1040473, 0.03490198, 0.01487297, 0.004373182, 0.002787965, 
    1.133455, 2.264122, 1.132061, 0, 0, 0, 3.513149e-05, 0.000163801, 
    0.0003408819, 0.00047816, 0.0005222964, 0.0005440575, 0.0001787618, 0, 0, 
    0, 0, 0, 2.834295e-05, 5.668591e-05, 2.834295e-05, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1.650628e-05, 3.301255e-05, 
    1.650628e-05, 0, 0.2853062, 2.8531, 15.28999, 92.98447, 1364.58, 
    3648.308, 3397.121, 2607.161, 787.4029, 50.64072, 37.1208, 35.10719, 
    166.4949, 297.8827, 157.2079, 16.53311, 25.69385, 34.85459, 17.4274, 
    6.980677e-05, 6.980681e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13.90419, 
    27.80837, 20.41499, 5.30679, 46.71128, 434.7813, 2177.342, 3361.273, 
    3304.844, 3139.021, 2777.711,
  2798.481, 2883.996, 3197.939, 3773.546, 3990.698, 3650.659, 2955.796, 
    3302.555, 4594.524, 7057.85, 7992.424, 7001.383, 4976.213, 5180.815, 
    5795.797, 7006.875, 7901.461, 7556.407, 6128.653, 3555.135, 1137.56, 
    239.5013, 45.98085, 4.598087, 0, 0, 0, 0.008941149, 0.0894115, 1874.706, 
    3749.152, 3372.39, 2143.157, 560.535, 0.01111815, 0.4614481, 3.485093, 
    17.23444, 108.5548, 658.7348, 1653.479, 2143.359, 2364.692, 2054.696, 
    1458.887, 393.7933, 5.240454e-05, 272.4314, 544.8627, 449.6443, 193.1852, 
    40.99731, 0, 0, 0, 0, 0, 1.209144, 2.418288, 1.209144, 0, 0, 0, 
    5.176115e-05, 0.0001868449, 0.0002444817, 0.0002691143, 0.0002662182, 
    0.0002448017, 7.520948e-05, 0, 0, 0, 0, 0, 0.0001294835, 0.000258967, 
    0.0001294835, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1.30343, 13.0343, 69.85155, 424.7953, 2017.401, 3833.937, 
    3544.717, 2623.077, 733.4944, 1.51457, 4.124999, 12.2731, 21.55268, 
    24.75148, 13.59293, 2.434386, 7.969119, 13.50385, 6.751925, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 15.67906, 31.35813, 22.86519, 5.510051, 42.6819, 
    394.9529, 1567.503, 2716.748, 3006.052, 3032.186, 2915.333,
  3146.159, 3337.506, 3669.111, 4624.111, 4995.323, 4349.717, 3030.436, 
    3317.411, 4337.346, 6442.463, 7253.312, 5973.439, 4693.566, 4907.979, 
    5122.393, 4236.249, 3350.106, 6712.072, 10074.04, 8927.722, 5602.771, 
    3276.257, 1315.809, 211.5402, 1.681701, 0.2179983, 0, 0.8691179, 
    10.93345, 2208.151, 4381.058, 3823.941, 2189.175, 767.2085, 136.3578, 
    18.35259, 0.7773394, 15.65745, 301.9497, 1483.923, 2497.566, 2569.964, 
    2581.36, 1719.931, 552.0558, 75.96044, 3.614852e-05, 568.2218, 1136.444, 
    786.5593, 149.5462, 14.95463, 0, 0, 0, 0, 0, 0.7693192, 1.538638, 
    0.7693192, 0, 0, 0, 1.53461e-06, 1.250261e-05, 4.13626e-05, 6.277838e-05, 
    6.335993e-05, 6.261342e-05, 2.027322e-05, 0, 0, 0, 0, 0, 0.0008889613, 
    0.001777923, 0.0008889613, 0, 0.002112539, 0.02312556, 9.889574, 
    19.70866, 9.854331, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.741549e-05, 
    0.0003551768, 0.0007484138, 0.001996229, 12.15271, 121.4894, 1389.047, 
    4024.524, 4789.604, 5004.968, 4495.55, 3466.814, 1960.181, 622.1638, 
    103.6114, 23.43749, 127.4412, 300.5322, 517.8714, 592.1988, 350.2883, 
    41.85721, 15.27838, 7.027122, 1.109856, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15.94776, 31.89551, 17.95914, 4.022761, 50.86862, 406.242, 1410.291, 
    2474.385, 2847.961, 3003.055, 3074.607,
  3505.861, 3990.457, 4555.207, 5497.607, 5832.835, 5089.543, 3570.642, 
    3728.667, 4317.05, 5942.38, 6593.081, 5325.458, 4057.836, 4271.623, 
    4485.409, 3818.49, 3151.572, 6805.579, 10459.59, 9339.036, 6031.552, 
    3556.465, 1429.988, 242.4903, 7.845005, 1.016945, 0, 3.929802, 49.75803, 
    2283.326, 4405.877, 3904.25, 2466.02, 1519.734, 715.46, 138.1839, 
    0.4641456, 243.093, 1284.783, 3269.954, 4390.773, 4032.827, 2920.009, 
    1620.176, 486.7438, 59.53434, 3.557985e-05, 584.5016, 1169.003, 761.7992, 
    121.4367, 12.14368, 0, 0, 0, 0, 0, 0.3460784, 0.6921567, 0.3460784, 0, 0, 
    0, 0, 0, 1.890259e-05, 5.752961e-05, 5.752961e-05, 5.752961e-05, 
    1.890259e-05, 0, 0, 0, 0, 0, 0.0009511314, 0.001902263, 0.0009511314, 0, 
    0.01075365, 0.1096766, 46.1314, 91.93938, 45.96969, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0.0002678388, 0.001656872, 0.003491293, 0.009312252, 
    56.69144, 566.7386, 5288.846, 8922.837, 7880.361, 5080.077, 3889.328, 
    2835.458, 925.0995, 165.276, 94.812, 77.76153, 177.2869, 345.8204, 
    568.2263, 645.2327, 385.033, 44.79547, 9.920557, 2.590956, 0.2590958, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15.95716, 31.91431, 17.7955, 3.676692, 
    49.49994, 403.7562, 1420.926, 2476.554, 2770.962, 2925.775, 3184.91,
  3947.784, 4884.947, 5714.624, 5946.043, 6081.72, 6443.153, 6800.868, 
    7120.741, 7298.335, 7118.652, 6408.584, 4259.421, 3410.694, 3704.322, 
    4270.735, 4310.516, 4350.297, 6654.436, 8685.79, 7047.512, 2938.849, 
    1922.171, 1432.307, 688.8167, 206.5414, 26.8974, 0.005406982, 21.45749, 
    165.4929, 1480.435, 3809.862, 3889.945, 3853.97, 3316.75, 2345.299, 
    974.0905, 195.2926, 893.5055, 3187.724, 6484.02, 7680.708, 6571.05, 
    3501.942, 1698.422, 491.8102, 85.31981, 37.34111, 171.9266, 306.5121, 
    187.0593, 23.15291, 2.315336, 2.833646e-05, 1.145432e-05, 8.939953e-06, 
    2.041203e-05, 0.0001495228, 0.04917838, 0.09789905, 0.04894952, 0, 
    4.129842e-06, 8.259684e-06, 4.129842e-06, 0, 0.0001463, 0.0004452608, 
    0.0004452608, 0.0004452608, 0.0001463, 0, 0, 0, 0, 0, 5.333416e-05, 
    0.0002138448, 0.000276295, 0.0004214681, 3.464522, 34.63869, 308.8356, 
    516.5272, 258.2636, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0005692889, 
    0.005692889, 0.2791401, 2.67185, 660.1484, 3934.786, 11907.54, 15003.42, 
    9489.372, 1625.082, 719.6503, 410.5088, 128.1859, 32.98808, 75.37637, 
    155.9979, 256.6574, 358.5266, 454.1994, 485.5933, 228.0917, 4.752932, 
    0.6611149, 0.08848646, 0.008848649, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.8572941, 3.557971, 4.766434, 7.649235, 447.6915, 1666.499, 2601.683, 
    2886.63, 2868.341, 2830.967, 3089.899,
  3824.517, 6056.245, 6929.729, 6923.127, 6909.637, 6932.657, 7066.99, 
    7439.724, 7586.3, 7135.491, 5671.63, 4053.458, 2989.572, 3128.725, 
    3614.048, 4648.153, 5927.678, 7402.206, 7884.749, 5437.397, 1866.032, 
    1496.164, 1322.628, 975.0575, 642.9659, 163.498, 0.02576605, 39.43296, 
    304.0241, 1615.611, 3649.179, 3948.31, 3965.906, 3390.174, 2427.249, 
    1357.411, 674.766, 1512.129, 4432.316, 9131.325, 10868.57, 9672.528, 
    6018.072, 2450.947, 575.8416, 213.7027, 175.5721, 194.1405, 203.2271, 
    123.0067, 14.65291, 1.4655, 0.0001350325, 5.458358e-05, 4.260182e-05, 
    9.727004e-05, 0.0007125252, 0.02715832, 0.05213546, 0.02606773, 0, 
    1.968006e-05, 3.936011e-05, 1.968006e-05, 0, 0.000161556, 0.0004916923, 
    0.0004916923, 0.0004916923, 0.000161556, 0, 0, 0, 0, 0, 2.807546e-08, 
    2.807546e-07, 0.0001838639, 0.001832743, 3.880234, 38.76386, 336.1305, 
    559.0748, 279.5374, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002146335, 
    0.02146335, 1.314533, 12.6946, 2649.912, 9743.349, 14349.52, 15772.11, 
    7523.326, 363.558, 117.5224, 50.08189, 23.48017, 14.5996, 65.53082, 
    158.0488, 284.4148, 369.1941, 349.0884, 268.4232, 75.42133, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.7542988, 7.542989, 480.9414, 
    1797.065, 2875.578, 3212.36, 3074.78, 2793.638, 2963.149,
  3063.713, 5375.327, 9158.326, 8986.179, 8785.229, 7563.489, 5949.667, 
    5486.23, 5275.521, 5135.257, 4925.098, 4002.273, 3007.864, 2378.491, 
    2158.417, 4473.621, 7800.61, 8108.284, 8215.079, 4205.859, 1623.052, 
    1379.341, 1273.869, 1159.398, 1036.204, 684.741, 433.8009, 381.0916, 
    354.3652, 2073.335, 3533.555, 3419.242, 3101.428, 2741.221, 2300.544, 
    1641.865, 1209.594, 1892.07, 4773.977, 9988.919, 13718.79, 13730.87, 
    13390.88, 6769.938, 3163.886, 3062.229, 2960.573, 2475.89, 1821.852, 
    678.1819, 99.48269, 10.83673, 0.3917537, 0.03695294, 0.006634294, 
    0.0408071, 0.08095843, 0.07350925, 0.0491767, 0.01316409, 0, 
    8.925902e-05, 0.000178518, 8.925902e-05, 0, 2.075344e-05, 6.316265e-05, 
    6.316265e-05, 6.316265e-05, 2.075344e-05, 0, 3.0129e-06, 2.324237e-05, 
    0.000113777, 0.0001698785, 0.00015665, 0.0001296179, 0.0009469871, 
    0.008330919, 0.5165862, 4.992137, 43.18823, 71.81859, 35.90929, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2.503395, 25.03395, 88.04689, 354.7559, 
    6004.943, 16409.19, 15509.86, 12546.42, 3742.923, 42.25773, 5.264567, 
    2.8305, 5.326696, 15.32724, 30.92193, 43.84749, 47.91269, 49.12563, 
    35.10263, 15.20442, 3.036953, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0.5427925, 5.427925, 366.3095, 1484.653, 2826.97, 3294.921, 
    3195.865, 2993.446, 2979.8,
  3055.147, 5109.396, 9307.208, 9146.649, 8966.816, 7453.676, 5253.157, 
    3567.171, 3072.659, 3428.544, 3602.701, 3417.587, 2882.715, 2420.951, 
    2273.853, 4343.434, 8572.577, 8345.433, 7586.683, 4262.282, 1355.831, 
    1133.536, 1189.682, 1726.767, 2300.862, 2381.619, 2416.113, 1453.18, 
    981.9581, 2164.802, 3463.696, 3352.932, 2993.123, 2519.884, 2195.393, 
    2303.091, 2806.405, 3640.717, 6162.927, 14929.24, 19148.79, 17773.22, 
    13375.82, 8162.993, 4407.082, 3639.264, 3293.916, 2860.534, 2352.018, 
    866.4679, 112.2928, 15.44104, 1.985828, 0.2083054, 0.01647816, 
    0.06649213, 0.09096705, 0.08039964, 0.04783211, 0.01217435, 0, 
    9.725224e-05, 0.0001945045, 9.725224e-05, 0, 0, 0, 0, 0, 0, 0, 
    2.531394e-05, 0.0001242813, 0.0003054829, 0.0003735587, 0.000263094, 
    0.0001526293, 0.005872489, 0.01159235, 0.009555552, 0.004078126, 
    0.00086129, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12.18207, 
    121.8207, 423.091, 1672.676, 10029.7, 15455.87, 13523.64, 7733.477, 
    1986.201, 32.31912, 4.189516, 0, 4.52128, 16.53511, 23.59781, 25.82513, 
    11.03286, 0.3144428, 0.03189252, 0.0002134402, 2.134403e-05, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.5116178, 5.116178, 162.6619, 
    896.613, 2372.922, 3530.032, 3646.353, 3634.577, 3245.531,
  3283.337, 3711.515, 4985.197, 6066.814, 6730.332, 6386.199, 5192.914, 
    3474.561, 2073.384, 1786.675, 1732.579, 1822.753, 2192.615, 3483.156, 
    5232.862, 7474.515, 8234.807, 7443.808, 5084.817, 2775.839, 2010.847, 
    6725.622, 11440.4, 10595.31, 8399.666, 7929.787, 7210.076, 4025.312, 
    1664.235, 1918.582, 2501.081, 3030.025, 4700.295, 12097.47, 22202.49, 
    28724.76, 30690.98, 22944.04, 19152.98, 24170.64, 29188.29, 23834.74, 
    10366.88, 6823.814, 5148.751, 3112.499, 2408.294, 2377.76, 2347.226, 
    1098.206, 25.29284, 13.28064, 8.536497, 1.760471, 0.04350151, 0.06927542, 
    0.09504934, 0.09526344, 0.090998, 0.02888825, 0, 1.458957e-05, 
    2.917915e-05, 1.458957e-05, 0, 0, 0, 0, 0, 0, 0, 0.0001814395, 
    0.000567019, 0.00059721, 0.0006058394, 0.0002144353, 2.289713e-05, 
    0.0008809784, 0.00173906, 0.001139889, 0.0001851772, 1.851773e-05, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01770066, 0.1770066, 49.13077, 
    487.5906, 2109.168, 5459.638, 12064.87, 14535.17, 11621, 4074.156, 
    850.9163, 66.31211, 14.0235, 9.63337, 18.59739, 28.65586, 31.15281, 
    32.28168, 10.67208, 0.03574489, 0.003598918, 1.163174e-05, 1.163174e-06, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.929339, 42.27567, 
    87.36065, 228.9771, 1444.881, 3686.241, 4424.486, 4561.776, 3703.396,
  4027.708, 3754.506, 3736.299, 4034.036, 4331.772, 4370.158, 4339.537, 
    2940.553, 1138.878, 922.5051, 913.3685, 943.7209, 1236.99, 3259.064, 
    5941.942, 7914.887, 8546.191, 6036.925, 2838.467, 2495.55, 2227.867, 
    9618.218, 13234.77, 11893.77, 10552.76, 11126.71, 11700.67, 9735.828, 
    4702.807, 2622.526, 1707.126, 5367.197, 13806.21, 29327.23, 42061.27, 
    45116.36, 45681.5, 37187.01, 33030.13, 35003.83, 36977.52, 27543.87, 
    9923.114, 7216.137, 6032.086, 2738.232, 1618.976, 1965.846, 2312.716, 
    1161.733, 10.7493, 20.46134, 30.17338, 15.17977, 0.1235669, 0.09482128, 
    0.09079064, 0.0906195, 0.09044836, 0.04463742, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0.0002050641, 0.0006241083, 0.0006241083, 0.0006241083, 
    0.0002050641, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0.08813155, 0.8813156, 106.8329, 1049.821, 4552.43, 9436.12, 13119.54, 
    14299.83, 10277.9, 3816.146, 1050.287, 228.8568, 69.41581, 53.20367, 
    63.91631, 74.62895, 69.70553, 51.20368, 14.19486, 0.01968144, 
    0.001968145, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16.16133, 56.56831, 61.52875, 68.03884, 990.4819, 3551.222, 5677.322, 
    6344.292, 5640.685,
  8334.229, 5538.318, 3378.479, 3013.114, 2811.058, 2200.346, 1573.707, 
    840.6031, 602.707, 657.8317, 712.9565, 455.4032, 197.8499, 1119.172, 
    3753.432, 5924.458, 6604.897, 4495.365, 2385.832, 6299.659, 13451.68, 
    13569.7, 13394.99, 11739.78, 10929.78, 13578.75, 16227.72, 14526.04, 
    10066.23, 7633.602, 6853.006, 22741.5, 44394.36, 47827.09, 48635.24, 
    48624.09, 48564.85, 47122.41, 44816.61, 43959.7, 42052.57, 30271.87, 
    13623.43, 9290.118, 7304.171, 3289.382, 1098.996, 756.032, 604.5485, 
    164.6514, 13.48431, 282.5078, 551.5313, 494.4341, 313.3124, 107.9023, 
    13.98646, 1.424052, 0.0120978, 0.00120978, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3.519355e-05, 0.0001071108, 0.0001071108, 0.0001071108, 3.519355e-05, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001968509, 
    0.01968509, 13.56637, 135.2504, 444.3691, 1603.711, 6276.943, 11771.95, 
    13725.86, 14202.6, 10259.48, 4705.362, 1885.401, 547.4364, 354.0567, 
    362.5631, 626.8765, 756.2214, 505.8356, 87.72078, 9.406565, 0.3009069, 
    0.0298042, 0, 0.00127336, 0.002546721, 0.00127336, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 12.81702, 25.63404, 24.74879, 22.93978, 318.791, 
    2217.82, 6941.589, 10430.18, 9912.614,
  9002.199, 6114.318, 3275.98, 2597.876, 2256.489, 1299.472, 576.6361, 
    386.071, 360.7826, 547.1066, 638.2865, 357.1578, 76.02911, 911.7817, 
    3309.571, 5316.399, 5948.852, 4131.548, 2314.243, 8350.698, 14459.67, 
    14127.1, 13026.46, 11502.5, 10954.16, 13796.59, 16639.01, 16472.96, 
    16133.64, 16289.65, 18040.31, 33199.76, 47644.46, 48929.42, 49188.43, 
    49063.76, 48692.7, 47697.13, 46044.05, 45014.1, 42529.75, 31021.44, 
    17027.11, 11808.49, 8588.955, 3826.261, 1005.783, 392.3622, 199.0922, 
    52.86374, 24.67838, 291.9814, 847.4424, 860.9953, 861.1076, 412.4296, 
    70.92799, 7.092802, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01002538, 0.1002538, 
    152.9566, 853.0485, 1587.328, 3499.364, 9809.842, 14504.59, 14363.61, 
    14092.87, 10626.83, 5743.709, 2864.277, 1235.472, 847.0808, 796.5154, 
    1502.504, 1847.987, 1322.484, 274.0869, 30.46671, 1.454713, 0.1451254, 0, 
    0.001537174, 0.003074347, 0.001537174, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2.806806, 5.738173, 5.756338, 5.774503, 118.3983, 1131.214, 
    5668.826, 10987.68, 10465.35,
  4453.382, 4444.296, 4312.858, 3320.154, 1980.198, 959.9561, 354.4422, 
    305.9574, 312.3501, 344.0156, 520.9127, 1420.691, 2639.379, 3387.924, 
    4107.581, 4888.621, 5812.975, 6799.593, 8218.118, 12174.11, 13697.18, 
    12913.94, 10990.04, 10418.88, 10224.3, 11353.37, 14068.08, 17728.52, 
    22680.87, 30614.99, 37902.17, 40172.58, 41395.4, 44523.77, 46910.95, 
    47699.56, 47935.88, 45343.47, 41748.73, 41151.15, 40239.11, 31532.68, 
    17890.93, 13176, 10023.83, 5019.011, 1446.483, 501.8279, 241.7507, 
    122.0243, 90.19643, 392.7239, 851.4245, 1118.041, 1366.701, 1783.907, 
    1928.138, 966.1382, 1.417285, 0.1417285, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.185668, 11.85668, 913.7239, 3845.933, 6575.704, 9720.66, 14176.46, 
    17450.35, 18440.54, 18841.76, 13334.33, 5881.481, 3427.567, 2402.509, 
    1504.389, 1251.98, 2317.755, 3383.53, 3129.682, 2288.295, 652.0761, 
    9.263658, 0.9262993, 0, 0.0002970998, 0.0005941995, 0.0002970998, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0.003956311, 0.03956312, 0.1558609, 0.7277833, 
    6.483573, 10.93317, 5.657239, 0.3813055, 0.3819115, 0.3859804, 17.15372, 
    168.0198, 2010.386, 4265.673, 4436.107,
  3338.927, 4065.967, 4337.894, 3589.309, 1625.064, 774.8335, 365.0817, 
    312.0392, 308.3446, 341.803, 521.8065, 2324.917, 5318.378, 6000.825, 
    6058.72, 5900.687, 5823.352, 9753.115, 13682.88, 12898.29, 10556.73, 
    8544.827, 7306.176, 7508.342, 8080.355, 8500.815, 9645.401, 14891.37, 
    23522.68, 35214.81, 39284.42, 35341.99, 31399.57, 32669.14, 36684.66, 
    41438.75, 43092.38, 40019.15, 34456.83, 34093.84, 33730.84, 27951.29, 
    18385.01, 14423.69, 11301.04, 7135.598, 3561.15, 1198.047, 441.0194, 
    488.6789, 574.2508, 712.0646, 919.9036, 1124.669, 1400.144, 2088.462, 
    2349.582, 1185.576, 7.386838, 0.7386842, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    6.126528, 61.26528, 2355.501, 8478.848, 11922.99, 14908.32, 17940.61, 
    19592.3, 19944.99, 20277.66, 14318.23, 6312.471, 3950.649, 3002.436, 
    1906.601, 1601.675, 2545.651, 3512.603, 3632.229, 3723.136, 1297.421, 
    40.58969, 4.058971, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01986783, 
    0.1986783, 1.178653, 4.184587, 10.95764, 13.55257, 6.776284, 0, 0, 0, 
    6.393955, 63.93956, 963.6639, 2851.163, 3175.456,
  4298.801, 2062.664, 920.8984, 814.0658, 798.3642, 791.5525, 835.8483, 
    1697.305, 2200.395, 1885.829, 1571.264, 2724.866, 5928.787, 7762.52, 
    9294.182, 9928.06, 10653.31, 13826.34, 15081.88, 10845.39, 2968.827, 
    1887.699, 1709.203, 1945.471, 2596.045, 3289.134, 5196.128, 11867.77, 
    20460.19, 30819.93, 34268.41, 28468.49, 15595.5, 14117.83, 14126.4, 
    17336.92, 22023.92, 25215.6, 26930.8, 25158.81, 21828.64, 16970.44, 
    13614.15, 13322.57, 13030.99, 10576.58, 7267.65, 2592.705, 966.6252, 
    1787.57, 2608.515, 2359.741, 1573.012, 641.9683, 318.1509, 785.4734, 
    1252.796, 667.6419, 28.24926, 2.824939, 5.526755e-06, 5.526757e-07, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 82.4919, 824.919, 5691.188, 14309.38, 16218.79, 17086.06, 
    19203.04, 20466.59, 20625.42, 20294.11, 14389.55, 6834.271, 4287.786, 
    3126.744, 2077.73, 1786.833, 2076.519, 2602.326, 3435.04, 3735.823, 
    2664.732, 549.7286, 65.51551, 5.020367, 0.5022584, 0.0001054785, 
    1.054786e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0551688, 0.551688, 5.58856, 
    13.9432, 13.95912, 13.88786, 4.543471, 0, 0, 0, 52.46457, 524.6458, 
    3636.868, 6349.467, 5861.98,
  4563.516, 1282.257, 72.51356, 203.6391, 646.0788, 957.9147, 1513.36, 
    3432.68, 4188.054, 3502.384, 2816.715, 3565.953, 5868.405, 7766.964, 
    9637.441, 11001.71, 12253.35, 14429.06, 15191.19, 8292.891, 1169.994, 
    1073.615, 1049.234, 1026.934, 1007.501, 1243.103, 2410.172, 7158.683, 
    14703.08, 22615.79, 25188.93, 22190.98, 14587.26, 12120.73, 11361.32, 
    11543.08, 12392.79, 17174.17, 19288.12, 18645.18, 16512.02, 13597.04, 
    12551.62, 12679.66, 12941.31, 12540.38, 10360.28, 4587.138, 2325.849, 
    2577.455, 3091.607, 3061.542, 2723.284, 830.9799, 8.564355, 395.6646, 
    782.7648, 550.3969, 108.9141, 10.89147, 2.949471e-05, 2.949472e-06, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 136.5073, 1365.073, 6943.611, 14940.53, 16572.86, 
    17305.41, 19310.99, 20534.92, 20680.79, 20296.63, 14385.51, 6875.251, 
    4394.726, 3298.972, 2331.375, 2002.168, 2050.769, 2250.732, 3307.589, 
    3761.17, 3200.79, 1622.428, 431.8878, 26.79226, 2.68041, 0.0005629089, 
    5.629091e-05, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.06003961, 0.6003962, 6.67866, 
    14.77644, 13.5287, 9.61285, 2.644635, 0, 0, 0, 65.0817, 650.817, 
    4248.739, 7354.995, 6696.75,
  4224.925, 3981.772, 3662.095, 2701.654, 2010.964, 1971.03, 2006.109, 
    3764.353, 4860.783, 4561.546, 3590.205, 2308.265, 1428.551, 1593.735, 
    2403.438, 4458.882, 6966.755, 9530.998, 10337.77, 5510.771, 683.7723, 
    865.2954, 1046.819, 938.2795, 716.4822, 787.249, 1457.103, 3855.34, 
    7372.632, 11296.75, 14742.92, 16392.32, 16921.34, 16120.37, 14620, 
    12069.85, 11135.44, 12469.96, 15220.94, 15163.83, 15071.9, 14149.7, 
    12759.06, 11550.1, 11183.77, 11287.68, 11391.6, 9434.746, 4498.341, 
    2848.219, 2576.234, 3359.484, 3742.776, 2714.771, 1042.511, 806.3749, 
    708.9637, 648.4571, 577.3096, 199.7574, 18.07093, 1.826424, 0.009204946, 
    0.000920495, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 150.0266, 1500.266, 6759.081, 13835.93, 
    15990.43, 17120.59, 19257.11, 20500.07, 19714.97, 16622.06, 11626.33, 
    6698.062, 4641.275, 3614.984, 2848.094, 2527.021, 2337.137, 2282.994, 
    2543.493, 2803.991, 2787.38, 2613.573, 1732.07, 677.5757, 271.1879, 
    107.6971, 31.05568, 7.525509, 1.043384, 0.3579758, 0.6649, 0.815097, 
    0.4075485, 0, 0, 0, 0.01421513, 0.1421513, 1.86291, 3.310738, 2.727193, 
    1.159313, 0.2441388, 0, 0, 0, 57.29291, 572.9291, 3393.192, 5113.431, 
    4875.333,
  3621.763, 4286.131, 4701.332, 4824.497, 4888.39, 3778.195, 3234.908, 
    3809.512, 4983.703, 4930.535, 4446.953, 1523.233, 237.1691, 222.8629, 
    329.214, 1138.249, 2307.146, 3640.61, 4081.329, 2198.348, 315.3671, 
    674.3353, 1033.303, 920.4101, 689.7151, 804.3731, 1476.213, 3140.122, 
    5241.853, 6358.244, 8103.128, 13756.99, 17795.9, 17268.36, 15686.33, 
    12309.32, 10988.81, 12145.79, 14683.5, 14896.49, 14907.46, 14333.81, 
    13240.59, 11344.13, 10648.92, 11095.93, 11542.93, 10327.66, 6782.411, 
    3596.262, 2567.729, 3238.345, 3908.961, 3440.149, 2110.567, 1105.044, 
    686.5446, 667.6371, 648.7297, 294.0605, 23.68432, 2.474126, 0.05032977, 
    0.00503298, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 151.1708, 1511.708, 6088.523, 11675.88, 
    14297.45, 16229.14, 19176.23, 20141.12, 17795.51, 11478.22, 8462.438, 
    6159.946, 4549.039, 3620.055, 3255.154, 3057.844, 2582.311, 2278.062, 
    2296.152, 2396.492, 2947.436, 3189.396, 2851.344, 1831.126, 971.5247, 
    304.7525, 109.1979, 47.67542, 8.969041, 1.9573, 3.635466, 4.456697, 
    2.228348, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 54.0519, 410.9632, 
    1293.429, 2327.227, 3023.014,
  1869.843, 2958.134, 4284.671, 6896.323, 7852.362, 7112.238, 5116.064, 
    3873.414, 3502.477, 4241.618, 4603.325, 3378.394, 803.2982, 511.2549, 
    524.5376, 850.378, 1176.218, 1140.456, 959.2375, 243.7763, -57.44519, 
    316.6017, 933.3474, 982.4276, 1031.508, 1205.234, 1669.086, 3043.192, 
    4705.797, 5711.383, 6895.949, 9335.889, 11570.17, 11981.15, 12350.31, 
    14420.31, 16258.99, 16510.73, 16688.62, 18036.86, 18572.96, 16699.52, 
    13078.75, 12726.38, 12419.12, 10700.18, 8925.619, 8504.798, 7872.035, 
    4131.751, 2620.707, 2823.513, 3026.32, 2841.689, 2359.529, 2268.011, 
    2100.098, 1032.432, 217.4225, 67.00245, 24.44584, 7.538375, 2.47066, 
    0.3227327, 0.01607235, 0.001607236, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6.84289e-08, 6.84289e-07, 0.2015235, 
    2.015221, 229.5406, 1643.73, 4932.104, 8718.222, 11475.9, 13626.65, 
    15240.85, 15755.6, 12844.1, 8713.724, 6861.263, 5555.59, 4291.986, 
    3607.958, 3534.449, 3472.963, 3008.378, 2664.546, 2697.526, 2831.432, 
    3241.15, 3570.126, 3354.302, 2580.564, 1462.56, 496.4689, 181.1405, 
    133.503, 365.1931, 478.5734, 256.5378, 11.81578, 1.181578, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 10.69416, 62.82728, 131.7627, 322.6013, 920.351,
  829.1974, 1772.112, 3279.751, 6890.893, 8296.772, 7620.572, 5536.924, 
    3302.836, 2540.577, 3585.618, 4623.03, 3366.501, 1338.294, 986.3846, 
    951.4275, 994.7183, 1014.666, 880.2568, 478.7102, 52.18144, -92.38046, 
    153.6995, 858.4072, 1386.925, 1812.816, 1891.273, 1976.18, 2835.739, 
    4252.836, 5389.513, 5743.698, 5304.422, 4741.751, 5874.729, 9726.579, 
    15580.22, 17780.96, 17744.36, 17691.8, 18780.72, 19828.5, 17039.68, 
    13307.66, 13112.02, 12936.96, 10550.52, 8089.253, 7901.796, 7710.904, 
    5027.749, 2770.005, 2667.455, 2689.251, 2888.474, 3086.545, 3027.797, 
    2573.429, 968.451, 133.0974, 44.82969, 24.49408, 20.10136, 17.58864, 
    5.212841, 0.1634679, 0.01008262, 0.0001341424, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.711185e-09, 4.292731e-07, 
    0.0168232, 1.264211, 14.84419, 276.9024, 1685.249, 4707.084, 8175.964, 
    11739.61, 12877.72, 12025.44, 9634.461, 8159.865, 6838.042, 5708.325, 
    4788.454, 4012.284, 3592.159, 3551.116, 3510.662, 3135.581, 2810.054, 
    2845.599, 2993.814, 3332.858, 3588.184, 3629.63, 3591.608, 2504.164, 
    1131.467, 635.0035, 567.1837, 617.8143, 639.1492, 341.4353, 18.27176, 
    1.518201, 0.02019863, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.0001242849, 
    0.009341695, 0.286461, 14.81096, 97.65171, 297.8567,
  616.1959, 933.5225, 1612.562, 3701.627, 4691.45, 4479.272, 3716.574, 
    2673.199, 2289.833, 2574.776, 2852.045, 2169.438, 1480.709, 1506.274, 
    1548.078, 1525.576, 1447.768, 1388.266, 1254.434, 703.4572, 376.046, 
    760.6616, 1804.532, 2548.383, 2768.372, 2477.158, 2199.089, 2948.907, 
    3784.274, 3851.289, 3849.51, 3444.168, 3073.368, 4567.198, 9201.229, 
    14842.15, 16892.97, 16603.57, 16301.97, 17762.5, 19139.77, 15407.61, 
    11315.25, 11033.39, 10823.42, 9671.521, 8253.874, 7887.806, 7514.805, 
    5882.668, 3732.122, 3016.707, 2926.87, 3953.965, 4966.728, 4270.909, 
    2310.015, 821.9142, 168.2393, 28.83576, 9.929073, 115.7448, 221.3261, 
    194.0541, 109.2159, 28.67975, 1.273596, 3.872284, 7.742311, 8.192957, 
    8.59605, 10.60003, 15.65613, 24.33968, 27.6294, 24.66513, 16.89874, 
    13.72892, 10.6173, 3.270801, 0.2223162, 0.02286031, 0.000575284, 
    1.488414e-05, 3.112247e-07, 0, 0, 0, 0.01117321, 0.5343521, 4.23234, 
    35.38763, 242.9999, 2402.458, 7454.373, 10502.33, 12218.21, 12841.35, 
    12902.82, 11240.89, 7870.032, 6824.058, 6162.082, 4974.22, 3971.849, 
    3511.869, 3422.505, 3417.08, 3405.382, 3054.527, 2208.838, 1866.73, 
    1810.518, 2266.319, 3533.789, 4627.536, 4980.069, 4604.185, 3520.005, 
    2732.957, 1962.776, 1201.872, 564.5768, 123.6271, 7.088471, 0.6687093, 
    0.0139826, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001609631, 0.07697967, 1.933839, 
    61.87172, 180.5434, 221.9014, 281.0804, 391.5906,
  472.0515, 467.3549, 477.9736, 804.7759, 1189.496, 1235.597, 1280.076, 
    1617.02, 1891.82, 1773.485, 1562.63, 1505.62, 1502.26, 1671.582, 
    1838.288, 1757.387, 1614.956, 1578.042, 1532.734, 1239.469, 1018.51, 
    1320.033, 2151.69, 2827.719, 3034.942, 2624.362, 2222.343, 2666.052, 
    3117.578, 2934.854, 2428.748, 2111.943, 2069.679, 3608.799, 7922.406, 
    12014.07, 13419.85, 13145.33, 12883.41, 14567.59, 16129.91, 12280.71, 
    8403.296, 9135.247, 9986.253, 9590.307, 8510.227, 8033.65, 7488.721, 
    6453.073, 5344.52, 4168.401, 3807.68, 4856.424, 5878.856, 4709.488, 
    1788.641, 608.9147, 175.2914, 25.8842, 10.06629, 276.5886, 587.8848, 
    624.8894, 619.4321, 316.5376, 13.61602, 6.608661, 10.75594, 11.38797, 
    11.96856, 14.77256, 21.81055, 33.76052, 38.35157, 35.27939, 32.25827, 
    38.0966, 43.35369, 23.17871, 1.594479, 0.1374372, 0.004354308, 
    8.952449e-05, 2.476268e-06, 0, 0, 0, 0.08889983, 3.213995, 25.31153, 
    197.6442, 1141.162, 4942.73, 10924.12, 13258.81, 13646.64, 13569.15, 
    12983.57, 9960.736, 6689.727, 5992.488, 5552.191, 4353.973, 3334.934, 
    3003.588, 2952.277, 3043.062, 3117.576, 2568.256, 1233.847, 677.5527, 
    589.5603, 1368.039, 3401.079, 4811.557, 5235.04, 5030.375, 4277.692, 
    3355.465, 2322.218, 1206.165, 381.2845, 56.45422, 1.753268, 0.03105236, 
    0.0008589154, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.003095225, 0.1119016, 
    2.381527, 55.92402, 233.828, 505.4794, 608.7241, 543.9604,
  357.0723, 120.6344, 61.34686, 127.3295, 304.7637, 404.9247, 522.8275, 
    714.3574, 930.5607, 1154.545, 1355.962, 1465.894, 1571.001, 1824.141, 
    1919.62, 1744.43, 1541.015, 1518.148, 1498.132, 1359.432, 1253.746, 
    1472.598, 2118.694, 2828.851, 3062.692, 2458.146, 1844.728, 1856.824, 
    1885.363, 1645.192, 1403.982, 1412.868, 1540.604, 2192.418, 3689.093, 
    5204.815, 6629.535, 7526.166, 8153.677, 8718.201, 8851.104, 8067.386, 
    7326.736, 8442.178, 10079.19, 10445.24, 10483.33, 10022.76, 8743.932, 
    7514.336, 7082.815, 7123.196, 7176.43, 7045.583, 6237.688, 3507.743, 
    923.0684, 226.389, 57.39295, 8.805112, 6.43089, 160.5515, 864.0469, 
    2444.178, 3042.025, 1613.436, 108.5752, 13.27877, 5.70259, 3.93312, 
    3.678826, 4.492989, 6.837564, 8.418112, 11.41802, 17.33771, 33.5055, 
    84.14813, 110.6598, 111.8053, 110.6831, 83.66249, 26.28082, 5.750628, 
    1.168366, 0.1664781, 0.009735069, 0.1198616, 1.366676, 19.59615, 
    151.2029, 1186.36, 4216.755, 8677.356, 11106.95, 11663.29, 11735.98, 
    11346.47, 9927.729, 7835.325, 5876.235, 5093.749, 4595.718, 3669.694, 
    2838.558, 2455.381, 2259.654, 2160.89, 2034.575, 1475.063, 633.4224, 
    321.5034, 297.8602, 1021.911, 2939.894, 4493.593, 5004.958, 4923.212, 
    4378.431, 3204.702, 1866.629, 715.5723, 168.1547, 24.35201, 0.8593246, 
    0.005372726, 0.0001826637, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002774625, 
    0.08161065, 1.49309, 29.88909, 196.2509, 703.3244, 964.2495, 796.1766,
  273.2705, 57.31008, 17.7017, 62.98434, 202.5874, 373.402, 435.0912, 
    366.1121, 306.4013, 552.2848, 1147.91, 1410.428, 1601.105, 1848.283, 
    1924.147, 1707.644, 1487.134, 1480.446, 1484.783, 1466.22, 1454.2, 
    1596.254, 2070.598, 2797.305, 3047.542, 2263.777, 1223.598, 1019.724, 
    989.7657, 991.3171, 1008.952, 1087.53, 1258.366, 1388.835, 1650.392, 
    2226.841, 3011.76, 4293.548, 4800.803, 4753.561, 4691.482, 4928.021, 
    6031.606, 8184, 10197.88, 11045.54, 11173.12, 10688.11, 9322.009, 
    7914.998, 7421.032, 7792.68, 8176.059, 7883.747, 6350.688, 2948.468, 
    736.2673, 114.9843, 8.000487, 1.014349, 11.24428, 245.3345, 1194.359, 
    3099.693, 3809.844, 2149.437, 253.1445, 31.55309, 4.15533, 0.5229882, 
    0.02118232, 5.223471e-05, 0.000136455, 0.003363488, 0.4076503, 8.618091, 
    35.89153, 61.49408, 120.3076, 304.2905, 401.0199, 337.516, 165.6502, 
    50.43607, 7.928592, 1.026524, 0.0705343, 0.739081, 7.870408, 94.50394, 
    636.2975, 3385.333, 8408.953, 10646.47, 11082.26, 10419.13, 8527.109, 
    6694.352, 5710.436, 5467.085, 5284.465, 4832.367, 4225.356, 3521.723, 
    2800.085, 2164.332, 1595.66, 1110.113, 709.1466, 364.0709, 198.316, 
    150.5752, 174.3104, 812.5056, 2418.88, 3461.276, 4057.604, 4276.913, 
    4262.92, 3231.851, 1041.487, 226.2125, 43.3772, 6.219241, 0.2633108, 
    0.00268155, 0.0001071255, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.001188917, 
    0.02976082, 0.9837314, 20.49695, 143.4929, 664.9965, 1019.288, 805.9467,
  199.5036, 559.7615, 1368.661, 1686.199, 1725.674, 1408.613, 651.2661, 
    228.2821, 122.2374, 274.7659, 603.1923, 729.853, 892.7899, 1373.532, 
    1624.816, 1555.445, 1470.548, 1469.892, 1490.243, 1524.607, 1611.448, 
    1799.698, 2044.824, 2385.378, 2471.687, 1745.904, 858.0121, 705.1477, 
    691.1343, 789.5295, 904.7668, 921.863, 936.338, 1023.349, 1266.476, 
    1543.889, 2019.145, 3183.455, 3695.904, 3648.986, 3582.719, 3789.23, 
    4540.41, 5584.257, 6835.241, 8551.154, 9194.319, 8810.062, 7824.618, 
    7378.58, 7084.922, 6918.388, 6674.649, 6111.888, 5274.389, 4067.579, 
    2751.276, 1275.281, 736.7509, 729.4831, 842.5641, 1063.176, 1403.018, 
    2015.808, 2215.978, 1384.851, 384.0168, 228.6789, 172.1617, 73.2657, 
    17.71258, 2.803346, 0.3051336, 0.192905, 0.4367617, 4.404183, 19.24811, 
    38.69632, 94.66923, 358.7358, 862.2708, 1243.353, 1339.862, 929.4676, 
    489.4691, 446.7501, 471.6281, 957.3195, 2310.904, 3366.78, 4988.295, 
    8958.783, 10710.58, 10812.86, 10721.12, 9351.945, 6366.034, 5168.224, 
    4503.483, 3963.251, 3825.768, 3975.202, 4118.369, 3874.093, 3051.106, 
    1987.783, 960.6908, 335.4461, 97.62226, 32.30099, 21.61102, 31.4383, 
    139.6652, 1058.974, 1894.134, 1857.467, 1793.484, 2206.535, 2573.738, 
    1775.337, 459.4362, 72.59965, 7.781445, 7.765491, 29.4802, 143.0737, 
    226.9517, 133.2316, 18.75097, 2.075993, 0.09453375, 0, 0, 0, 0, 0, 
    0.0001945202, 0.004271728, 0.2617964, 5.255436, 53.29734, 435.3299, 
    760.0071, 479.5158,
  98.68642, 603.4781, 1980.055, 3357.826, 3829.68, 3201.024, 1595.411, 
    470.4556, 121.6332, 260.681, 474.8007, 523.0399, 570.9604, 800.0818, 
    1199.682, 1380.767, 1448.484, 1470.433, 1491.768, 1546.767, 1642.768, 
    1789.715, 1954.038, 2138.024, 2157.042, 1507.49, 770.5862, 662.5842, 
    657.8714, 747.992, 838.4329, 841.4561, 841.5451, 907.1511, 1138.242, 
    1424.872, 1917.049, 3067.011, 3570.299, 3527.668, 3468.949, 3718.174, 
    4090.479, 4190.989, 4324.411, 5123.824, 5779.889, 5491.065, 5176.29, 
    5485.419, 5776.465, 5227.023, 4653.114, 4634.53, 4821.782, 5789.817, 
    6474.552, 5195.113, 3567.834, 3267.032, 3055.764, 2424.587, 1817.742, 
    1629.752, 1491.239, 1094.804, 872.0292, 926.1841, 969.0388, 604.6012, 
    123.55, 17.69025, 1.969334, 1.15446, 1.384266, 3.339799, 11.25138, 
    27.03794, 83.48055, 387.8696, 1177.545, 2351.454, 2815.144, 2541.7, 
    2238.275, 2273.491, 2629.855, 4037.555, 6481.199, 7840.586, 9106.954, 
    11263.74, 12124.95, 11744.09, 10014.66, 6867.471, 4585.398, 3828.121, 
    3610.006, 3534.759, 3538.54, 3770.008, 3992.125, 3840.986, 3170.267, 
    2008.129, 847.829, 187.8159, 16.59301, 1.321063, 0.8789353, 13.75641, 
    126.1771, 850.4488, 1473.657, 1397.517, 1282.843, 1398.084, 1478.856, 
    904.0096, 170.8742, 22.3856, 2.611001, 24.86806, 180.9864, 879.3412, 
    1366.793, 807.7869, 120.6417, 13.13582, 0.6670913, 0, 0, 0, 0, 0, 0, 0, 
    0.1022, 2.012439, 23.78635, 197.8849, 347.1036, 211.8065,
  46.07317, 460.2399, 1764.575, 3674.762, 4476.393, 4409.362, 3686.29, 
    1583.041, 346.7863, 364.2673, 636.6653, 772.4763, 865.0372, 935.4399, 
    1000.869, 1087.15, 1185.448, 1295.854, 1411.62, 1529.62, 1637.146, 
    1701.615, 1796.47, 2048.812, 2125.245, 1461.631, 774.5488, 705.654, 
    707.4476, 749.3987, 800.3044, 810.3776, 819.8871, 879.0637, 1096.375, 
    1489.464, 2097.43, 3186.153, 3665.126, 3705.81, 3721.98, 3863.985, 
    3997.289, 3966.496, 3834.5, 3690.227, 3455.574, 2935.934, 2704.578, 
    2725.281, 2926.85, 3422.395, 4057.387, 4451.314, 5294.912, 8289.92, 
    10311.86, 10317.95, 9558.956, 8045.896, 6392.046, 5210.026, 4420.378, 
    4095.688, 3819.334, 3034.82, 2579.514, 2687.193, 2785.549, 2182.657, 
    824.7855, 203.0802, 60.96211, 49.62323, 49.2061, 50.90456, 59.30486, 
    79.65081, 153.286, 498.878, 1300.311, 2200.948, 3279.279, 4599.774, 
    5920.161, 6971.718, 7917.793, 8961.377, 9636.501, 9866.497, 10160.95, 
    11498.19, 12491.41, 11700.48, 8980.263, 5157.008, 3272.001, 2935.585, 
    2917.721, 3230.637, 3603.329, 3672.176, 3667.097, 3472.032, 2809.673, 
    1834.003, 872.0687, 280.2261, 80.48344, 39.80149, 34.162, 45.94137, 
    131.2656, 553.2593, 1174.478, 1403.821, 1445.537, 1439.234, 1345.224, 
    697.6266, 105.3467, 51.32418, 108.9836, 951.3167, 4054.419, 9714.545, 
    11758.11, 6768.73, 989.0098, 103.1369, 9.409161, 0.7968252, 0.2380682, 
    2.891445, 52.67084, 486.5985, 898.1776, 870.2485, 635.548, 215.6295, 
    33.11486, 44.89764, 68.59998, 43.4179,
  16.62835, 217.5286, 1193.975, 3441.465, 4521.975, 4548.044, 4098.187, 
    2398.798, 1136.582, 1022.143, 1080.246, 1287.132, 1415.474, 1228.779, 
    988.8677, 939.8303, 936.3417, 973.6841, 1123.628, 1418.596, 1552.076, 
    1548.906, 1563.51, 1851.755, 2073.905, 1442.779, 782.816, 723.2269, 
    730.5637, 724.4543, 718.6313, 732.7651, 784.8634, 859.6174, 1054.082, 
    1620.962, 2555.095, 3584.615, 4161.685, 4327.568, 4345.479, 4224.834, 
    4003.324, 3912.083, 3784.002, 3448.906, 2964.08, 2413.278, 2194.168, 
    2186.653, 2279.853, 2841.909, 3996.177, 4627.846, 5832.009, 9195.511, 
    11130.83, 11247.5, 10865.84, 9434.872, 7138.947, 6077.322, 5535.896, 
    5270.646, 5073.761, 4654.472, 4275.379, 4120.647, 3919.965, 3285.203, 
    2178.84, 905.1539, 358.598, 290.6724, 268.0109, 206.6077, 171.3408, 
    195.655, 339.9518, 746.574, 1505.753, 2466.854, 3671.717, 5196.743, 
    6768.64, 8151.192, 9275.109, 10043.58, 10265.68, 10248.2, 10328.9, 
    11453.73, 12449.07, 11020.29, 7285.467, 4241.289, 3009.939, 2805.905, 
    2822.355, 3229.45, 3626.365, 3522.884, 3100.042, 2606.253, 2051.809, 
    1460.398, 939.5403, 625.395, 426.3898, 279.4995, 205.0284, 177.8034, 
    185.0101, 339.7383, 820.8521, 1526.845, 1827.368, 1773.961, 1388.065, 
    504.9514, 82.67303, 69.74248, 297.1117, 1923.769, 7016.029, 15609.27, 
    18812.02, 12693.02, 3336.474, 549.5848, 56.06853, 5.184972, 1.658843, 
    18.84082, 155.3661, 823.313, 1379.476, 1375.859, 1080.378, 393.0328, 
    46.71139, 8.392272, 5.09085, 3.538113,
  3.189973, 43.26501, 247.5215, 827.3576, 1910.177, 3416.357, 4062.477, 
    3980.53, 3421.723, 2368.784, 1882.761, 1893.715, 1923.486, 1644.721, 
    1156.257, 972.0522, 881.2635, 741.1612, 710.3987, 950.2469, 1188.533, 
    1155.991, 1143.992, 1554.414, 1949.042, 1763.875, 1232.036, 872.9573, 
    628.2666, 504.3598, 475.7788, 480.0254, 510.8569, 596.5566, 881.8436, 
    1737.472, 3244.69, 5041.789, 5778.716, 5689.595, 5230.574, 4654.532, 
    4258.872, 4120.839, 3987.121, 3628.733, 3075.683, 2454.515, 2210.814, 
    2343.929, 3153.906, 5145.851, 6224.607, 6158.832, 6214.339, 8181.402, 
    10151.63, 10138.75, 9008.122, 6661.284, 4824.422, 4138.307, 4011.619, 
    4088.826, 4339.273, 4673.167, 4803.193, 4655.706, 4233.21, 3811.907, 
    3331.023, 2775.828, 2151.803, 1419.217, 770.3688, 393.4391, 298.7045, 
    360.2911, 666.5513, 1310.365, 2209.688, 3230.128, 4336.919, 5515.042, 
    6542.624, 7122.479, 7590.257, 8350.04, 8652.084, 8392.514, 8104.088, 
    8104.814, 8033.252, 6965.617, 4654.517, 3361.601, 2970.992, 2914.944, 
    2932.381, 3128.184, 3292.64, 2993.403, 2258.472, 1747.515, 1410.898, 
    1261.827, 1247.987, 1392.803, 1526.611, 1401.782, 995.9667, 466.6673, 
    240.371, 255.2905, 492.0869, 1373.093, 2287.282, 2549.907, 2466.805, 
    1410.428, 353.0215, 255.4157, 512.5297, 2206.35, 7456.12, 16290.79, 
    20059.1, 17600.54, 11099.42, 6674.449, 3373.823, 1265.786, 534.97, 
    374.3105, 405.1931, 882.3669, 1357.932, 1366.143, 1110.378, 452.7195, 
    56.14806, 3.641754, 0.7297399, 0.3827748,
  0.00019263, 0.002654472, 1.512194, 20.69162, 313.4001, 1973.182, 3766.928, 
    4169.855, 4078.754, 3115.94, 2153.481, 2044.479, 2041.631, 1781.921, 
    1252.329, 994.0853, 786.8528, 440.858, 304.2137, 462.5173, 649.933, 
    683.9755, 742.6394, 1106.454, 1473.159, 1533.787, 1478.919, 1047.49, 
    475.7748, 302.95, 276.814, 291.8497, 350.8531, 453.5312, 753.3114, 
    1688.614, 3420.076, 5493.839, 6361.09, 6156.231, 5439.334, 4805.814, 
    4406.888, 4255.662, 4106.241, 3724.411, 3138.657, 2483.915, 2227.66, 
    2462.542, 3678.045, 6280.396, 7500.283, 6871.093, 6188.502, 6806.564, 
    7457.128, 6829.553, 4911.86, 2692.858, 1568.691, 1323.245, 1321.587, 
    1642.301, 2637.786, 4129.272, 4801.271, 4697.392, 4270.684, 3905.067, 
    3582.229, 3371.015, 2992.121, 2022.301, 916.8237, 425.5467, 328.4216, 
    402.7943, 753.4113, 1478.917, 2451.026, 3523.56, 4492.267, 5137.377, 
    5292.199, 4983.503, 4703.68, 4999.292, 5295.68, 4924.557, 3852.985, 
    2673.365, 2176.463, 2158.16, 2332.393, 2707.115, 2929.605, 2977.771, 
    2976.97, 2895.478, 2583.401, 2024.531, 1427.105, 975.2735, 834.9758, 
    970.2535, 1351.409, 1758.172, 1913.777, 1787.441, 1342.081, 678.2991, 
    370.9211, 340.0984, 433.0469, 1107.382, 2441.325, 3127.526, 3114.02, 
    1822.62, 522.2054, 417.5632, 893.4777, 2861.363, 8151.65, 16908.27, 
    21074.54, 21562.21, 21271.72, 18631.14, 12439.07, 7031.637, 3236.584, 
    1592.772, 1243.611, 1257.498, 1296.75, 1271.76, 1087.526, 507.3484, 
    69.78669, 2.887185, 0.2095176, 0,
  0.216404, 0.0003266071, 0.2196097, 2.740807, 69.55715, 529.4813, 1580.506, 
    2609.531, 2976.833, 2610.672, 1986.323, 1735.874, 1561.534, 1200.464, 
    781.2496, 492.8106, 285.7652, 127.3487, 74.98228, 109.6848, 233.5777, 
    415.7253, 498.0275, 474.8238, 458.4267, 560.6987, 646.0306, 517.4575, 
    311.3895, 236.1087, 225.9978, 255.2029, 340.3347, 449.4733, 719.8087, 
    1494.848, 2892.712, 4571.32, 5293.75, 5072.652, 4428.445, 4031.108, 
    3821.837, 3731.018, 3603.844, 3147.78, 2435.585, 2068.309, 2003.125, 
    2236.228, 3141.135, 4783.87, 5499.745, 4864.38, 3935.071, 3641.809, 
    3394.217, 2611.72, 1483.829, 926.2589, 649.5906, 441.8269, 375.1197, 
    428.7629, 782.3915, 1780.196, 2460.109, 2291.22, 2034.99, 2144.353, 
    2290.885, 2203.998, 1780.178, 1012.875, 413.094, 178.7615, 139.4555, 
    235.8232, 602.0186, 1252.497, 1958.499, 2502.681, 2807.951, 2923.053, 
    3037.968, 3315.118, 3487.8, 3359.797, 2770.459, 1695.784, 946.0918, 
    696.9707, 671.3004, 844.8635, 1306.145, 1860.1, 2190.042, 2290.459, 
    2296.799, 2190.416, 1858.531, 1357.345, 834.9147, 432.463, 351.9552, 
    725.8671, 1116.593, 1180.042, 1189.339, 1264.08, 1327.967, 1273.93, 
    1273.738, 1677.681, 2207.464, 2375.803, 2365.213, 2074.816, 1348.859, 
    546.2054, 209.042, 363.9451, 1338.644, 4164.042, 9535.196, 16507.45, 
    22941.61, 26567.97, 27522.47, 27135.7, 24875.03, 19242.75, 11784.89, 
    6472.699, 3029.191, 1310.271, 724.5215, 552.8309, 431.2688, 187.2048, 
    34.87221, 8.705995, 5.681057, 1.924034,
  0.6389964, 0, 0.02108463, 0.2405119, 2.683905, 21.35813, 123.2247, 
    456.0099, 986.4002, 1372.093, 1460.924, 1169.373, 619.2632, 316.0235, 
    163.4594, 59.44799, 19.75106, 12.55798, 13.57558, 32.64716, 125.4425, 
    329.489, 433.6435, 312.9021, 167.8647, 136.9972, 140.0782, 154.3781, 
    169.6036, 173.713, 180.829, 224.8049, 321.7685, 427.4502, 641.6324, 
    1098.956, 1812.771, 2726.913, 3110.586, 2833.208, 2500.31, 2499.151, 
    2577.237, 2597.494, 2465.471, 1839.474, 1223.298, 1162.64, 1355.259, 
    1610.309, 1802.674, 1883.253, 1812.876, 1398.917, 987.2664, 917.7213, 
    877.5862, 603.9479, 327.1125, 271.9744, 259.2685, 180.161, 95.62258, 
    74.34053, 101.8407, 236.7227, 350.7336, 280.9894, 214.7369, 345.1332, 
    490.3671, 476.0885, 340.6914, 145.5025, 32.50022, 5.00176, 8.300686, 
    67.9511, 289.7647, 677.0028, 859.8763, 764.5149, 641.1469, 671.7164, 
    980.2689, 1726.771, 2182.945, 1773.719, 825.6232, 261.6711, 102.5192, 
    102.6006, 187.3868, 395.0137, 693.1738, 969.6382, 1172.977, 1269.331, 
    1290.79, 1269.335, 1155.505, 853.8105, 453.3684, 223.5125, 221.3925, 
    507.7046, 784.7928, 769.7751, 725.3423, 925.1078, 1348.317, 1662.291, 
    2112.944, 2940.48, 3369.624, 3100.642, 2146.601, 861.3702, 175.1358, 
    37.70462, 73.68847, 554.6742, 2498.554, 6627.016, 12317.3, 18600.09, 
    24173.39, 27644.58, 28756.52, 28783.93, 28052.47, 25072.68, 18973.12, 
    12089.03, 5954.311, 2081.914, 521.4187, 91.26953, 9.264935, 5.871143, 
    10.41281, 10.99227, 8.935199, 4.073005,
  0.4243007, 0, 0.03756952, 0.389131, 2.44396, 12.0915, 40.25931, 93.58552, 
    188.0685, 317.9208, 368.973, 277.4405, 125.5978, 46.17498, 20.08062, 
    7.281125, 2.4337, 1.520232, 3.698236, 25.08646, 153.7794, 455.6624, 
    697.8214, 744.2251, 680.3508, 512.7038, 295.8246, 166.0785, 103.6099, 
    65.65932, 62.02406, 119.7663, 229.8941, 334.1563, 502.8368, 810.3132, 
    1240.672, 1715.066, 1896.44, 1694.344, 1489.131, 1585.405, 1773.205, 
    1843.328, 1743.242, 1294.634, 726.2303, 476.7737, 438.1512, 451.73, 
    461.9936, 421.9794, 326.802, 231.6194, 196.1508, 222.9951, 242.573, 
    190.2422, 114.535, 81.71344, 64.47827, 36.75955, 15.90992, 9.630474, 
    13.08005, 28.4264, 40.76617, 33.7415, 27.23098, 41.44395, 57.8413, 
    56.69011, 40.43542, 18.08325, 4.351353, 0.6529179, 1.787781, 14.35539, 
    59.34385, 132.0752, 163.2566, 128.216, 85.80041, 82.27062, 146.4635, 
    315.1256, 427.5367, 319.9697, 124.2403, 30.48876, 12.20618, 14.01656, 
    43.48259, 163.5527, 413.8749, 710.1328, 927.644, 1022.937, 1037.008, 
    977.9457, 800.5988, 536.2912, 332.2169, 247.5068, 274.9326, 456.1331, 
    668.45, 754.6471, 860.2905, 1243.385, 1820.953, 2153.133, 2208.673, 
    2052.604, 1710.461, 1339.997, 930.2275, 488.1713, 259.9942, 243.8892, 
    504.7442, 1907.184, 5704.826, 11677.85, 17820.93, 22301.88, 25433.91, 
    27589.06, 28428.74, 28356.5, 27455.85, 25012.35, 20863.42, 15971.65, 
    10754.41, 5644.089, 2049.034, 471.3907, 66.91194, 9.222707, 3.746444, 
    3.49807, 3.420794, 1.970172,
  0, 0.02292627, 0.3008365, 2.105643, 8.260301, 18.6011, 26.84878, 27.94549, 
    22.56685, 13.98377, 6.265257, 1.947727, 0.4289651, 0.07363721, 
    0.01007101, 0.0007674962, 0, 0.4501646, 5.907019, 45.31225, 200.1676, 
    512.1604, 845.0907, 1024.092, 999.4446, 776.0785, 457.8493, 220.5621, 
    100.2566, 40.29335, 21.84847, 45.1614, 104.0891, 192.6287, 320.2918, 
    494.3143, 694.3882, 867.5245, 957.2852, 972.2366, 985.1082, 1039.357, 
    1099.642, 1108.919, 1003.223, 726.6381, 381.5195, 155.6277, 73.68423, 
    50.92696, 37.77018, 23.06181, 13.9731, 18.38814, 35.14465, 54.37976, 
    62.60059, 53.94534, 36.60741, 22.46825, 13.49127, 6.785456, 2.42991, 
    0.5844054, 0.09024583, 0.007181752, 7.483396e-05, 5.70298e-06, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.01306407, 
    0.1714255, 2.890372, 23.55266, 102.6457, 277.2658, 507.2904, 689.1707, 
    771.919, 767.0975, 674.9398, 511.9892, 355.1158, 272.6285, 270.1862, 
    339.3355, 482.6144, 675.0828, 934.2108, 1414.033, 2090.372, 2591.64, 
    2658.125, 2240.125, 1445.477, 715.0067, 385.9046, 386.1033, 609.2662, 
    991.1838, 1550.458, 2838.724, 5700.763, 10134.67, 15136.56, 19670.09, 
    23151.14, 25460.41, 26724.78, 27079.77, 26617.79, 25424.19, 23536.96, 
    20727.86, 16820.81, 12113.76, 7314.173, 3434.925, 1177.738, 291.134, 
    55.10716, 7.952444, 0.6145499, 0.002092234, 0.0001594459,
  1.539552, 9.494467, 42.60406, 148.8519, 376.3348, 665.2653, 860.758, 
    881.8467, 749.0692, 517.6072, 280.5029, 120.743, 44.21815, 14.0353, 
    3.831038, 1.498572, 1.638375, 3.626983, 10.13899, 34.12737, 108.8737, 
    252.0609, 411.3943, 510.9113, 529.1339, 478.1214, 373.571, 245.5744, 
    129.7869, 51.46415, 16.65203, 12.29538, 23.10783, 44.38027, 80.38461, 
    143.5744, 253.932, 415.6334, 595.1274, 741.6502, 826.8279, 856.3439, 
    834.387, 733.4067, 538.4658, 306.8488, 129.4861, 41.48085, 13.22829, 
    6.84712, 4.771609, 3.005729, 2.249371, 3.808788, 7.566432, 11.51238, 
    12.91372, 10.76464, 6.984301, 4.087089, 2.463241, 1.348861, 0.5547107, 
    0.1568347, 0.028417, 0.002794967, 0.0001177264, 9.772384e-06, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0.002237674, 
    0.02695691, 0.473429, 4.500376, 23.79343, 74.83298, 152.5101, 222.448, 
    257.7247, 257.2993, 233.0039, 204.9987, 190.7024, 197.3507, 242.7679, 
    363.3904, 594.6749, 954.8204, 1434.409, 1994.828, 2584.181, 3140.48, 
    3497.938, 3341.577, 2614.877, 1843.768, 1574.511, 1944.784, 2968.304, 
    4532.467, 6465.117, 8932.212, 12021.14, 15182.64, 17920.14, 20446.65, 
    22888.96, 24731.47, 25613.2, 25648.73, 24958.96, 23711.5, 22051.05, 
    19658.27, 16159.69, 11764.12, 7216.296, 3529.223, 1343.757, 416.4416, 
    110.7744, 23.08969, 3.292629, 0.3950406, 0.1957537,
  5.213823, 26.20424, 102.6427, 308.7534, 689.1858, 1142.569, 1458.484, 
    1503.771, 1289.478, 915.4044, 529.4497, 252.5878, 104.8308, 39.44173, 
    13.77657, 6.355107, 7.440219, 13.67901, 23.33481, 33.94624, 44.18747, 
    55.09484, 70.73323, 101.7577, 159.6926, 230.6901, 267.3786, 234.2467, 
    151.1544, 70.40108, 23.36855, 6.115491, 2.898563, 6.113542, 20.59903, 
    61.18555, 143.9865, 274.1564, 435.5238, 585.6744, 674.1574, 672.032, 
    575.4656, 407.4914, 228.0344, 99.03681, 34.4919, 10.14694, 2.410491, 
    0.3920935, 0.04347607, 0.05639257, 0.246078, 0.706645, 1.401263, 2.01366, 
    2.142337, 1.707394, 1.063077, 0.5929514, 0.3539842, 0.2166755, 0.1131063, 
    0.04527956, 0.01314663, 0.002635191, 0.0003604439, 3.638089e-05, 
    2.420401e-06, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1.646813e-05, 0.0002475313, 0.006493859, 0.07983672, 0.5784287, 2.710253, 
    8.498638, 18.57947, 29.92297, 38.0874, 41.87165, 45.28305, 57.45543, 
    88.32388, 143.7047, 238.569, 413.6485, 713.0751, 1141.855, 1654.341, 
    2189.634, 2741.761, 3343.454, 3896.156, 4160.716, 4063.888, 3833.285, 
    3763.49, 4091.242, 5052.567, 6759.861, 9068.749, 11700.47, 14358.63, 
    16743.38, 18663.47, 20108.63, 21112.34, 21676.13, 21837.79, 21599.79, 
    20861.01, 19585.64, 17850.8, 15660.28, 12940.27, 9743.437, 6415.075, 
    3550.571, 1617.407, 611.0378, 195.9883, 53.60022, 12.28754, 2.403743, 
    1.085929,
  5.214683, 21.08001, 69.69033, 179.9967, 360.2772, 567.3036, 726.3879, 
    786.3427, 738.7462, 603.0378, 421.4787, 249.2514, 124.5554, 53.06929, 
    20.60192, 10.53441, 12.0768, 20.4143, 32.92693, 47.13588, 61.55175, 
    76.05445, 91.65887, 110.8155, 134.4909, 155.3025, 157.6989, 132.0477, 
    87.40575, 44.57181, 17.57524, 6.314337, 4.590349, 10.23435, 29.04996, 
    71.90106, 144.428, 235.5232, 318.2069, 363.6631, 354.1961, 291.0337, 
    198.0642, 110.3659, 50.68176, 19.68314, 6.68064, 2.015849, 0.5279037, 
    0.1102427, 0.01822097, 0.01360318, 0.0422155, 0.1026484, 0.184904, 
    0.2532462, 0.2677625, 0.2215791, 0.1483506, 0.0873197, 0.05089048, 
    0.03022827, 0.01656469, 0.007622583, 0.002849794, 0.0008647623, 
    0.0002117067, 3.970982e-05, 4.947156e-06, 2.928852e-07, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.664335e-07, 9.567691e-06, 
    0.0002398694, 0.00317127, 0.02526394, 0.1333581, 0.4879802, 1.284991, 
    2.532116, 3.900855, 4.958539, 5.669187, 7.038516, 12.35728, 29.81673, 
    76.80862, 182.4011, 379.4872, 686.0176, 1091.691, 1564.91, 2077.55, 
    2628.463, 3230.766, 3855.981, 4399.659, 4727.863, 4778.814, 4647.221, 
    4570.614, 4793.324, 5431.228, 6470.95, 7839.814, 9408.732, 10947.95, 
    12168.34, 12885.97, 13154.12, 13184.5, 13124.59, 12935.36, 12474.18, 
    11652.16, 10493.21, 9078.924, 7490.601, 5810.371, 4149.307, 2655.737, 
    1478.404, 695.6431, 271.1368, 87.28819, 23.66577, 5.63564, 2.021181,
  1.495067, 2.24579, 4.922228, 10.02801, 18.80852, 33.34372, 56.32339, 
    88.90589, 126.4694, 156.3481, 163.3904, 141.6704, 100.8215, 59.03258, 
    29.98407, 16.96084, 16.70107, 25.113, 39.22828, 56.62119, 74.86304, 
    91.2951, 102.7175, 105.5087, 97.06274, 78.21076, 54.18163, 32.01642, 
    16.34617, 7.659519, 4.025781, 3.743267, 7.108542, 17.38551, 40.25843, 
    79.58349, 130.068, 174.0665, 190.1693, 169.3202, 122.6453, 72.16795, 
    34.51572, 13.48118, 4.343651, 1.168371, 0.2636507, 0.04954094, 
    0.007635429, 0.0009338066, 8.136653e-05, 3.67264e-06, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3.085674e-07, 6.836244e-06, 
    9.244484e-05, 0.0009514221, 0.009025623, 0.08055032, 0.5926363, 3.338771, 
    14.31892, 47.62589, 125.9627, 272.3336, 496.4528, 791.024, 1147.585, 
    1578.437, 2116.75, 2781.491, 3528.607, 4232.202, 4720.301, 4846.326, 
    4557.482, 3930.029, 3150.718, 2441.845, 1968.141, 1783.769, 1843.01, 
    2052.464, 2330.575, 2644.672, 3001.466, 3395.558, 3764.387, 3999.748, 
    4007.715, 3762.333, 3317.293, 2778.571, 2254.513, 1806.879, 1433.821, 
    1098.474, 778.0626, 488.015, 262.2835, 118.2121, 44.12704, 13.60628, 
    3.657094,
  2.702178, 1.251308, 1.284701, 2.179508, 3.980809, 7.111449, 12.0729, 
    18.96877, 26.96257, 34.13276, 38.13166, 37.43576, 32.33397, 24.87972, 
    17.84955, 13.49838, 12.88296, 15.91025, 21.74875, 29.19403, 36.83191, 
    43.09019, 46.38872, 45.54792, 40.36107, 31.92462, 22.32023, 13.71361, 
    7.469125, 3.891431, 2.672643, 3.603363, 7.005666, 13.56108, 23.52724, 
    35.75586, 47.31322, 54.38022, 54.19434, 46.73166, 34.77337, 22.25749, 
    12.21423, 5.731743, 2.298985, 0.7911898, 0.2360549, 0.06206518, 
    0.01459717, 0.003070969, 0.0005655367, 8.804737e-05, 1.115496e-05, 
    1.090764e-06, 7.351246e-08, 2.530961e-09, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    2.12646e-10, 6.176361e-09, 1.012836e-07, 1.217211e-06, 1.341428e-05, 
    0.0001440908, 0.001355847, 0.0103037, 0.0621437, 0.3004976, 1.185, 
    3.87765, 10.70464, 25.3408, 52.3517, 96.34958, 161.9971, 256.0914, 
    390.7543, 583.4502, 849.0876, 1184.835, 1556.485, 1898.068, 2129.536, 
    2185.997, 2045.114, 1739.575, 1347.129, 960.7145, 653.186, 455.8252, 
    360.3786, 337.9569, 359.32, 405.2141, 465.3385, 531.5333, 592.2277, 
    632.4552, 639.1589, 607.796, 545.5119, 468.3992, 393.9854, 333.1616, 
    286.3933, 246.3806, 204.9067, 158.8608, 111.5796, 69.57468, 37.9509, 
    17.91308, 7.300492,
  0.01720216, 0.007134988, 0.002748055, 0.0009810849, 0.0003240056, 
    9.875001e-05, 2.769835e-05, 7.126376e-06, 1.67518e-06, 3.5806e-07, 
    6.918829e-08, 1.200131e-08, 1.85277e-09, 2.519483e-10, 2.980704e-11, 
    3.023391e-12, 2.584144e-13, 1.820687e-14, 1.022538e-15, 4.299969e-17, 
    1.203479e-18, 2.052644e-20, 4.119906e-22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5.27e-20, 2.625651e-18, 
    7.057653e-17, 1.346764e-15, 2.007508e-14, 2.444474e-13, 2.499678e-12, 
    2.19168e-11, 1.675506e-10, 1.13213e-09, 6.835349e-09, 3.7197e-08, 
    1.837231e-07, 8.283488e-07, 3.425768e-06, 1.305021e-05, 4.596037e-05, 
    0.0001501208, 0.0004560057, 0.001291075, 0.003413274, 0.008438042, 
    0.01952671, 0.04233364, 0.08603706, 0.1640046, 0.293362, 0.4926459, 
    0.7770787, 1.151924, 1.605646, 2.105614, 2.599134, 3.021201, 3.307919, 
    3.411966, 3.31508, 3.033181, 2.612199, 2.116059, 1.611047, 1.151707, 
    0.7723033, 0.4852658, 0.2853864, 0.1569097, 0.08055878, 0.03857289,
  0.0544402, 0.03951677, 0.02799566, 0.01935524, 0.01305729, 0.008594061, 
    0.00551794, 0.00345563, 0.002110497, 0.001256846, 0.0007297065, 
    0.0004129611, 0.000227765, 0.0001224055, 6.408632e-05, 3.268073e-05, 
    1.622884e-05, 7.846116e-06, 3.69226e-06, 1.690806e-06, 7.532645e-07, 
    3.263903e-07, 1.37512e-07, 5.631566e-08, 2.241138e-08, 8.663989e-09, 
    3.252582e-09, 1.185342e-09, 4.19179e-10, 1.43788e-10, 4.782231e-11, 
    1.541452e-11, 4.813012e-12, 1.455043e-12, 4.25675e-13, 1.204429e-13, 
    3.294035e-14, 8.702527e-15, 2.219433e-15, 5.460194e-16, 1.294831e-16, 
    2.95736e-17, 6.499856e-18, 1.373434e-18, 2.787295e-19, 5.427057e-20, 
    1.012632e-20, 1.808451e-21, 3.087086e-22, 5.029789e-23, 7.809636e-24, 
    1.153598e-24, 1.618154e-25, 2.151056e-26, 2.70392e-27, 3.206235e-28, 
    3.576841e-29, 3.745608e-30, 3.959941e-31, 3.434672e-31, 3.018101e-30, 
    2.749692e-29, 2.358987e-28, 1.909362e-27, 1.461746e-26, 1.060899e-25, 
    7.314778e-25, 4.800424e-24, 3.003764e-23, 1.794957e-22, 1.025848e-21, 
    5.61491e-21, 2.946989e-20, 1.484896e-19, 7.190601e-19, 3.349838e-18, 
    1.502727e-17, 6.497036e-17, 2.709483e-16, 1.090758e-15, 4.241841e-15, 
    1.594629e-14, 5.798569e-14, 2.040791e-13, 6.955651e-13, 2.297043e-12, 
    7.353758e-12, 2.2833e-11, 6.878951e-11, 2.011723e-10, 5.713091e-10, 
    1.576129e-09, 4.22553e-09, 1.101239e-08, 2.790793e-08, 6.879316e-08, 
    1.649886e-07, 3.850937e-07, 8.749615e-07, 1.935629e-06, 4.170241e-06, 
    8.751777e-06, 1.789422e-05, 3.565268e-05, 6.92327e-05, 0.000131052, 
    0.0002418571, 0.0004352345, 0.0007638368, 0.001307527, 0.002183391, 
    0.003557108, 0.005654572, 0.0087718, 0.01328039, 0.01962504, 0.02830932, 
    0.03986637, 0.0548124, 0.07358344, 0.09645882, 0.123479, 0.1543689, 
    0.1884802, 0.2247662, 0.2618024, 0.2978575, 0.331015, 0.3593354, 
    0.3810408, 0.394698, 0.3993745, 0.3947428, 0.3811187, 0.3594256, 
    0.3310912, 0.2978932, 0.2617753, 0.2246623, 0.1882955, 0.1541096, 
    0.1231596, 0.09609957, 0.0732069,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 lat = -90, -88.1052631578947, -86.2105263157895, -84.3157894736842, 
    -82.4210526315789, -80.5263157894737, -78.6315789473684, 
    -76.7368421052632, -74.8421052631579, -72.9473684210526, 
    -71.0526315789474, -69.1578947368421, -67.2631578947368, 
    -65.3684210526316, -63.4736842105263, -61.578947368421, 
    -59.6842105263158, -57.7894736842105, -55.8947368421053, -54, 
    -52.1052631578947, -50.2105263157895, -48.3157894736842, 
    -46.421052631579, -44.5263157894737, -42.6315789473684, 
    -40.7368421052632, -38.8421052631579, -36.9473684210526, 
    -35.0526315789474, -33.1578947368421, -31.2631578947368, 
    -29.3684210526316, -27.4736842105263, -25.5789473684211, 
    -23.6842105263158, -21.7894736842105, -19.8947368421053, -18, 
    -16.1052631578947, -14.2105263157895, -12.3157894736842, 
    -10.421052631579, -8.52631578947369, -6.63157894736843, 
    -4.73684210526316, -2.8421052631579, -0.947368421052636, 
    0.947368421052627, 2.84210526315789, 4.73684210526315, 6.63157894736842, 
    8.52631578947368, 10.4210526315789, 12.3157894736842, 14.2105263157895, 
    16.1052631578947, 18, 19.8947368421053, 21.7894736842105, 
    23.6842105263158, 25.578947368421, 27.4736842105263, 29.3684210526316, 
    31.2631578947368, 33.1578947368421, 35.0526315789474, 36.9473684210526, 
    38.8421052631579, 40.7368421052632, 42.6315789473684, 44.5263157894737, 
    46.4210526315789, 48.3157894736842, 50.2105263157895, 52.1052631578947, 
    54, 55.8947368421053, 57.7894736842105, 59.6842105263158, 
    61.578947368421, 63.4736842105263, 65.3684210526316, 67.2631578947368, 
    69.1578947368421, 71.0526315789474, 72.9473684210526, 74.8421052631579, 
    76.7368421052632, 78.6315789473684, 80.5263157894737, 82.4210526315789, 
    84.3157894736842, 86.2105263157895, 88.1052631578947, 90 ;

 lon = 0, 2.5, 5, 7.5, 10, 12.5, 15, 17.5, 20, 22.5, 25, 27.5, 30, 32.5, 35, 
    37.5, 40, 42.5, 45, 47.5, 50, 52.5, 55, 57.5, 60, 62.5, 65, 67.5, 70, 
    72.5, 75, 77.5, 80, 82.5, 85, 87.5, 90, 92.5, 95, 97.5, 100, 102.5, 105, 
    107.5, 110, 112.5, 115, 117.5, 120, 122.5, 125, 127.5, 130, 132.5, 135, 
    137.5, 140, 142.5, 145, 147.5, 150, 152.5, 155, 157.5, 160, 162.5, 165, 
    167.5, 170, 172.5, 175, 177.5, 180, 182.5, 185, 187.5, 190, 192.5, 195, 
    197.5, 200, 202.5, 205, 207.5, 210, 212.5, 215, 217.5, 220, 222.5, 225, 
    227.5, 230, 232.5, 235, 237.5, 240, 242.5, 245, 247.5, 250, 252.5, 255, 
    257.5, 260, 262.5, 265, 267.5, 270, 272.5, 275, 277.5, 280, 282.5, 285, 
    287.5, 290, 292.5, 295, 297.5, 300, 302.5, 305, 307.5, 310, 312.5, 315, 
    317.5, 320, 322.5, 325, 327.5, 330, 332.5, 335, 337.5, 340, 342.5, 345, 
    347.5, 350, 352.5, 355, 357.5 ;

 time = 0 ;
}
