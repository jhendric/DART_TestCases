netcdf wc13_ecco_bry {
dimensions:
	xi_rho = 56 ;
	eta_rho = 55 ;
	xi_u = 55 ;
	eta_u = 55 ;
	xi_v = 56 ;
	eta_v = 54 ;
	s_rho = 30 ;
	s_w = 31 ;
	zeta_time = 2 ;
	v2d_time = 2 ;
	v3d_time = 2 ;
	temp_time = 2 ;
	salt_time = 2 ;
variables:
	int spherical ;
		spherical:long_name = "grid type logical switch" ;
		spherical:flag_values = 0, 1 ;
		spherical:flag_meanings = "Cartesian spherical" ;
	int Vtransform ;
		Vtransform:long_name = "vertical terrain-following transformation equation" ;
	int Vstretching ;
		Vstretching:long_name = "vertical terrain-following stretching function" ;
	double theta_s ;
		theta_s:long_name = "S-coordinate surface control parameter" ;
	double theta_b ;
		theta_b:long_name = "S-coordinate bottom control parameter" ;
	double Tcline ;
		Tcline:long_name = "S-coordinate surface/bottom layer width" ;
		Tcline:units = "meter" ;
	double hc ;
		hc:long_name = "S-coordinate parameter, critical depth" ;
		hc:units = "meter" ;
	double s_rho(s_rho) ;
		s_rho:long_name = "S-coordinate at RHO-points" ;
		s_rho:valid_min = -1. ;
		s_rho:valid_max = 0. ;
		s_rho:positive = "up" ;
		s_rho:standard_name = "ocean_s_coordinate_g1" ;
		s_rho:formula_terms = "s: s_rho C: Cs_r eta: zeta depth: h depth_c: hc" ;
	double s_w(s_w) ;
		s_w:long_name = "S-coordinate at W-points" ;
		s_w:valid_min = -1. ;
		s_w:valid_max = 0. ;
		s_w:positive = "up" ;
		s_w:standard_name = "ocean_s_coordinate_g1" ;
		s_w:formula_terms = "s: s_w C: Cs_w eta: zeta depth: h depth_c: hc" ;
	double Cs_r(s_rho) ;
		Cs_r:long_name = "S-coordinate stretching curves at RHO-points" ;
		Cs_r:valid_min = -1. ;
		Cs_r:valid_max = 0. ;
	double Cs_w(s_w) ;
		Cs_w:long_name = "S-coordinate stretching curves at W-points" ;
		Cs_w:valid_min = -1. ;
		Cs_w:valid_max = 0. ;
	double h(eta_rho, xi_rho) ;
		h:long_name = "bathymetry at RHO-points" ;
		h:units = "meter" ;
		h:coordinates = "lon_rho lat_rho" ;
	double lon_rho(eta_rho, xi_rho) ;
		lon_rho:long_name = "longitude of RHO-points" ;
		lon_rho:units = "degree_east" ;
		lon_rho:standard_name = "longitude" ;
	double lat_rho(eta_rho, xi_rho) ;
		lat_rho:long_name = "latitude of RHO-points" ;
		lat_rho:units = "degree_north" ;
		lat_rho:standard_name = "latitude" ;
	double lon_u(eta_u, xi_u) ;
		lon_u:long_name = "longitude of U-points" ;
		lon_u:units = "degree_east" ;
		lon_u:standard_name = "longitude" ;
	double lat_u(eta_u, xi_u) ;
		lat_u:long_name = "latitude of U-points" ;
		lat_u:units = "degree_north" ;
		lat_u:standard_name = "latitude" ;
	double lon_v(eta_v, xi_v) ;
		lon_v:long_name = "longitude of V-points" ;
		lon_v:units = "degree_east" ;
		lon_v:standard_name = "longitude" ;
	double lat_v(eta_v, xi_v) ;
		lat_v:long_name = "latitude of V-points" ;
		lat_v:units = "degree_north" ;
		lat_v:standard_name = "latitude" ;
	double zeta_time(zeta_time) ;
		zeta_time:long_name = "free-surface time" ;
		zeta_time:units = "seconds since 1968-05-23 00:00:00 GMT" ;
		zeta_time:calendar = "gregorian" ;
	double v2d_time(v2d_time) ;
		v2d_time:long_name = "2D momentum time" ;
		v2d_time:units = "seconds since 1968-05-23 00:00:00 GMT" ;
		v2d_time:calendar = "gregorian" ;
	double v3d_time(v3d_time) ;
		v3d_time:long_name = "3D momentum time" ;
		v3d_time:units = "seconds since 1968-05-23 00:00:00 GMT" ;
		v3d_time:calendar = "gregorian" ;
	double temp_time(temp_time) ;
		temp_time:long_name = "potential temperature time" ;
		temp_time:units = "seconds since 1968-05-23 00:00:00 GMT" ;
		temp_time:calendar = "gregorian" ;
	double salt_time(salt_time) ;
		salt_time:long_name = "surface net heat flux time" ;
		salt_time:units = "seconds since 1968-05-23 00:00:00 GMT" ;
		salt_time:calendar = "gregorian" ;
	float zeta_west(zeta_time, eta_rho) ;
		zeta_west:long_name = "free-surface western boundary condition" ;
		zeta_west:units = "meter" ;
		zeta_west:time = "zeta_time" ;
	float zeta_east(zeta_time, eta_rho) ;
		zeta_east:long_name = "free-surface eastern boundary condition" ;
		zeta_east:units = "meter" ;
		zeta_east:time = "zeta_time" ;
	float zeta_south(zeta_time, xi_rho) ;
		zeta_south:long_name = "free-surface southern boundary condition" ;
		zeta_south:units = "meter" ;
		zeta_south:time = "zeta_time" ;
	float zeta_north(zeta_time, xi_rho) ;
		zeta_north:long_name = "free-surface northern boundary condition" ;
		zeta_north:units = "meter" ;
		zeta_north:time = "zeta_time" ;
	float ubar_west(v2d_time, eta_u) ;
		ubar_west:long_name = "2D u-momentum western boundary condition" ;
		ubar_west:units = "meter second-1" ;
		ubar_west:time = "v2d_time" ;
	float ubar_east(v2d_time, eta_u) ;
		ubar_east:long_name = "2D u-momentum eastern boundary condition" ;
		ubar_east:units = "meter second-1" ;
		ubar_east:time = "v2d_time" ;
	float ubar_south(v2d_time, xi_u) ;
		ubar_south:long_name = "2D u-momentum southern boundary condition" ;
		ubar_south:units = "meter second-1" ;
		ubar_south:time = "v2d_time" ;
	float ubar_north(v2d_time, xi_u) ;
		ubar_north:long_name = "2D u-momentum northern boundary condition" ;
		ubar_north:units = "meter second-1" ;
		ubar_north:time = "v2d_time" ;
	float vbar_west(v2d_time, eta_v) ;
		vbar_west:long_name = "2D v-momentum western boundary condition" ;
		vbar_west:units = "meter second-1" ;
		vbar_west:time = "v2d_time" ;
	float vbar_east(v2d_time, eta_v) ;
		vbar_east:long_name = "2D v-momentum eastern boundary condition" ;
		vbar_east:units = "meter second-1" ;
		vbar_east:time = "v2d_time" ;
	float vbar_south(v2d_time, xi_v) ;
		vbar_south:long_name = "2D v-momentum southern boundary condition" ;
		vbar_south:units = "meter second-1" ;
		vbar_south:time = "v2d_time" ;
	float vbar_north(v2d_time, xi_v) ;
		vbar_north:long_name = "2D v-momentum northern boundary condition" ;
		vbar_north:units = "meter second-1" ;
		vbar_north:time = "v2d_time" ;
	float u_west(v3d_time, s_rho, eta_u) ;
		u_west:long_name = "3D u-momentum western boundary condition" ;
		u_west:units = "meter second-1" ;
		u_west:time = "v3d_time" ;
	float u_east(v3d_time, s_rho, eta_u) ;
		u_east:long_name = "3D u-momentum eastern boundary condition" ;
		u_east:units = "meter second-1" ;
		u_east:time = "v3d_time" ;
	float u_south(v3d_time, s_rho, xi_u) ;
		u_south:long_name = "3D u-momentum southern boundary condition" ;
		u_south:units = "meter second-1" ;
		u_south:time = "v3d_time" ;
	float u_north(v3d_time, s_rho, xi_u) ;
		u_north:long_name = "3D u-momentum northern boundary condition" ;
		u_north:units = "meter second-1" ;
		u_north:time = "v3d_time" ;
	float v_west(v3d_time, s_rho, eta_v) ;
		v_west:long_name = "3D v-momentum western boundary condition" ;
		v_west:units = "meter second-1" ;
		v_west:time = "v3d_time" ;
	float v_east(v3d_time, s_rho, eta_v) ;
		v_east:long_name = "3D v-momentum eastern boundary condition" ;
		v_east:units = "meter second-1" ;
		v_east:time = "v3d_time" ;
	float v_south(v3d_time, s_rho, xi_v) ;
		v_south:long_name = "3D v-momentum southern boundary condition" ;
		v_south:units = "meter second-1" ;
		v_south:time = "v3d_time" ;
	float v_north(v3d_time, s_rho, xi_v) ;
		v_north:long_name = "3D v-momentum northern boundary condition" ;
		v_north:units = "meter second-1" ;
		v_north:time = "v3d_time" ;
	float temp_west(temp_time, s_rho, eta_rho) ;
		temp_west:long_name = "potential temperature western boundary condition" ;
		temp_west:units = "Celsius" ;
		temp_west:time = "temp_time" ;
	float temp_east(temp_time, s_rho, eta_rho) ;
		temp_east:long_name = "potential temperature eastern boundary condition" ;
		temp_east:units = "Celsius" ;
		temp_east:time = "temp_time" ;
	float temp_south(temp_time, s_rho, xi_rho) ;
		temp_south:long_name = "potential temperature southern boundary condition" ;
		temp_south:units = "Celsius" ;
		temp_south:time = "temp_time" ;
	float temp_north(temp_time, s_rho, xi_rho) ;
		temp_north:long_name = "potential temperature northern boundary condition" ;
		temp_north:units = "Celsius" ;
		temp_north:time = "temp_time" ;
	float salt_west(salt_time, s_rho, eta_rho) ;
		salt_west:long_name = "salinity western boundary condition" ;
		salt_west:time = "salt_time" ;
	float salt_east(salt_time, s_rho, eta_rho) ;
		salt_east:long_name = "salinity eastern boundary condition" ;
		salt_east:time = "salt_time" ;
	float salt_south(salt_time, s_rho, xi_rho) ;
		salt_south:long_name = "salinity southern boundary condition" ;
		salt_south:time = "salt_time" ;
	float salt_north(salt_time, s_rho, xi_rho) ;
		salt_north:long_name = "salinity northern boundary condition" ;
		salt_north:time = "salt_time" ;

// global attributes:
		:type = "BOUNDARY FORCING" ;
		:Conventions = "CF-1.4" ;
		:title = "California Current System, 1/3 degree resolution (WC13)" ;
		:grd_file = "wc13_grd.nc" ;
		:history = "Thursday - February 8, 2007 -  11:00:00 AM" ;
data:

 spherical = 1 ;

 Vtransform = 1 ;

 Vstretching = 1 ;

 theta_s = 5 ;

 theta_b = 0.4 ;

 Tcline = 10 ;

 hc = 10 ;

 s_rho = -0.983333333333333, -0.95, -0.916666666666667, -0.883333333333333, 
    -0.85, -0.816666666666667, -0.783333333333333, -0.75, -0.716666666666667, 
    -0.683333333333333, -0.65, -0.616666666666667, -0.583333333333333, -0.55, 
    -0.516666666666667, -0.483333333333333, -0.45, -0.416666666666667, 
    -0.383333333333333, -0.35, -0.316666666666667, -0.283333333333333, -0.25, 
    -0.216666666666667, -0.183333333333333, -0.15, -0.116666666666667, 
    -0.0833333333333333, -0.05, -0.0166666666666667 ;

 s_w = -1, -0.966666666666667, -0.933333333333333, -0.9, -0.866666666666667, 
    -0.833333333333333, -0.8, -0.766666666666667, -0.733333333333333, -0.7, 
    -0.666666666666667, -0.633333333333333, -0.6, -0.566666666666667, 
    -0.533333333333333, -0.5, -0.466666666666667, -0.433333333333333, -0.4, 
    -0.366666666666667, -0.333333333333333, -0.3, -0.266666666666667, 
    -0.233333333333333, -0.2, -0.166666666666667, -0.133333333333333, -0.1, 
    -0.0666666666666667, -0.0333333333333333, 0 ;

 Cs_r = -0.951533875009937, -0.865525766528738, -0.792044761269449, 
    -0.728914353094819, -0.674204624279983, -0.626170729989037, 
    -0.583200287133593, -0.543774115119252, -0.506448977195438, 
    -0.469875433493012, -0.432865580628998, -0.39451827877102, 
    -0.354386434772583, -0.312632258634705, -0.270082002827858, 
    -0.228100664712844, -0.188284024260942, -0.15207318852824, 
    -0.1204487484324, -0.0938097782858442, -0.0720351699264823, 
    -0.0546479652981894, -0.0409944497135269, -0.0303842518734395, 
    -0.022176433349889, -0.0158196793238963, -0.0108619873876149, 
    -0.00694371576956987, -0.00378353920774699, -0.00116283376462356 ;

 Cs_w = -1, -0.9068164336607, -0.827361959419869, -0.759311373494851, 
    -0.700619627249543, -0.649456534986167, -0.604149373019713, 
    -0.563136150071506, -0.524935972281481, -0.488147475821263, 
    -0.451489928129714, -0.41389976586145, -0.374680938702067, 
    -0.333675595048554, -0.291381088924103, -0.248921369578993, 
    -0.207823725744927, -0.169653369247619, -0.135649074479394, 
    -0.106503119630948, -0.0823381033977505, -0.0628317602307056, 
    -0.0473980529834848, -0.0353508120779761, -0.026016827357272, 
    -0.0187972226760524, -0.0131904457723761, -0.00879215816914654, 
    -0.00528382012336189, -0.00241737715547015, -2.22044604925031e-17 ;

 h =
  4544.23173916444, 4544.23173916444, 4544.79426389874, 4575.27187875418, 
    4627.88387506815, 4656.53924392246, 4631.08347903984, 4577.49706734492, 
    4552.47814461172, 4565.54221912462, 4586.18364719751, 4594.30447609547, 
    4574.39206650845, 4527.69684711849, 4495.83801948936, 4492.14709328146, 
    4467.64380074904, 4399.44136055673, 4327.49472148068, 4302.29688279779, 
    4320.35897876608, 4343.08814634039, 4358.20738541416, 4349.46475029001, 
    4289.75441283314, 4215.81804710384, 4185.22222271129, 4187.05275653615, 
    4189.38818301993, 4186.4490169725, 4175.66341773197, 4142.07739985843, 
    4075.70044918496, 3997.00312800151, 3944.25371901054, 3935.16549206096, 
    3951.2558047985, 3958.64548793587, 3943.45989706591, 3911.34708277734, 
    3862.1715666883, 3780.79737664238, 3678.11557646457, 3595.67176022016, 
    3501.49492621635, 3289.25979329267, 2896.58205795875, 2352.40586806033, 
    1772.09928153261, 1302.56677967285, 960.976870860982, 711.196259578647, 
    522.555355162128, 395.323088498131, 323.662451586529, 323.662451586529,
  4544.23173916444, 4544.23173916444, 4544.79426389874, 4575.27187875418, 
    4627.88387506815, 4656.53924392246, 4631.08347903984, 4577.49706734492, 
    4552.47814461172, 4565.54221912462, 4586.18364719751, 4594.30447609547, 
    4574.39206650845, 4527.69684711849, 4495.83801948936, 4492.14709328146, 
    4467.64380074904, 4399.44136055673, 4327.49472148068, 4302.29688279779, 
    4320.35897876608, 4343.08814634039, 4358.20738541416, 4349.46475029001, 
    4289.75441283314, 4215.81804710384, 4185.22222271129, 4187.05275653615, 
    4189.38818301993, 4186.4490169725, 4175.66341773197, 4142.07739985843, 
    4075.70044918496, 3997.00312800151, 3944.25371901054, 3935.16549206096, 
    3951.2558047985, 3958.64548793587, 3943.45989706591, 3911.34708277734, 
    3862.1715666883, 3780.79737664238, 3678.11557646457, 3595.67176022016, 
    3501.49492621635, 3289.25979329267, 2896.58205795875, 2352.40586806033, 
    1772.09928153261, 1302.56677967285, 960.976870860982, 711.196259578647, 
    522.555355162128, 395.323088498131, 323.662451586529, 323.662451586529,
  4581.20306850219, 4581.20306850219, 4581.05443610493, 4604.71946120312, 
    4646.54670934288, 4668.91718302023, 4642.97795096356, 4589.43046853591, 
    4562.31846514785, 4574.72143430655, 4598.07616632174, 4608.02692384179, 
    4587.5322195804, 4538.40625260849, 4498.02567931232, 4481.39651749719, 
    4448.80703087107, 4375.58943533342, 4294.01949303288, 4259.57370812034, 
    4280.9909609781, 4321.60253935474, 4357.0287159001, 4362.45089786222, 
    4311.35787693119, 4235.03204846224, 4189.87261251325, 4180.88537292758, 
    4180.97041782351, 4171.26804870582, 4146.13681235275, 4103.17921234677, 
    4046.36081877392, 3997.51670687154, 3978.95990758941, 3987.28481777666, 
    3999.29846022342, 3992.84820420204, 3963.40744799293, 3922.91335533047, 
    3878.55474333038, 3809.91438417508, 3702.02941591236, 3569.16450006744, 
    3373.21026382655, 3037.25614865833, 2559.08504641728, 2018.77701672062, 
    1508.65439707269, 1101.85843894156, 804.857064242746, 589.420523815565, 
    432.405454431678, 327.867105788503, 270.561290302579, 270.561290302579,
  4623.48833534044, 4623.48833534044, 4625.14308297671, 4638.80853527542, 
    4659.10093049708, 4664.876579305, 4636.29923315107, 4586.95346909775, 
    4559.88098009503, 4569.42963393316, 4592.64138892843, 4602.2119480859, 
    4578.84784914869, 4525.46862983985, 4475.64605906825, 4446.28825789006, 
    4409.6961336633, 4343.22514035204, 4268.75493274308, 4235.30178810939, 
    4256.20727567624, 4300.30483051158, 4341.06981543873, 4355.63545056018, 
    4320.84189534038, 4250.86150468709, 4189.93962693495, 4165.34013134978, 
    4163.87865036288, 4153.10365452407, 4121.53069379165, 4078.59485956991, 
    4038.31985303755, 4014.94129633134, 4013.96482627076, 4024.25773046066, 
    4026.96701675567, 4008.19534275141, 3968.61092777677, 3925.89555819141, 
    3889.10678853173, 3815.03229319934, 3652.32423194131, 3403.83859850201, 
    3048.63099772166, 2567.14694332822, 2033.12121939942, 1549.58325861452, 
    1149.410358201, 833.849817994801, 605.111913755601, 441.745291281403, 
    325.709794087748, 248.1380027957, 206.709043091792, 206.709043091792,
  4652.49641856838, 4652.49641856838, 4658.5461386928, 4662.93531597116, 
    4657.56341975582, 4640.42860451954, 4608.81642327584, 4571.97481931722, 
    4553.27888378034, 4559.03073255249, 4572.42395869682, 4572.33661759364, 
    4543.54532272951, 4489.45676601025, 4436.98801095366, 4401.77185089924, 
    4368.26614983131, 4322.03878856609, 4275.39563775351, 4255.77206939713, 
    4262.12073770524, 4270.89520606311, 4282.30934941684, 4297.82260378007, 
    4292.73002600475, 4249.92511298711, 4190.16411093688, 4155.80925090521, 
    4152.98117612948, 4148.64273940564, 4127.72165322691, 4101.17960632973, 
    4079.27211849663, 4060.8538276248, 4043.02344561869, 4027.71648229933, 
    4011.3481185846, 3983.18480503743, 3942.4715340666, 3901.76154164396, 
    3843.27458580368, 3685.46003687713, 3384.03405107853, 2990.73822956482, 
    2524.82272759487, 2005.92978069869, 1524.47099468206, 1144.66824908798, 
    846.049317940853, 610.484254076365, 442.456197990811, 323.9578135515, 
    239.886940147896, 183.087521960577, 152.880194252125, 152.880194252125,
  4659.13365936528, 4659.13365936528, 4675.43398069902, 4680.91745536224, 
    4657.66545888755, 4616.97801431754, 4579.62166961895, 4558.72163052341, 
    4554.67947359429, 4557.09097731079, 4553.84507677578, 4538.80438734522, 
    4508.69910722481, 4464.94124411728, 4419.78874711566, 4383.70059947938, 
    4352.531597622, 4315.71217121884, 4279.26319547345, 4264.80249812204, 
    4255.28910969561, 4220.77925907525, 4195.4200373486, 4215.46374165356, 
    4250.20252577742, 4251.82402282647, 4217.24173710575, 4186.55755234997, 
    4179.09714390133, 4176.52566650864, 4167.57510472287, 4157.86750123282, 
    4149.69353671237, 4132.89991472317, 4099.23465982375, 4054.36492033476, 
    4005.39597026007, 3953.25007095246, 3898.19546619301, 3821.44278441447, 
    3651.28505169201, 3311.16691219192, 2843.15538265381, 2362.62555133848, 
    1901.79030526253, 1465.89892099186, 1101.2866479768, 824.843822806377, 
    606.941334723719, 439.458989396382, 321.98879850632, 237.517464793998, 
    175.947038438146, 133.294688359389, 109.884937990091, 109.884937990091,
  4647.63529134803, 4647.63529134803, 4681.35148584362, 4700.55364451643, 
    4670.25970768922, 4607.61855649259, 4555.94730699649, 4536.8265102513, 
    4534.06571154281, 4527.24178105183, 4512.46491043904, 4493.88426033577, 
    4472.97585543645, 4447.24280229628, 4417.65876141512, 4390.84235993417, 
    4361.44573105093, 4301.58012341757, 4221.80030742787, 4191.51282768478, 
    4205.43577850412, 4193.82916410683, 4175.47459867039, 4202.14147844874, 
    4254.5132421351, 4285.25796122482, 4279.75955338952, 4259.27367699597, 
    4243.37739999847, 4232.64894977857, 4222.03372015607, 4211.33917252256, 
    4202.71346119134, 4190.03262671499, 4159.8625352122, 4102.99413920884, 
    4023.22836404036, 3932.55425236281, 3817.39975844179, 3612.52282600939, 
    3244.67739026829, 2734.00318511326, 2202.4614281815, 1747.57433009297, 
    1370.64878144944, 1048.11980560431, 787.951232380888, 587.759925055099, 
    429.667825556643, 313.14237482486, 231.94229675481, 171.8256163584, 
    126.946473875121, 94.7817862435477, 76.6650168625554, 76.6650168625554,
  4637.68969497669, 4637.68969497669, 4677.52803120923, 4692.73412900199, 
    4651.63967498131, 4588.19028259844, 4539.38068468956, 4510.11573477237, 
    4485.20928962466, 4459.68061337293, 4441.86485429655, 4433.39421457502, 
    4428.37308665449, 4421.83206469579, 4413.81411909414, 4407.98611895634, 
    4385.720936857, 4296.76810484593, 4163.08967015618, 4112.91227510697, 
    4170.96318975353, 4229.84071062217, 4255.28755154373, 4284.0517524371, 
    4322.53333122122, 4353.06468929402, 4361.85029231426, 4346.32875071427, 
    4319.39222334353, 4295.89375871934, 4272.12995894136, 4243.75772320817, 
    4220.99251678725, 4205.55370015074, 4180.28050399216, 4124.31391812456, 
    4029.62070005339, 3884.35765879391, 3627.65277117482, 3210.64769654756, 
    2666.51653057594, 2111.10050803224, 1636.34089602099, 1268.69199028966, 
    984.177998675156, 750.852294306836, 564.164699106238, 418.910247037904, 
    305.411496577657, 223.314271548412, 165.078777990805, 121.594604096877, 
    89.4592573763288, 66.1016868210483, 52.9644744472566, 52.9644744472566,
  4655.11660036142, 4655.11660036142, 4670.71017112609, 4640.2033972255, 
    4578.48435599508, 4555.73206062764, 4556.74475142744, 4528.66197025972, 
    4476.18024170199, 4431.52143962979, 4410.04166580416, 4406.15450279078, 
    4410.44737587045, 4419.12953263844, 4430.91037105882, 4442.69928865785, 
    4433.08713903214, 4359.98417850935, 4243.02753461369, 4191.54003458094, 
    4238.09651438767, 4302.58231814134, 4341.70731665728, 4368.51072827602, 
    4394.65775758866, 4421.48649514877, 4436.78299307274, 4420.79392651344, 
    4382.48971757325, 4347.61675794033, 4311.86659266128, 4267.78157218745, 
    4230.98244048305, 4203.45544599825, 4165.04368089032, 4095.17624398876, 
    3969.78509514393, 3721.36659555542, 3260.14276258651, 2660.39777091905, 
    2062.90760035477, 1572.30440162224, 1194.1278121366, 912.869622010108, 
    700.487004202836, 529.815402810136, 394.779509869509, 291.559155614352, 
    213.270111252041, 156.945280733921, 115.840190262992, 84.9505239394382, 
    62.5787481068954, 46.5053157320914, 37.6536739418347, 37.6536739418347,
  4722.17499895874, 4722.17499895874, 4711.72505206442, 4648.95236897551, 
    4589.95841975627, 4618.0849854606, 4665.92878030228, 4640.80534759011, 
    4573.59132227387, 4521.43144949398, 4494.05507496239, 4481.67958954755, 
    4478.87686643682, 4483.87423316343, 4493.58353364064, 4502.37703498201, 
    4499.81523266211, 4469.49207647492, 4413.90362619637, 4370.18203777397, 
    4358.29582978939, 4364.60689649414, 4379.85412032965, 4401.33306252238, 
    4426.24355326677, 4456.31380503157, 4479.31480120011, 4466.27910799341, 
    4421.69480901602, 4377.66805770294, 4336.62967611443, 4290.87854499481, 
    4249.24786919094, 4205.62996030446, 4129.87435582875, 3989.11344011646, 
    3749.44565231115, 3333.71377326732, 2707.39215845518, 2066.84332325927, 
    1533.4063370843, 1137.51387586013, 846.518820470319, 638.219763078127, 
    484.524898946922, 364.86949581633, 271.047325791245, 200.655914745441, 
    148.528742712036, 110.450993728711, 81.8217421229109, 60.0664150976212, 
    44.39150007444, 33.2283846328971, 27.1455914382647, 27.1455914382647,
  4839.197637147, 4839.197637147, 4833.20613518488, 4801.29393291243, 
    4785.08356147458, 4828.43249278775, 4863.26510967357, 4826.50193817306, 
    4762.91104655535, 4717.54642191982, 4686.17511130547, 4659.47704694789, 
    4634.40152762302, 4609.6371402811, 4590.58506774037, 4580.92455758778, 
    4574.48352202061, 4561.09053613555, 4531.59048054844, 4486.21162143848, 
    4439.53578308103, 4411.6966868979, 4410.32633597315, 4425.42114582258, 
    4445.71469973072, 4472.81246759508, 4498.17248118439, 4490.88682500138, 
    4445.49244773682, 4391.73051521803, 4348.32178645424, 4312.30383890512, 
    4271.68361300608, 4199.60689726054, 4039.12679141241, 3734.62510038382, 
    3291.31385317629, 2719.9800418162, 2076.29148568086, 1541.85372600583, 
    1130.96582493334, 822.176542462913, 596.974285161318, 442.382119308157, 
    331.452595963358, 249.050390407283, 185.464703758093, 138.466926437112, 
    104.011387437909, 78.0292501844521, 57.9614899389249, 42.6572007825565, 
    31.6454058609897, 23.8642346370132, 19.6604871852787, 19.6604871852787,
  4970.66419408737, 4970.66419408737, 4975.1587636182, 4982.44464757379, 
    5001.46833408445, 5030.23970843441, 5031.67364608269, 4992.92680239878, 
    4950.01298633855, 4916.42676778564, 4878.37902257174, 4834.80398179935, 
    4785.1867957837, 4728.50368077253, 4684.44128994845, 4666.14613894863, 
    4657.02876733997, 4638.94145816627, 4606.57786254995, 4561.77123589576, 
    4515.78390701885, 4486.13536541385, 4482.40245163123, 4496.40249647202, 
    4511.83478368329, 4526.04849492881, 4536.66631291294, 4522.4078719028, 
    4471.49269377475, 4405.39131088651, 4358.63802729304, 4333.11171033397, 
    4282.7337667682, 4139.38324482518, 3822.40794773347, 3297.5027851464, 
    2669.50595564834, 2052.3693377238, 1518.54720504216, 1127.47844918619, 
    828.075997332773, 594.219763613423, 421.987403819266, 307.341369845669, 
    227.067799567441, 169.488750048895, 126.464245699632, 95.4213355999122, 
    72.5806101206411, 54.8664994530235, 41.0314297053813, 30.5919710750778, 
    22.9923757922265, 17.5226730036082, 14.563966661654, 14.563966661654,
  5071.78968633837, 5071.78968633837, 5071.26768457787, 5078.95756132154, 
    5095.01037700239, 5107.42625091151, 5101.81445138946, 5081.97710501549, 
    5062.2563244778, 5032.71694318789, 4981.12649542033, 4922.90080226929, 
    4863.73787752757, 4799.57683135895, 4755.19735635622, 4744.04211661822, 
    4738.10320181809, 4719.04868696445, 4693.05417092001, 4663.40329183095, 
    4629.08626498677, 4598.70044222693, 4589.27088805911, 4601.03343159064, 
    4611.5360000834, 4607.68492192521, 4590.25656654651, 4553.51533591393, 
    4489.10246928203, 4411.32751206983, 4358.95876454559, 4328.21443151194, 
    4230.21445944968, 3955.78039263282, 3449.26310649583, 2755.11619613271, 
    2062.23614660648, 1501.13286080552, 1092.34349880951, 802.92410049247, 
    583.348716844789, 416.747059981793, 293.335353246967, 210.128482888655, 
    153.07836771147, 114.019792684054, 85.7988988319871, 65.5563766715868, 
    50.425537292467, 38.585086499834, 29.2690563082526, 22.250764294712, 
    17.1184670858479, 13.5187279623415, 11.6699447476716, 11.6699447476716,
  5123.6037491913, 5123.6037491913, 5114.98082386404, 5108.13546112219, 
    5107.43143459747, 5111.18561269296, 5113.94560251188, 5113.12016054178, 
    5103.95373683565, 5066.9858340723, 4999.25517723011, 4934.34500773128, 
    4884.41875751488, 4836.32584331279, 4805.14664663132, 4800.43567708298, 
    4796.05471248216, 4781.55536295418, 4769.2285492328, 4758.08073197528, 
    4736.05652541613, 4704.18424551834, 4682.35257080251, 4678.71262119273, 
    4674.20509152265, 4651.44770526897, 4609.10376095326, 4549.97174305126, 
    4472.46334737095, 4387.23521323761, 4323.09654640801, 4252.33889775095, 
    4044.2089370089, 3591.15778156123, 2934.65519077142, 2200.04145574465, 
    1568.09496054666, 1107.79128336172, 790.433250015548, 566.679079229781, 
    404.088477087324, 289.051310596887, 204.766845173323, 145.25349312548, 
    104.341975527756, 77.452359634942, 58.7784672768897, 45.5126595684195, 
    35.4903783850075, 27.5711601191515, 21.2350821651204, 16.4750942128851, 
    13.1996423965538, 11.2415790576685, 10.409478761505, 10.409478761505,
  5146.21917865266, 5146.21917865266, 5130.5142314379, 5111.45367395597, 
    5098.66022087426, 5099.38474696456, 5111.07325669628, 5122.69199744876, 
    5116.84029818707, 5071.59309554911, 4992.31657389434, 4922.65026436163, 
    4880.75897154188, 4849.25680825932, 4829.06982285497, 4824.11821546715, 
    4817.9895359485, 4807.30427498796, 4802.63851679231, 4800.47860369378, 
    4786.56429461038, 4756.71252659308, 4725.94913540466, 4705.57636932373, 
    4685.38639863575, 4649.34244850199, 4591.86038780602, 4517.82591387005, 
    4430.41260237482, 4336.33917868715, 4243.39811826083, 4086.08625529088, 
    3712.99188964242, 3082.46617377548, 2363.74045082882, 1700.02083959312, 
    1181.05917326087, 816.179419198417, 566.530139165009, 396.590716460574, 
    279.266599916123, 199.152883508988, 141.004320834194, 99.1288898794317, 
    70.6338321356094, 52.3837883832172, 40.1896894301902, 31.5995748748693, 
    25.0565945490081, 19.8574133551127, 15.7259832375162, 12.7859964397438, 
    11.0518349948811, 10.2800747563701, 10.0549181389887, 10.0549181389887,
  5162.88918317251, 5162.88918317251, 5137.45214422988, 5105.24156387863, 
    5083.20388945779, 5083.30833025408, 5101.94116544786, 5121.80875134795, 
    5120.09511952797, 5076.64032326632, 4997.86645060181, 4922.27382395131, 
    4871.77628850713, 4838.61491421393, 4819.90348010959, 4813.12007411494, 
    4805.75069982894, 4796.8403012922, 4794.03612663521, 4793.12417743015, 
    4781.43080943953, 4754.17220459011, 4723.49046337874, 4700.60039593835, 
    4677.97598602367, 4637.64098156932, 4570.63339318825, 4484.20027901151, 
    4383.61300523262, 4266.82282893864, 4114.89468148605, 3832.23348024767, 
    3294.11742427269, 2552.28931008592, 1849.48421544287, 1290.50808114165, 
    875.981588372673, 590.375783525561, 399.93392619858, 275.312605870548, 
    192.0469031884, 135.790008706509, 95.1757032073565, 66.2786027706133, 
    47.0576688794302, 35.0387804028303, 27.4226014978858, 22.0640038541592, 
    17.9562040835183, 14.7674378660872, 12.3789868551569, 10.8949028043696, 
    10.2223264155853, 10.0310955856371, 10.0029839377891, 10.0029839377891,
  5176.15916541235, 5176.15916541235, 5143.10547454374, 5099.77308200526, 
    5069.28913238004, 5065.84832059337, 5082.19850684781, 5098.68134721257, 
    5097.4598669813, 5065.19578460196, 5002.89617090307, 4930.95147344904, 
    4866.81387930512, 4817.38321972187, 4790.13190073947, 4781.45742887454, 
    4774.65741142494, 4767.27899810242, 4767.12367988064, 4768.96490446636, 
    4759.27665670042, 4733.92776066712, 4706.08030959187, 4687.70558738151, 
    4670.3384629767, 4631.41761354207, 4557.75671859636, 4456.37143674168, 
    4330.48344391035, 4163.63318405878, 3909.41132926724, 3467.10107177856, 
    2794.92068100642, 2026.83916048148, 1396.59999751819, 952.981885836902, 
    640.426000845145, 427.458484169389, 286.950241446432, 194.490278002865, 
    133.095631723312, 92.7924469017267, 64.475721731366, 44.8174204035951, 
    31.917084413833, 23.9754864126556, 19.3027225302532, 16.1003788893387, 
    13.6551729265486, 11.880080649277, 10.7359352604221, 10.1860477045788, 
    10.0224076750767, 10.0005131170989, 10.0001248664912, 10.0001248664912,
  5190.49000271153, 5190.49000271153, 5154.04106075283, 5101.66983316406, 
    5059.89609810296, 5045.48383366365, 5047.98922608201, 5049.38722622769, 
    5043.56773764359, 5025.41741844366, 4988.74703613935, 4934.83347015575, 
    4869.76620993803, 4807.15467022898, 4769.04117307282, 4757.46417456461, 
    4750.35513134789, 4743.95695448364, 4748.79768189956, 4756.51604654305, 
    4749.23608844465, 4722.91705974371, 4692.9392359658, 4673.6785440653, 
    4658.15870992903, 4622.16393645736, 4546.21137357283, 4428.11076013958, 
    4258.81831383792, 4000.66583884069, 3595.59658158535, 2981.33218784106, 
    2238.65068576824, 1543.1353088323, 1036.88391925549, 703.1331436664, 
    471.554918465099, 311.204526462214, 206.176962460931, 137.666248330503, 
    92.9415810233869, 64.2791451281258, 44.657596877656, 31.3521396018396, 
    22.6673925198056, 17.2855829930371, 14.3301018868186, 12.5535014641448, 
    11.3240329459503, 10.540456048312, 10.1447411855493, 10.0181871666948, 
    10, 10.000019806029, 10, 10,
  5199.52300481727, 5199.52300481727, 5163.56116209495, 5104.42198191636, 
    5049.46722240014, 5020.21690163272, 5006.65335648548, 4993.47638321382, 
    4983.42893008031, 4976.68810447706, 4962.96201999946, 4932.19502389073, 
    4879.78324856891, 4817.32271840589, 4774.50265584544, 4759.51480393845, 
    4749.45383624614, 4741.91772240244, 4749.52713660876, 4759.54742330249, 
    4749.60826114169, 4716.50008334076, 4678.02411533748, 4649.55459298059, 
    4625.78018022577, 4586.6159596643, 4510.50943325523, 4375.61146176183, 
    4135.48775609206, 3732.78859107865, 3161.29302314604, 2442.96767456191, 
    1733.64569739517, 1170.40157220408, 784.529739221816, 526.873764273077, 
    348.036801595876, 224.862756509542, 146.501563078794, 97.5599921298659, 
    66.3908246073321, 45.923354479416, 31.9393025583426, 22.698991026034, 
    16.8322121265398, 13.3322223580698, 11.5983456481262, 10.7812121114461, 
    10.3295129060452, 10.0954833024034, 10.0130965956596, 10, 10, 10, 10, 10,
  5172.77885125431, 5172.77885125431, 5146.95971893599, 5094.40749613154, 
    5036.40458001211, 4998.44596839565, 4976.11602561955, 4957.40656247379, 
    4947.28311547567, 4948.42766996238, 4949.89363590525, 4935.12888535496, 
    4894.03057068821, 4837.25897468012, 4794.75005608659, 4776.64399203855, 
    4763.45455115915, 4753.26239410765, 4756.71723175367, 4760.32042929743, 
    4741.7520204705, 4698.43287393831, 4649.11120138805, 4606.46587495899, 
    4562.79351333728, 4506.87073710926, 4422.31677705593, 4252.63889255741, 
    3895.44488278705, 3318.42290261877, 2633.86384511762, 1927.73197336663, 
    1328.05421995354, 890.66084410437, 589.23412466988, 384.645701229384, 
    248.658245023644, 158.66733086782, 102.942452550315, 68.9917714809962, 
    47.5674038312381, 32.9722252501071, 23.1307091696819, 16.8766766793574, 
    13.1580387477077, 11.2182888505073, 10.4255437263116, 10.155987335909, 
    10.0483464689256, 10.0075820262996, 10, 10, 10, 10, 10, 10,
  5111.14634555927, 5111.14634555927, 5106.26684250578, 5076.24515755, 
    5027.88540409757, 4987.39338863837, 4959.8107474887, 4940.52219438317, 
    4935.88819921325, 4947.27902198854, 4959.27361352726, 4949.05825277259, 
    4908.21957176732, 4853.43283294704, 4811.93323156036, 4791.46126498583, 
    4776.68428685794, 4763.34789424196, 4757.06393648163, 4748.41402147964, 
    4719.91122597929, 4668.12686599268, 4609.93657049945, 4554.56446228579, 
    4491.31270741627, 4411.97153202787, 4286.89088754598, 4014.06849099919, 
    3491.77267499983, 2789.38780962284, 2099.26261300059, 1487.40770222521, 
    1012.06684866134, 675.234849259198, 437.281121230085, 277.144768883424, 
    176.620238729104, 112.895663801299, 73.6599108387008, 49.3232344050752, 
    34.0271065418672, 23.7321368206641, 17.1527504144492, 13.2571637164537, 
    11.2016697522007, 10.3392195191824, 10.0756837160021, 10.0176576270894, 
    10.0031038825953, 10, 10, 10, 10, 10, 10, 10,
  5049.67138595013, 5049.67138595013, 5067.60542406193, 5063.89751079851, 
    5027.89791006065, 4983.53545629374, 4946.16700208192, 4923.72299755764, 
    4927.27133349758, 4951.89349447876, 4970.83309546978, 4956.52677131828, 
    4908.95898213139, 4854.58766776207, 4816.06694550385, 4794.74130811645, 
    4777.76876993947, 4760.60980808219, 4746.04567094837, 4727.83896141457, 
    4692.66132560991, 4636.28879526445, 4572.80886105318, 4511.3712003401, 
    4439.94461384366, 4329.14045770584, 4102.02256111553, 3649.22205601242, 
    2977.10289873391, 2255.68701552403, 1639.63288075758, 1137.09911118288, 
    761.641712868952, 498.854936350624, 315.368254462607, 197.198806933474, 
    126.258718727844, 82.0493841141155, 54.1239438784196, 36.1478147737722, 
    24.9594624553114, 17.7929160663186, 13.5674415653257, 11.3434302398691, 
    10.3733786617825, 10.0688613757661, 10.0074899455388, 10.0007299190201, 
    10, 10, 10, 10, 10, 10, 10, 10,
  4999.03556930938, 4999.03556930938, 5032.14086251412, 5048.28484582927, 
    5023.73569218206, 4978.24449098455, 4934.20304861928, 4908.61071313013, 
    4914.21514607438, 4940.79083122903, 4955.49329669772, 4931.13782760769, 
    4877.5424232746, 4828.98293610024, 4799.90633385549, 4780.44608713745, 
    4758.79576844505, 4737.09632226665, 4720.53233062683, 4700.08086456384, 
    4661.60660176137, 4602.69040983417, 4536.59002524094, 4471.45651343746, 
    4385.51001397637, 4210.34160397227, 3836.85759572864, 3216.67430934666, 
    2482.76587414399, 1812.79939294674, 1275.45036422527, 862.196272294677, 
    568.017740600984, 364.966557312296, 227.183842455158, 142.025400143616, 
    91.7879620845661, 60.5475569673054, 40.2515336648567, 26.9127192972148, 
    18.7547685381955, 13.964586045641, 11.5041184744298, 10.4367013737252, 
    10.0824245746129, 10.0075873411873, 10.0000621687022, 10, 10, 10, 10, 10, 
    10, 10, 10, 10,
  4960.7524801354, 4960.7524801354, 4994.57084579647, 5015.13350185835, 
    4997.99025716321, 4961.20480882811, 4925.8566001965, 4904.17746400561, 
    4902.9481481801, 4914.51958764567, 4913.98546717604, 4878.82474845302, 
    4824.26765752253, 4787.30532704934, 4772.03206176317, 4756.36639128958, 
    4729.57470277127, 4703.70081063454, 4688.20473373084, 4668.13877617017, 
    4626.96933598358, 4566.77400091861, 4499.44130537502, 4422.43737009986, 
    4290.39912446114, 4005.9601969358, 3486.12931013106, 2770.44371614665, 
    2051.15653682688, 1455.25519795456, 988.931305351921, 647.01502956072, 
    418.469072263054, 265.673439604375, 165.100743160168, 103.717307122545, 
    67.1538768619968, 44.4043874423909, 29.6576088912538, 20.1279260834423, 
    14.550396109898, 11.6859547903259, 10.4875128482173, 10.0957659248058, 
    10.0091708644146, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  4936.11912035897, 4936.11912035897, 4955.26915695677, 4960.5002022062, 
    4940.47641760816, 4916.1464097819, 4899.13078528273, 4885.16938159534, 
    4872.31578361781, 4865.37498957917, 4856.38731906834, 4822.71797097881, 
    4774.88373098531, 4748.59270822205, 4742.77001795915, 4730.41738926457, 
    4702.28637805698, 4674.10539449487, 4656.23361632123, 4632.98593479284, 
    4590.44720348649, 4533.11814210648, 4464.8656257746, 4362.05977661571, 
    4145.05030563499, 3710.00894683796, 3062.62802228546, 2318.68245452405, 
    1652.64714112384, 1139.06739681325, 754.005083347575, 480.980258901242, 
    305.566020361594, 191.768871485782, 118.573747201614, 74.5667938930242, 
    48.6774959836614, 32.4361987813435, 21.9168141024988, 15.4326363392078, 
    12.0063423297871, 10.5616434608605, 10.1079274632098, 10.0105873126637, 
    10.0000186791801, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  4887.2560406231, 4887.2560406231, 4886.85201609211, 4872.30271956829, 
    4845.41117668184, 4824.62265897612, 4813.35993617845, 4794.51654393397, 
    4760.33559603793, 4737.99048339646, 4741.34995380856, 4733.1603489658, 
    4702.60013007058, 4682.99510572864, 4679.02690860183, 4668.76873511235, 
    4644.41727821069, 4616.97270816365, 4594.8122023315, 4570.48653589544, 
    4535.84551212804, 4488.70785586877, 4416.70936019091, 4267.84999953574, 
    3928.05440160251, 3326.93224784872, 2602.3534324532, 1903.86770962884, 
    1318.65799925866, 878.724020912957, 567.370566240149, 356.420286038599, 
    224.384368864872, 140.388440220965, 86.6043816278155, 54.4864586683328, 
    36.0163989181802, 24.3523960305856, 16.9100698003414, 12.6953358416383, 
    10.7854145450795, 10.1538714924126, 10.016322574306, 10.0003510627118, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  4801.79829678032, 4801.79829678032, 4785.51058290586, 4760.27810161887, 
    4731.89302069667, 4704.12957670381, 4677.87149238163, 4637.64797039214, 
    4576.49610753292, 4543.10628480412, 4569.3320150847, 4597.44133554402, 
    4588.37273592226, 4570.95688228334, 4560.99418593481, 4547.75532645776, 
    4526.48514915931, 4501.56227442719, 4479.63115942357, 4464.47190245198, 
    4449.58271634254, 4415.25625921267, 4323.48379599903, 4093.9535581332, 
    3613.50625994771, 2891.45755600271, 2159.08970711296, 1544.57184634539, 
    1049.44547308013, 677.205531527741, 427.456807627975, 266.603101496854, 
    166.82201155934, 103.777496806263, 63.8559358322598, 40.4197198224133, 
    27.2239126381836, 18.9252187079723, 13.8459601936894, 11.2712268461851, 
    10.2901542475205, 10.0386291354675, 10.0019966973595, 10, 10, 10, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 10,
  4727.02285991146, 4727.02285991146, 4700.09419700867, 4669.80933413962, 
    4644.47163112952, 4613.04518300323, 4573.79041006497, 4521.68505216492, 
    4456.60375689636, 4426.78738177263, 4462.52369024686, 4505.23214129452, 
    4507.25153800635, 4486.0186349032, 4460.61721341729, 4433.37625374002, 
    4406.76041372769, 4382.44744662599, 4364.97764915308, 4362.49232863653, 
    4363.75760168316, 4326.65549809419, 4181.76299396045, 3837.92591288345, 
    3236.56927857968, 2478.44917265539, 1788.36256914993, 1244.14215094085, 
    824.585568336075, 518.778090443587, 322.10498843693, 199.737512531272, 
    124.077253582492, 76.9107029059059, 47.7679686550082, 30.8773733078067, 
    21.3615529599495, 15.4812555338298, 12.0779116061839, 10.5547135738679, 
    10.089561163426, 10.0063246827668, 10, 10, 10, 10, 10, 10, 10, 10, 10, 
    10, 10, 10, 10, 10,
  4616.05449450345, 4616.05449450345, 4601.03653710479, 4586.22050354798, 
    4574.76344804034, 4552.14367188861, 4519.22691564942, 4482.91941923461, 
    4447.09309708272, 4437.32644167042, 4468.88797284249, 4506.15544018085, 
    4513.58556342406, 4490.63935297604, 4451.72445858854, 4410.87017159726, 
    4376.48254456304, 4350.4134254351, 4335.19351656813, 4334.74092718997, 
    4330.1295967234, 4259.6738474441, 4023.73375463756, 3540.83502032133, 
    2835.44619178622, 2091.26124286338, 1471.35991090596, 993.821038231705, 
    642.080148015422, 399.589818434971, 246.931965177376, 152.587296351689, 
    94.4736174182958, 58.9581120114086, 37.3573099043511, 24.6803019014494, 
    17.4346756049812, 13.2064277319777, 11.0139187523135, 10.2001808377869, 
    10.0194124334715, 10.0004873000753, 10.0000163860455, 10, 10, 10, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 10,
  4388.45499413225, 4388.45499413225, 4412.69757254262, 4440.76188122343, 
    4454.32642340893, 4443.77695655915, 4424.46768529927, 4413.32664300872, 
    4409.57122898848, 4418.14821171211, 4447.08789598383, 4482.15217749897, 
    4495.30518449382, 4473.64010733752, 4437.19847774213, 4407.34070341218, 
    4380.62483518681, 4353.02347285656, 4330.59419387152, 4315.90856727412, 
    4285.70621593811, 4160.74555217737, 3814.28253741995, 3200.28907781825, 
    2431.78566404984, 1734.79638011504, 1200.67737018551, 799.319378354336, 
    509.612915096757, 315.219875520945, 193.706380174743, 119.702740590367, 
    74.2576921658226, 46.669016521812, 30.1132972141873, 20.2981912957317, 
    14.6621559315857, 11.6881776614399, 10.4203373138598, 10.0609453682501, 
    10.0045036418369, 10.0002203215302, 10, 10, 10, 10, 10, 10, 10, 10, 10, 
    10, 10, 10, 10, 10,
  4149.01571339975, 4149.01571339975, 4191.11783336121, 4234.2288353717, 
    4250.47238350395, 4237.75698057301, 4218.22134864859, 4208.4366488055, 
    4204.09362988181, 4205.28522337295, 4219.46656473449, 4237.1296682332, 
    4229.27669817631, 4189.14028064601, 4161.62444589177, 4169.09854893174, 
    4170.94919985913, 4141.98212772406, 4098.96990739928, 4060.95489038577, 
    4010.76472146909, 3852.84221657056, 3442.31324699904, 2784.20820042765, 
    2049.46686233756, 1435.57960024816, 981.344750877847, 647.782117235577, 
    409.57694668889, 251.592217689998, 154.366489527467, 96.4991507057383, 
    60.3806643385852, 37.9789708407552, 24.7196635371172, 17.0299890653755, 
    12.7863374491214, 10.826809723809, 10.162936549461, 10.0191001679898, 
    10.0011720352377, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  4011.82008535928, 4011.82008535928, 4022.77013449021, 4024.52799336808, 
    4010.78749904848, 3985.41248286322, 3953.91220086486, 3919.22495296686, 
    3881.89234099429, 3844.30611396935, 3810.79752490424, 3777.46961865125, 
    3724.85186977377, 3658.5723129732, 3638.39722250391, 3680.9218484277, 
    3712.13401644999, 3678.15102469608, 3601.67619379714, 3537.70342723393, 
    3494.63771680641, 3369.43022728182, 2998.76586075633, 2402.19150986505, 
    1760.48797606723, 1222.70201868364, 823.400597087819, 537.986253902339, 
    337.879047583519, 206.748290785476, 127.237959422347, 80.7134230333706, 
    51.1939192039835, 32.3088767537537, 21.1801595174696, 14.8887054020675, 
    11.6544994903164, 10.3885464101792, 10.0561648541273, 10.0039138060888, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3923.12609855637, 3923.12609855637, 3897.27893508507, 3857.74517083855, 
    3822.88815990133, 3796.59583501158, 3760.55006921451, 3702.87291545834, 
    3631.02544026278, 3546.51799708542, 3452.41398045105, 3368.12896878141, 
    3299.58195181178, 3247.90923595321, 3243.95261704729, 3292.21983622061, 
    3326.61324852029, 3279.24864302443, 3163.02321652507, 3070.35644726451, 
    3046.01107933634, 2983.92055337905, 2694.8276608548, 2175.56065571925, 
    1608.58668972091, 1114.74849759263, 742.356287198545, 480.891512511174, 
    302.19965160457, 185.384163831752, 113.77572585922, 72.3094678372059, 
    46.42866874255, 29.5464977727653, 19.4295727901744, 13.7534319267703, 
    11.0665614626471, 10.190052993248, 10.0181144689625, 10.000671067418, 
    10.0000219641831, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3830.14602593956, 3830.14602593956, 3796.77393253335, 3753.43012995293, 
    3722.95904793933, 3704.97085505299, 3667.14149475081, 3593.38049263348, 
    3502.37885758472, 3397.16478963598, 3278.20865563353, 3180.62448664423, 
    3131.50456221156, 3122.42693791535, 3139.40436342407, 3171.80441522109, 
    3185.25358566856, 3118.93934036762, 2971.38382772115, 2850.60827525239, 
    2827.24903922201, 2803.84146300579, 2573.32233960731, 2094.26522599658, 
    1558.12500290486, 1083.06340921438, 718.22429956445, 459.655875840931, 
    287.326002896674, 176.654020009561, 108.330064043346, 68.4542851635969, 
    44.1676615910654, 28.5025092075394, 18.8260300336639, 13.294449866969, 
    10.8350610039873, 10.1280246815522, 10.010377638874, 10.0003480749477, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3756.17000237666, 3756.17000237666, 3731.59775036371, 3697.89985381481, 
    3673.44729274386, 3659.06736079483, 3616.522612787, 3530.44847371164, 
    3436.42169729927, 3347.12230889334, 3253.16641624978, 3175.35734826599, 
    3142.18137237787, 3151.82462844282, 3176.83620189116, 3194.83473797697, 
    3185.66539703096, 3105.60199465358, 2951.16214430058, 2815.29884462757, 
    2765.79002043676, 2721.5564003064, 2484.97052859275, 2005.30229549282, 
    1483.8020090508, 1034.9483369041, 685.534354371935, 432.531750335323, 
    267.720081221938, 164.848639243923, 101.399602204598, 63.7789489994822, 
    41.1964088088524, 27.1192355027574, 18.2721508752003, 13.0352800675696, 
    10.7484588459055, 10.1163292253955, 10.0108887368136, 10.0005269121419, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3720.24622881651, 3720.24622881651, 3695.54889929353, 3655.3178991069, 
    3624.11154851884, 3615.2774174082, 3587.00269735964, 3514.62787944754, 
    3436.57113291195, 3372.37081772538, 3307.85480079123, 3247.79033189277, 
    3213.85813625765, 3214.52395771136, 3232.01116241345, 3240.22188594625, 
    3216.59664886538, 3134.97923687234, 2997.61521045526, 2862.94380882712, 
    2774.33067701416, 2667.35003963622, 2378.71191870917, 1884.97711330584, 
    1376.95492747365, 954.356378739467, 627.758077957933, 392.102709787848, 
    241.472409867714, 148.547981560455, 91.3425243066205, 57.5082062153008, 
    37.285122085822, 24.9647786970087, 17.2894918025721, 12.6383929758253, 
    10.6177444727306, 10.0842063575763, 10.0052652755136, 10, 10, 10, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3716.99767974781, 3716.99767974781, 3678.25832845059, 3619.3481973661, 
    3578.98294620222, 3580.66382591329, 3582.46677093211, 3546.74692074078, 
    3494.89193962983, 3442.79013746363, 3383.50459174402, 3324.26536892205, 
    3283.71319416693, 3270.7649196346, 3274.62306323157, 3272.03484565554, 
    3239.09967630765, 3159.91708456433, 3040.53870222754, 2914.42136531486, 
    2799.83284512515, 2629.85572292145, 2272.60277944449, 1759.53226880811, 
    1264.68362608744, 864.450358355574, 564.588416286183, 352.71030742076, 
    217.840121577415, 134.238343526031, 82.6648845486766, 52.2208072088846, 
    33.8973636624134, 22.8031994445339, 16.1051298486417, 12.1401899689354, 
    10.4797250943687, 10.0645052237544, 10.0052237701732, 10.0002766630273, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3736.28565796575, 3736.28565796575, 3683.85251007521, 3615.95814850175, 
    3576.4561970644, 3581.73833716013, 3595.63839706645, 3582.16942632036, 
    3546.37228134537, 3497.84373656117, 3438.04372236093, 3377.12961270603, 
    3330.73820049205, 3307.07070025587, 3299.09884507364, 3287.33571702546, 
    3247.77171976569, 3164.9535493562, 3046.99423822845, 2923.57069301325, 
    2798.1523242531, 2586.94181610343, 2178.71239155108, 1662.17362922171, 
    1187.79618214915, 803.992203700001, 522.539859712086, 327.775364220996, 
    202.705972496952, 124.106734267115, 76.1232537808751, 48.4713930723974, 
    31.8959471079217, 21.6209966503862, 15.3594947519482, 11.7901869316948, 
    10.3819289178249, 10.0480937502139, 10.0029210821302, 10, 10, 10, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3766.43139210862, 3766.43139210862, 3711.06324913093, 3647.06758155152, 
    3612.36560926698, 3610.32555351616, 3613.48694024747, 3597.28754875667, 
    3561.59773327584, 3514.83617485023, 3461.32958366229, 3403.86920943719, 
    3352.35273834959, 3319.09448395071, 3302.33672306021, 3284.63474608588, 
    3242.33810390076, 3159.85853279641, 3046.21335938782, 2931.27604315517, 
    2809.19845032487, 2576.97316288632, 2132.5644272541, 1613.04675549634, 
    1153.82176914793, 779.560088771833, 504.299154919435, 316.075452833303, 
    195.567909773856, 119.593407756097, 73.3284296905944, 46.8801858944773, 
    31.0865143622674, 21.0405844248915, 14.814413826028, 11.4585970066919, 
    10.2696036699213, 10.0277665914582, 10.0015117598835, 10.0000644610775, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3785.97291950549, 3785.97291950549, 3735.47128349476, 3677.72400805657, 
    3643.28818126647, 3631.10779813846, 3620.56070608258, 3593.7420938922, 
    3550.20151471266, 3501.57446042461, 3454.21813534855, 3403.29615594604, 
    3351.71756966819, 3312.05053561855, 3285.11726821828, 3256.89411721658, 
    3210.83734364855, 3138.32030975494, 3047.37269968776, 2957.42172230504, 
    2848.48203807726, 2605.29489710413, 2134.95632716296, 1607.2927402674, 
    1152.63687469323, 779.831588123358, 499.787673613171, 310.108315876548, 
    191.719631113694, 118.150306165818, 72.7527866488589, 46.319504692059, 
    30.6444410651756, 20.6318629126344, 14.486368689276, 11.3010873725727, 
    10.2267215032046, 10.0210294100446, 10.0008019045596, 10, 10, 10, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3779.09992050158, 3779.09992050158, 3733.31021054086, 3679.86662343366, 
    3644.63435538579, 3626.01537761518, 3608.18520875199, 3575.0867819061, 
    3522.37510243825, 3462.27413769126, 3408.30167413314, 3361.13412303453, 
    3316.9444779573, 3273.87790446115, 3228.74522142682, 3178.93079666831, 
    3125.16525359895, 3066.06640326213, 3004.88653409442, 2950.78708672352, 
    2869.83867834626, 2637.11394303528, 2162.20937799443, 1623.67061799859, 
    1164.25694904175, 790.624043431336, 505.030056301288, 310.513012869916, 
    190.248297208593, 117.49229935716, 72.8915574395726, 46.2716199110048, 
    30.4900634115824, 20.5213283760692, 14.5349065320772, 11.397090433298, 
    10.2733049609116, 10.0311343506842, 10.0016709838558, 10, 10, 10, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3770.37106395758, 3770.37106395758, 3727.66262426148, 3677.79487182195, 
    3641.82973694807, 3616.61817776818, 3593.8714076632, 3559.62947989686, 
    3496.21506893784, 3405.93796086025, 3315.24705610092, 3250.74421773149, 
    3207.06345318788, 3154.64134846657, 3083.4690277705, 3013.87613723076, 
    2969.4752968327, 2944.60187941578, 2924.74619928355, 2910.88413079755, 
    2864.04190116884, 2655.15334139847, 2186.00261124401, 1626.13337927985, 
    1155.21826990411, 788.021990387383, 508.847757219354, 315.307610754392, 
    191.852692729502, 117.55591976617, 73.1582144671892, 46.3645595194407, 
    30.4747314208694, 20.5937897053354, 14.7030713228801, 11.5157501208775, 
    10.3139902368163, 10.0395225961707, 10.0030038841453, 10.0001466653355, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3787.00453013841, 3787.00453013841, 3748.18155478593, 3701.74353082747, 
    3662.60429189536, 3627.60236257049, 3598.03407212345, 3559.8422170101, 
    3475.08027485218, 3331.75251145273, 3174.85727707907, 3069.22497822846, 
    3014.70174070946, 2953.66596259823, 2869.81141533781, 2804.87034301405, 
    2797.29527579928, 2828.80917568083, 2859.89167364941, 2880.73457821072, 
    2860.08164813801, 2677.31779950809, 2214.53284012439, 1620.66902439342, 
    1126.22091088626, 764.405815633645, 498.435624770413, 313.877451018635, 
    192.040428231099, 116.943125070791, 72.4457974204533, 45.8601525100039, 
    30.2627637243165, 20.6150265827902, 14.7619088353863, 11.534693347568, 
    10.3132324214944, 10.0375027418047, 10.0022000483977, 10, 10, 10, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3810.90452121907, 3810.90452121907, 3774.04564659813, 3728.77663965445, 
    3687.14784112389, 3646.33529705733, 3608.20328049974, 3551.12354545534, 
    3424.74582532088, 3219.52203722426, 3003.67622809467, 2867.81591998379, 
    2816.06137915023, 2776.80662871119, 2723.7470652982, 2693.3691659231, 
    2718.04750395417, 2777.98846288656, 2832.95102779353, 2868.50567497877, 
    2857.79125886445, 2691.70776270657, 2244.98255873436, 1647.72272806123, 
    1144.11751237036, 776.883691224685, 506.803288714702, 319.834764285614, 
    196.799145528879, 120.39241749602, 74.7232356686049, 47.2925849000243, 
    31.1673149998432, 21.2292384939373, 15.0484224300297, 11.6057301119406, 
    10.3130137126761, 10.033150608172, 10.0017039022688, 10.0000784029565, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3826.24917714508, 3826.24917714508, 3785.20530745337, 3734.48102224701, 
    3690.21602185763, 3648.20898339941, 3596.96854340373, 3503.36913372661, 
    3325.41562825746, 3078.19039210233, 2844.60241076616, 2708.46733948161, 
    2675.11539980514, 2684.3773088691, 2696.39135222079, 2712.79359651867, 
    2745.47165199874, 2789.85047035293, 2832.26740029155, 2862.61839969347, 
    2848.78836997392, 2687.39212418284, 2262.7314139474, 1695.0171320809, 
    1202.51645685028, 823.584910375753, 538.120248992009, 341.23550597022, 
    212.448270831842, 130.67927067047, 81.0151634184398, 51.0240930345213, 
    33.4061189932241, 22.722988316686, 15.9439132355225, 12.0313295356759, 
    10.4500524224869, 10.0588453255851, 10.0036634033917, 10, 10, 10, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3836.67970979765, 3836.67970979765, 3788.82657344893, 3726.89409667394, 
    3671.66182768311, 3618.13599571289, 3542.76337736069, 3409.14858692464, 
    3196.47440012559, 2945.08151768468, 2730.53022747171, 2603.16004228534, 
    2575.30557134341, 2624.1802720423, 2697.54571719374, 2752.69194474371, 
    2785.69800274958, 2811.73165315974, 2840.31268238535, 2863.42456006567, 
    2844.82887796461, 2686.41494420883, 2279.6090590975, 1736.08155520326, 
    1253.10555290749, 866.173066508666, 569.752058839368, 364.088643152935, 
    229.115634933454, 141.390835052224, 87.6105056749991, 55.0660960151001, 
    35.9739055743272, 24.5105924984576, 17.1136321767876, 12.645879402195, 
    10.6633023964596, 10.1042280834232, 10.0097735490412, 10.000499057799, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3830.06558168122, 3830.06558168122, 3783.0639687308, 3713.90435324358, 
    3636.77288851886, 3550.36493408301, 3440.58824222145, 3281.70588278163, 
    3063.28772790563, 2829.55400187284, 2637.11158882882, 2507.46407039906, 
    2470.37265893751, 2544.92525306347, 2665.56066518311, 2750.32071640152, 
    2789.55245219945, 2814.00585764589, 2840.90777973695, 2858.00485841671, 
    2829.3642668483, 2667.57576174616, 2270.55191960345, 1739.65932049677, 
    1263.34925892018, 881.678577116521, 586.007485622678, 375.083865648626, 
    236.320602510571, 146.191076122639, 90.9251041023366, 57.3284031190375, 
    37.3524302418679, 25.3441585345462, 17.7189592063586, 13.0430857551887, 
    10.8180111709486, 10.134317589676, 10.0116261986514, 10.0003634929987, 
    10.0000077554596, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3802.15204034138, 3802.15204034138, 3765.37841647344, 3695.28613457666, 
    3591.98235145781, 3465.6869152746, 3325.52728755556, 3158.99436835873, 
    2950.15257112809, 2728.00079121552, 2538.10336899804, 2403.79224667504, 
    2369.80785373108, 2466.29852420229, 2616.84642755758, 2723.12301422135, 
    2772.9972479066, 2801.39109430931, 2826.50783475358, 2836.21006000407, 
    2799.3461496401, 2635.38896832646, 2242.69427422312, 1712.73200389932, 
    1234.05471749743, 863.135349584512, 580.14021345108, 372.145411064465, 
    234.088969871937, 145.360034676313, 91.1085020748485, 57.8197958120538, 
    37.5484813533953, 25.2773242726104, 17.6758885870166, 13.068173079907, 
    10.8459652836869, 10.146477390609, 10.0148185461538, 10.000754886756, 10, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3778.79804664165, 3778.79804664165, 3749.51731090375, 3673.54179673781, 
    3547.95752239168, 3401.30301800498, 3250.04604783059, 3080.35133726789, 
    2874.73340300715, 2652.60001972522, 2461.80935754064, 2346.00433934281, 
    2340.74775561861, 2444.8267981641, 2588.28823886034, 2696.59827242508, 
    2754.96417188183, 2784.71065685748, 2801.44717945349, 2799.86693885243, 
    2755.25156495193, 2591.69398952333, 2210.95913516617, 1694.50290515394, 
    1218.42463872552, 851.521640458071, 574.90267282433, 368.662331793596, 
    231.39046020866, 144.588940642391, 91.3151914610899, 58.0951746126923, 
    37.5617429706909, 25.0859508418192, 17.4454620269941, 12.8870792776797, 
    10.7646489808304, 10.1252404242766, 10.0111946193702, 10.0004077381162, 
    10.00001021067, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3775.75040791738, 3775.75040791738, 3741.07336528078, 3647.74614660853, 
    3505.19457721095, 3358.7677354454, 3211.53441498699, 3035.32872085853, 
    2825.02480738228, 2612.29454028369, 2450.48882910879, 2382.20482743985, 
    2408.07134722317, 2491.28885594068, 2591.2435670627, 2678.71649033686, 
    2736.43831046074, 2764.15425642932, 2771.70247040671, 2761.04008684235, 
    2709.92135043171, 2539.29237224339, 2157.99471976666, 1650.47990524466, 
    1181.65780962268, 821.827098054605, 555.031993283505, 356.811640410843, 
    224.248164734375, 140.816453305406, 89.1263373423167, 56.6274641078605, 
    36.575325548786, 24.3992077521229, 16.9555841202019, 12.5605295559016, 
    10.6256451085232, 10.0939515003336, 10.0082518048884, 10.0004013520705, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3774.30511713892, 3774.30511713892, 3722.02640881132, 3605.41496372113, 
    3451.58898334925, 3312.19679722677, 3172.67559623672, 2994.80101367257, 
    2793.77998452109, 2620.47657089486, 2519.20931071974, 2499.44239741186, 
    2528.98933732804, 2568.85861413317, 2614.02226648085, 2667.6995882277, 
    2713.38178167589, 2737.22233270413, 2740.15343597967, 2721.52909247901, 
    2652.04718110552, 2449.09415721091, 2047.70891556169, 1548.70978045019, 
    1096.34821832724, 748.902504035678, 498.954798698815, 321.117181967121, 
    202.889334595096, 127.623465685258, 80.536246372159, 51.2392610399217, 
    33.4764074806315, 22.7593612192297, 16.1248213438673, 12.1854695927934, 
    10.4943208558286, 10.0639125527817, 10.003890674263, 10, 10, 10, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3742.40937917281, 3742.40937917281, 3667.69075306153, 3528.27410023643, 
    3371.07941690616, 3247.55436341361, 3125.9853104461, 2967.26750473498, 
    2807.34210342743, 2695.15554399751, 2644.18742684887, 2638.16198709892, 
    2643.98038120119, 2639.72551657288, 2638.55931407973, 2657.15506296265, 
    2686.67163136688, 2708.45186909086, 2710.59432879473, 2682.28908123772, 
    2581.24081035262, 2321.76704424462, 1883.59757088458, 1394.30263904459, 
    974.27632570438, 653.548843780523, 427.569942456387, 274.236644860368, 
    174.074694317573, 109.879597521087, 69.3922829327741, 44.5589996490174, 
    29.5673381041828, 20.5462905163687, 14.9761426442559, 11.8200462381412, 
    10.4197005037409, 10.0514105035682, 10.0030731138246, 10.0001515995651, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3678.16706666471, 3678.16706666471, 3583.1160127628, 3419.68120110938, 
    3258.44143191066, 3160.59244636033, 3077.50086962804, 2962.86082775365, 
    2862.54632466184, 2803.70451593646, 2765.93473287466, 2738.68239844681, 
    2713.2354872079, 2677.48856314253, 2644.37821930449, 2636.89874970066, 
    2656.5345246997, 2681.2150274215, 2685.42970320551, 2647.17720795862, 
    2509.10193124951, 2186.15419201617, 1712.04226026979, 1234.8336194334, 
    854.655321566952, 567.513976303326, 364.695214906096, 231.157001123888, 
    146.532970017859, 93.006650417408, 59.1388770168702, 38.6344737926224, 
    25.9440851325094, 18.3545612424267, 13.9577118579068, 11.8229992606818, 
    10.5904440576501, 10.1023153257052, 10.0072103617416, 10, 10, 10, 10, 10, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3622.09305312564, 3622.09305312564, 3513.76371953439, 3328.96359973774, 
    3158.13340086309, 3080.8872902217, 3037.9168517577, 2966.38732203885, 
    2908.49674186499, 2875.07392406226, 2830.70040541757, 2780.20857818542, 
    2733.93431995471, 2680.96660286269, 2631.30069423572, 2612.02933430543, 
    2630.16699876587, 2660.16377423538, 2668.13889771827, 2625.35782064925, 
    2464.39136222717, 2102.99587955717, 1609.87547148693, 1137.52055598363, 
    779.499670452809, 512.842704047382, 323.574143185544, 201.987686189467, 
    127.708746679929, 81.6421785162741, 52.3561318136806, 34.754320370818, 
    23.5644375662486, 17.0099337252208, 13.5588512666172, 12.2295888913736, 
    10.9841414746609, 10.2366097670953, 10.0288442602251, 10.0014422130113, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10,
  3622.09305312564, 3622.09305312564, 3513.76371953439, 3328.96359973774, 
    3158.13340086309, 3080.8872902217, 3037.9168517577, 2966.38732203885, 
    2908.49674186499, 2875.07392406226, 2830.70040541757, 2780.20857818542, 
    2733.93431995471, 2680.96660286269, 2631.30069423572, 2612.02933430543, 
    2630.16699876587, 2660.16377423538, 2668.13889771827, 2625.35782064925, 
    2464.39136222717, 2102.99587955717, 1609.87547148693, 1137.52055598363, 
    779.499670452809, 512.842704047382, 323.574143185544, 201.987686189467, 
    127.708746679929, 81.6421785162741, 52.3561318136806, 34.754320370818, 
    23.5644375662486, 17.0099337252208, 13.5588512666172, 12.2295888913736, 
    10.9841414746609, 10.2366097670953, 10.0288442602251, 10.0014422130113, 
    10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10, 10 ;

 lon_rho =
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667 ;

 lat_rho =
  30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30,
  30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333,
  30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667,
  31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 
    31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 
    31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31,
  31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333,
  31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667,
  32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 
    32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 
    32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32,
  32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333,
  32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667,
  33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 
    33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 
    33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33,
  33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333,
  33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667,
  34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 
    34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 
    34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34,
  34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333,
  34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333,
  35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667,
  36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 
    36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 
    36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36,
  36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333,
  36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667,
  37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 
    37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 
    37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37,
  37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333,
  37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667,
  38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 
    38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 
    38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38,
  38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333,
  38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667,
  39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 
    39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 
    39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39,
  39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333,
  39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667,
  40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 
    40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 
    40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40,
  40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333,
  40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667,
  41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 
    41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 
    41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41,
  41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333,
  41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667,
  42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 
    42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 
    42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42,
  42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333,
  42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667,
  43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 
    43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 
    43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43,
  43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333,
  43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667,
  44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 
    44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 
    44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44,
  44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333,
  44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667,
  45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 
    45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 
    45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45,
  45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333,
  45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667,
  46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 
    46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 
    46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46,
  46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333,
  46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667,
  47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 
    47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 
    47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47,
  47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333,
  47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667,
  48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 
    48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 
    48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48 ;

 lon_u =
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333,
  -133.833333333333, -133.5, -133.166666666667, -132.833333333333, -132.5, 
    -132.166666666667, -131.833333333333, -131.5, -131.166666666667, 
    -130.833333333333, -130.5, -130.166666666667, -129.833333333333, -129.5, 
    -129.166666666667, -128.833333333333, -128.5, -128.166666666667, 
    -127.833333333333, -127.5, -127.166666666667, -126.833333333333, -126.5, 
    -126.166666666667, -125.833333333333, -125.5, -125.166666666667, 
    -124.833333333333, -124.5, -124.166666666667, -123.833333333333, -123.5, 
    -123.166666666667, -122.833333333333, -122.5, -122.166666666667, 
    -121.833333333333, -121.5, -121.166666666667, -120.833333333333, -120.5, 
    -120.166666666667, -119.833333333333, -119.5, -119.166666666667, 
    -118.833333333333, -118.5, -118.166666666667, -117.833333333333, -117.5, 
    -117.166666666667, -116.833333333333, -116.5, -116.166666666667, 
    -115.833333333333 ;

 lat_u =
  30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 
    30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30, 30,
  30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333, 30.3333333333333, 
    30.3333333333333, 30.3333333333333, 30.3333333333333,
  30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667, 30.6666666666667, 
    30.6666666666667, 30.6666666666667, 30.6666666666667,
  31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 
    31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 
    31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31, 31,
  31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333, 31.3333333333333, 
    31.3333333333333, 31.3333333333333, 31.3333333333333,
  31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667, 31.6666666666667, 
    31.6666666666667, 31.6666666666667, 31.6666666666667,
  32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 
    32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 
    32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32, 32,
  32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333, 32.3333333333333, 
    32.3333333333333, 32.3333333333333, 32.3333333333333,
  32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667, 32.6666666666667, 
    32.6666666666667, 32.6666666666667, 32.6666666666667,
  33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 
    33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 
    33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33, 33,
  33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333, 33.3333333333333, 
    33.3333333333333, 33.3333333333333, 33.3333333333333,
  33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667, 33.6666666666667, 
    33.6666666666667, 33.6666666666667, 33.6666666666667,
  34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 
    34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 
    34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34, 34,
  34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333, 34.3333333333333, 
    34.3333333333333, 34.3333333333333, 34.3333333333333,
  34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667, 34.6666666666667, 
    34.6666666666667, 34.6666666666667, 34.6666666666667,
  35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 
    35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35, 35,
  35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333, 35.3333333333333, 
    35.3333333333333, 35.3333333333333, 35.3333333333333,
  35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667, 35.6666666666667, 
    35.6666666666667, 35.6666666666667, 35.6666666666667,
  36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 
    36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 
    36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36, 36,
  36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333, 36.3333333333333, 
    36.3333333333333, 36.3333333333333, 36.3333333333333,
  36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667, 36.6666666666667, 
    36.6666666666667, 36.6666666666667, 36.6666666666667,
  37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 
    37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 
    37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37, 37,
  37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333, 37.3333333333333, 
    37.3333333333333, 37.3333333333333, 37.3333333333333,
  37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667, 37.6666666666667, 
    37.6666666666667, 37.6666666666667, 37.6666666666667,
  38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 
    38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 
    38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38, 38,
  38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333, 38.3333333333333, 
    38.3333333333333, 38.3333333333333, 38.3333333333333,
  38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667, 38.6666666666667, 
    38.6666666666667, 38.6666666666667, 38.6666666666667,
  39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 
    39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 
    39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39, 39,
  39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333, 39.3333333333333, 
    39.3333333333333, 39.3333333333333, 39.3333333333333,
  39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667, 39.6666666666667, 
    39.6666666666667, 39.6666666666667, 39.6666666666667,
  40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 
    40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 
    40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40, 40,
  40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333, 40.3333333333333, 
    40.3333333333333, 40.3333333333333, 40.3333333333333,
  40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667, 40.6666666666667, 
    40.6666666666667, 40.6666666666667, 40.6666666666667,
  41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 
    41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 
    41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41, 41,
  41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333, 41.3333333333333, 
    41.3333333333333, 41.3333333333333, 41.3333333333333,
  41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667, 41.6666666666667, 
    41.6666666666667, 41.6666666666667, 41.6666666666667,
  42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 
    42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 
    42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42, 42,
  42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333, 42.3333333333333, 
    42.3333333333333, 42.3333333333333, 42.3333333333333,
  42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667, 42.6666666666667, 
    42.6666666666667, 42.6666666666667, 42.6666666666667,
  43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 
    43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 
    43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43, 43,
  43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333, 43.3333333333333, 
    43.3333333333333, 43.3333333333333, 43.3333333333333,
  43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667, 43.6666666666667, 
    43.6666666666667, 43.6666666666667, 43.6666666666667,
  44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 
    44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 
    44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44, 44,
  44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333, 44.3333333333333, 
    44.3333333333333, 44.3333333333333, 44.3333333333333,
  44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667, 44.6666666666667, 
    44.6666666666667, 44.6666666666667, 44.6666666666667,
  45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 
    45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 
    45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45, 45,
  45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333, 45.3333333333333, 
    45.3333333333333, 45.3333333333333, 45.3333333333333,
  45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667, 45.6666666666667, 
    45.6666666666667, 45.6666666666667, 45.6666666666667,
  46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 
    46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 
    46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46, 46,
  46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333, 46.3333333333333, 
    46.3333333333333, 46.3333333333333, 46.3333333333333,
  46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667, 46.6666666666667, 
    46.6666666666667, 46.6666666666667, 46.6666666666667,
  47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 
    47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 
    47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47, 47,
  47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333, 47.3333333333333, 
    47.3333333333333, 47.3333333333333, 47.3333333333333,
  47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667, 47.6666666666667, 
    47.6666666666667, 47.6666666666667, 47.6666666666667,
  48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 
    48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 
    48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48, 48 ;

 lon_v =
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667,
  -134, -133.666666666667, -133.333333333333, -133, -132.666666666667, 
    -132.333333333333, -132, -131.666666666667, -131.333333333333, -131, 
    -130.666666666667, -130.333333333333, -130, -129.666666666667, 
    -129.333333333333, -129, -128.666666666667, -128.333333333333, -128, 
    -127.666666666667, -127.333333333333, -127, -126.666666666667, 
    -126.333333333333, -126, -125.666666666667, -125.333333333333, -125, 
    -124.666666666667, -124.333333333333, -124, -123.666666666667, 
    -123.333333333333, -123, -122.666666666667, -122.333333333333, -122, 
    -121.666666666667, -121.333333333333, -121, -120.666666666667, 
    -120.333333333333, -120, -119.666666666667, -119.333333333333, -119, 
    -118.666666666667, -118.333333333333, -118, -117.666666666667, 
    -117.333333333333, -117, -116.666666666667, -116.333333333333, -116, 
    -115.666666666667 ;

 lat_v =
  30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667, 
    30.1666666666667, 30.1666666666667, 30.1666666666667, 30.1666666666667,
  30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 
    30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 
    30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 
    30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 
    30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5, 30.5,
  30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333, 
    30.8333333333333, 30.8333333333333, 30.8333333333333, 30.8333333333333,
  31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667, 
    31.1666666666667, 31.1666666666667, 31.1666666666667, 31.1666666666667,
  31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 
    31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 
    31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 
    31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 
    31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5, 31.5,
  31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333, 
    31.8333333333333, 31.8333333333333, 31.8333333333333, 31.8333333333333,
  32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667, 
    32.1666666666667, 32.1666666666667, 32.1666666666667, 32.1666666666667,
  32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 
    32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 
    32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 
    32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 
    32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5, 32.5,
  32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333, 
    32.8333333333333, 32.8333333333333, 32.8333333333333, 32.8333333333333,
  33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667, 
    33.1666666666667, 33.1666666666667, 33.1666666666667, 33.1666666666667,
  33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 
    33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 
    33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 
    33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 
    33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5, 33.5,
  33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333, 
    33.8333333333333, 33.8333333333333, 33.8333333333333, 33.8333333333333,
  34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667, 
    34.1666666666667, 34.1666666666667, 34.1666666666667, 34.1666666666667,
  34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 
    34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 
    34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 
    34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 
    34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5, 34.5,
  34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333, 
    34.8333333333333, 34.8333333333333, 34.8333333333333, 34.8333333333333,
  35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667, 
    35.1666666666667, 35.1666666666667, 35.1666666666667, 35.1666666666667,
  35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 
    35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 
    35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 
    35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 
    35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5, 35.5,
  35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333, 
    35.8333333333333, 35.8333333333333, 35.8333333333333, 35.8333333333333,
  36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667, 
    36.1666666666667, 36.1666666666667, 36.1666666666667, 36.1666666666667,
  36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 
    36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 
    36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 
    36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 
    36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5, 36.5,
  36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333, 
    36.8333333333333, 36.8333333333333, 36.8333333333333, 36.8333333333333,
  37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667, 
    37.1666666666667, 37.1666666666667, 37.1666666666667, 37.1666666666667,
  37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 
    37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 
    37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 
    37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 
    37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5, 37.5,
  37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333, 
    37.8333333333333, 37.8333333333333, 37.8333333333333, 37.8333333333333,
  38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667, 
    38.1666666666667, 38.1666666666667, 38.1666666666667, 38.1666666666667,
  38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 
    38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 
    38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 
    38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 
    38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5, 38.5,
  38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333, 
    38.8333333333333, 38.8333333333333, 38.8333333333333, 38.8333333333333,
  39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667, 
    39.1666666666667, 39.1666666666667, 39.1666666666667, 39.1666666666667,
  39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 
    39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 
    39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 
    39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 
    39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5, 39.5,
  39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333, 
    39.8333333333333, 39.8333333333333, 39.8333333333333, 39.8333333333333,
  40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667, 
    40.1666666666667, 40.1666666666667, 40.1666666666667, 40.1666666666667,
  40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 
    40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 
    40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 
    40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 
    40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5, 40.5,
  40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333, 
    40.8333333333333, 40.8333333333333, 40.8333333333333, 40.8333333333333,
  41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667, 
    41.1666666666667, 41.1666666666667, 41.1666666666667, 41.1666666666667,
  41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 
    41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 
    41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 
    41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 
    41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5, 41.5,
  41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333, 
    41.8333333333333, 41.8333333333333, 41.8333333333333, 41.8333333333333,
  42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667, 
    42.1666666666667, 42.1666666666667, 42.1666666666667, 42.1666666666667,
  42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 
    42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 
    42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 
    42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 
    42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5, 42.5,
  42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333, 
    42.8333333333333, 42.8333333333333, 42.8333333333333, 42.8333333333333,
  43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667, 
    43.1666666666667, 43.1666666666667, 43.1666666666667, 43.1666666666667,
  43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 
    43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 
    43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 
    43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 
    43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5, 43.5,
  43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333, 
    43.8333333333333, 43.8333333333333, 43.8333333333333, 43.8333333333333,
  44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667, 
    44.1666666666667, 44.1666666666667, 44.1666666666667, 44.1666666666667,
  44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 
    44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 
    44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 
    44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 
    44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5, 44.5,
  44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333, 
    44.8333333333333, 44.8333333333333, 44.8333333333333, 44.8333333333333,
  45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667, 
    45.1666666666667, 45.1666666666667, 45.1666666666667, 45.1666666666667,
  45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 
    45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 
    45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 
    45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 
    45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5, 45.5,
  45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333, 
    45.8333333333333, 45.8333333333333, 45.8333333333333, 45.8333333333333,
  46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667, 
    46.1666666666667, 46.1666666666667, 46.1666666666667, 46.1666666666667,
  46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 
    46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 
    46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 
    46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 
    46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5, 46.5,
  46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333, 
    46.8333333333333, 46.8333333333333, 46.8333333333333, 46.8333333333333,
  47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667, 
    47.1666666666667, 47.1666666666667, 47.1666666666667, 47.1666666666667,
  47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 
    47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 
    47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 
    47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 
    47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5, 47.5,
  47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333, 
    47.8333333333333, 47.8333333333333, 47.8333333333333, 47.8333333333333 ;

 zeta_time = 1123204320, 1125839520 ;

 v2d_time = 1123204320, 1125839520 ;

 v3d_time = 1123204320, 1125839520 ;

 temp_time = 1123204320, 1125839520 ;

 salt_time = 1123204320, 1125839520 ;

 zeta_west =
  0.1945676, 0.1911008, 0.1886568, 0.1872354, 0.184538, 0.1813965, 0.1778111, 
    0.1749165, 0.1702828, 0.1639102, 0.1572976, 0.1491248, 0.1393919, 
    0.1309063, 0.1212435, 0.1104036, 0.09756559, 0.08629598, 0.0765948, 
    0.06374691, 0.05341868, 0.04561009, 0.04148169, 0.03774762, 0.03440788, 
    0.03019939, 0.02458951, 0.01757825, 0.01312846, 0.006773788, 
    -0.001485771, -0.006856885, -0.0105803, -0.01265601, -0.01573393, 
    -0.01499586, -0.0104418, -0.006481897, -0.004119, -0.00335311, 
    -0.001812206, -0.005742479, -0.01514393, -0.02444928, -0.03660941, 
    -0.05162434, -0.06495959, -0.07825489, -0.09151025, -0.103099, 
    -0.1146492, -0.1261611, -0.1368219, -0.1473367, -0.1577057,
  0.1951549, 0.192003, 0.1894616, 0.1875308, 0.1852772, 0.1822626, 0.1784867, 
    0.1747626, 0.1694345, 0.1625024, 0.1554828, 0.1471121, 0.1373906, 
    0.1277605, 0.1170785, 0.1053445, 0.09261651, 0.08148928, 0.0719628, 
    0.05915555, 0.04898652, 0.04145573, 0.03755954, 0.03387873, 0.03041329, 
    0.02674029, 0.02202684, 0.01627295, 0.01282705, 0.007923776, 0.001563141, 
    -0.00328981, -0.007894522, -0.012251, -0.01633475, -0.01837307, 
    -0.01836595, -0.01956202, -0.02190558, -0.02539662, -0.0263586, 
    -0.03145717, -0.04069231, -0.04962564, -0.06122154, -0.07548001, 
    -0.0871397, -0.09905261, -0.1112187, -0.1208228, -0.1302656, -0.1395469, 
    -0.148397, -0.1571029, -0.1656648 ;

 zeta_east =
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0 ;

 zeta_south =
  0.1945676, 0.1913858, 0.1885075, 0.1859328, 0.1827619, 0.1802939, 
    0.1785288, 0.1762543, 0.1743248, 0.1727402, 0.1721051, 0.1716063, 
    0.1712438, 0.1700035, 0.1685078, 0.1667569, 0.1645189, 0.1612801, 
    0.1570406, 0.1527299, 0.1476703, 0.1418619, 0.1355231, 0.1292078, 
    0.1229162, 0.116244, 0.1099082, 0.1039089, 0.09854188, 0.0941123, 
    0.09062021, 0.08581141, 0.08191128, 0.0789198, 0.0769787, 0.07482707, 
    0.07246492, 0.06862932, 0.06378215, 0.0579234, 0.05401693, 0.04924937, 
    0.0436207, 0.03663502, 0.02921179, 0.02135102, 0.01405958, 0.005809117, 
    -0.003400377, -0.01275739, -0.02060301, -0.02693722, -0.03802665, 
    -0.03990405, -0.03256943, 0,
  0.1951549, 0.1912799, 0.1876969, 0.1844061, 0.1808648, 0.1781546, 
    0.1762755, 0.173883, 0.1717958, 0.1700139, 0.1694019, 0.1689055, 
    0.1685247, 0.167017, 0.1655804, 0.1642149, 0.1621823, 0.1593458, 
    0.1557053, 0.1517138, 0.1467316, 0.1407588, 0.1344837, 0.1280809, 
    0.1215505, 0.1144281, 0.1080283, 0.102351, 0.09680924, 0.09243736, 
    0.08923532, 0.08489908, 0.08112877, 0.07792439, 0.07620013, 0.07407444, 
    0.07154734, 0.06701269, 0.06151551, 0.0550558, 0.05055283, 0.04495985, 
    0.03827687, 0.03027446, 0.0223276, 0.01443629, 0.006397631, 
    -0.0006230123, -0.00662564, -0.01456061, -0.02048834, -0.02440883, 
    -0.03345758, -0.03535367, -0.03009711, 0 ;

 zeta_north =
  -0.1577057, -0.15413, -0.1503812, -0.1464594, -0.1433677, -0.1403997, 
    -0.1375553, -0.134531, -0.1320268, -0.1300428, -0.1274975, -0.1245822, 
    -0.1212967, -0.1206422, -0.1217769, -0.1247008, -0.1244928, -0.1260299, 
    -0.1293122, -0.1283505, -0.1190652, -0.1014563, -0.09761346, -0.08200509, 
    -0.05463113, -0.04198333, -0.04150527, -0.05319695, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -0.1656648, -0.1627909, -0.1597072, -0.1564135, -0.1531284, -0.1504281, 
    -0.1483127, -0.1458311, -0.1439497, -0.1426683, -0.1412403, -0.1382686, 
    -0.1337532, -0.1323863, -0.1309955, -0.129581, -0.123249, -0.1188593, 
    -0.1164119, -0.1102338, -0.1006279, -0.08759432, -0.08209626, 
    -0.07432818, -0.06429006, -0.05579513, -0.05357947, -0.05764308, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ubar_west =
  -0.0006678975, -0.0006789418, -0.0005143251, -0.0004785315, -0.0004512053, 
    -0.0005631825, -0.0005696236, -0.0005752319, -0.0003281413, 0.000385789, 
    0.00112311, 0.002211783, 0.003617904, 0.004993822, 0.005837638, 
    0.006583156, 0.007330678, 0.007377854, 0.006723282, 0.006079467, 
    0.005490072, 0.004789858, 0.004079824, 0.003782501, 0.003417528, 
    0.003050125, 0.002706425, 0.0023379, 0.001962804, 0.0017354, 0.001536858, 
    0.001327009, 0.001014114, 0.000600455, 0.0001827057, -0.0001674389, 
    -0.0004019918, -0.0006281966, -0.0006753055, -0.0004176237, 
    -0.0001686754, 9.742409e-05, 0.0005219372, 0.0009406779, 0.001313346, 
    0.001724551, 0.002141546, 0.002468072, 0.002691254, 0.002903633, 
    0.003064252, 0.00305954, 0.003076572, 0.002928334, 0.002697593,
  -0.0005773077, -0.0006865971, -0.0007935485, -0.0009777711, -0.001168132, 
    -0.001342944, -0.001363853, -0.001383598, -0.001136337, -0.0005008977, 
    0.0001555522, 0.001058109, 0.002183117, 0.00328482, 0.003963977, 
    0.004583369, 0.005203748, 0.005335466, 0.004977832, 0.004629301, 
    0.004293595, 0.003917004, 0.003535836, 0.003518185, 0.003381468, 
    0.00324757, 0.003058961, 0.002786923, 0.002505706, 0.002332514, 
    0.00226648, 0.002196437, 0.002064368, 0.001909205, 0.001755282, 
    0.001614091, 0.001463287, 0.001314355, 0.001201604, 0.001191301, 
    0.001178929, 0.00115285, 0.001244041, 0.00133141, 0.001426991, 
    0.001621732, 0.001820963, 0.001946644, 0.001988816, 0.002022952, 
    0.002078814, 0.001991602, 0.001918952, 0.001738258, 0.001550777 ;

 ubar_east =
  0.005035975, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.003648904, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 ubar_south =
  -0.0006678975, -0.0006568531, -0.0003181022, -2.85883e-05, 0.0001999014, 
    0.0005586869, 0.0009310374, 0.001350019, 0.001853967, 0.002450457, 
    0.003127038, 0.003358196, 0.003644508, 0.003986313, 0.004086371, 
    0.004164411, 0.004232616, 0.004249408, 0.004195256, 0.004060653, 
    0.003978458, 0.003854235, 0.003692679, 0.003508163, 0.003376184, 
    0.003285046, 0.003098401, 0.002956955, 0.002866965, 0.002858127, 
    0.002874998, 0.002924636, 0.002900392, 0.002881713, 0.002853606, 
    0.002881385, 0.002903544, 0.002932447, 0.002996576, 0.00302816, 
    0.00303291, 0.002970122, 0.002875475, 0.002742677, 0.002629007, 
    0.002599201, 0.002786038, 0.003255715, 0.004127074, 0.004946665, 
    0.005852672, 0.007403719, 0.009793968, 0.01007195, 0.005035975,
  -0.0005773077, -0.0004680182, -0.000258686, -7.717728e-05, 7.27586e-05, 
    0.0003320517, 0.000603229, 0.0009057491, 0.001183249, 0.001508892, 
    0.001875915, 0.002067238, 0.002245549, 0.002408562, 0.002480771, 
    0.002499738, 0.002474272, 0.00247291, 0.0024292, 0.00233542, 0.002263934, 
    0.002179781, 0.002086157, 0.002002521, 0.001964942, 0.001964915, 
    0.001903146, 0.001886241, 0.001919485, 0.002014858, 0.002130859, 
    0.002274836, 0.002388245, 0.002499121, 0.002595554, 0.002657089, 
    0.00265517, 0.002601024, 0.002728608, 0.002750837, 0.002668596, 
    0.002399823, 0.002089445, 0.001720773, 0.001327257, 0.001051181, 
    0.001004981, 0.0009570346, 0.00166285, 0.002639964, 0.00348053, 
    0.004713247, 0.006793123, 0.007297809, 0.003648904 ;

 ubar_north =
  0.002697593, 0.002466853, 0.002428511, 0.002325701, 0.002123974, 
    0.00203703, 0.001901265, 0.00171725, 0.001466567, 0.001156317, 
    0.0007914217, 0.0004056503, 3.552365e-05, -0.0003238022, -0.0008845667, 
    -0.001270135, -0.001469915, -0.00180607, -0.001982081, -0.002044724, 
    -0.002568687, -0.003229219, -0.003973703, -0.005820477, -0.007560776, 
    -0.008428942, -0.0119987, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.001550777, 0.001363297, 0.00136214, 0.001393568, 0.00144256, 0.001457369, 
    0.001448067, 0.001415759, 0.001445137, 0.001365172, 0.001171764, 
    0.0009618172, 0.0007014336, 0.0003851004, -5.072015e-05, -0.0003655516, 
    -0.0005513782, -0.0006643839, -0.0006518112, -0.0005317631, 
    -0.0006611814, -0.0009316272, -0.001390741, -0.002336815, -0.003406594, 
    -0.004384436, -0.005952768, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 vbar_west =
  -0.002459162, -0.002522481, -0.002835823, -0.003255516, -0.003797391, 
    -0.004396621, -0.00476712, -0.004904747, -0.005226149, -0.005296425, 
    -0.005143276, -0.004950647, -0.004690541, -0.004350128, -0.003987409, 
    -0.003456859, -0.002751504, -0.00240326, -0.002114364, -0.001895412, 
    -0.001372296, -0.001084445, -0.00102034, -0.0008522703, -0.0007888064, 
    -0.0008351636, -0.0007076785, -0.0007273715, -0.000886076, -0.0009655363, 
    -0.001107838, -0.001322039, -0.00156809, -0.00174535, -0.001842041, 
    -0.002084627, -0.002290328, -0.002459306, -0.002491765, -0.002510578, 
    -0.002514322, -0.002621479, -0.002590537, -0.002435136, -0.002229578, 
    -0.001947263, -0.001589791, -0.001277189, -0.0009596358, -0.0006404914, 
    -0.0004028559, -0.0001298274, 0.0001901424, 0.0002938875,
  -0.002106344, -0.002155531, -0.002346569, -0.002604415, -0.002941107, 
    -0.003229328, -0.003428823, -0.003536057, -0.003654312, -0.003663589, 
    -0.003580265, -0.003479105, -0.003345131, -0.003166744, -0.003033771, 
    -0.00271199, -0.002197865, -0.001978066, -0.001764969, -0.00156714, 
    -0.001106289, -0.0008500108, -0.0007903349, -0.0006887648, -0.0006952091, 
    -0.0008164975, -0.000797425, -0.0008966147, -0.001102451, -0.001199234, 
    -0.001318527, -0.001469449, -0.00160189, -0.001732545, -0.001850907, 
    -0.001923962, -0.002002945, -0.002090001, -0.002256716, -0.002346153, 
    -0.00235765, -0.002606835, -0.00264249, -0.002477853, -0.002293762, 
    -0.001978543, -0.001531945, -0.001224783, -0.0008818972, -0.0005069438, 
    -0.0003108298, -6.700175e-05, 0.0002313026, 0.0003113857 ;

 vbar_east =
  -0.005849799, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0,
  -0.003928086, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 vbar_south =
  -0.002459162, -0.002395843, -0.002675301, -0.003016448, -0.003366251, 
    -0.003787647, -0.004292216, -0.004813739, -0.005178574, -0.005399574, 
    -0.005619864, -0.005442299, -0.004981169, -0.004519816, -0.004134614, 
    -0.003823246, -0.003513574, -0.003165237, -0.003074588, -0.002981987, 
    -0.002812849, -0.00257026, -0.002328485, -0.002002461, -0.00162721, 
    -0.001248831, -0.0008821379, -0.000468913, -5.605029e-05, 0.0002055604, 
    0.0004252014, 0.0006500555, 0.000687491, 0.0005791098, 0.0004675596, 
    0.0001879225, -0.0002963109, -0.000779553, -0.001198042, -0.001677274, 
    -0.00216987, -0.002503135, -0.00267194, -0.002832052, -0.00284977, 
    -0.002871372, -0.003052966, -0.003506596, -0.004180436, -0.00508651, 
    -0.005776213, -0.006271932, -0.006747437, -0.008893793, -0.0116996, 
    -0.005849799,
  -0.002106344, -0.002057157, -0.002158357, -0.002237846, -0.002325681, 
    -0.002485726, -0.002679693, -0.002880517, -0.003067274, -0.00323595, 
    -0.003404372, -0.003383978, -0.003272907, -0.003162332, -0.003075343, 
    -0.003009686, -0.002947022, -0.002813406, -0.002832531, -0.002846407, 
    -0.002812135, -0.002735443, -0.002659855, -0.002529846, -0.002349148, 
    -0.002169572, -0.002008091, -0.001774797, -0.00154165, -0.001430438, 
    -0.001319112, -0.00120654, -0.001159771, -0.001230003, -0.001307322, 
    -0.001417369, -0.001733423, -0.002048881, -0.002202294, -0.002429564, 
    -0.00266505, -0.002676524, -0.002452962, -0.002209491, -0.001825889, 
    -0.001395585, -0.0009274452, -0.0007143891, -0.0005168433, -0.0003126854, 
    -0.0008457602, -0.00186458, -0.003175716, -0.005463152, -0.007856172, 
    -0.003928086 ;

 vbar_north =
  0.0002938875, 0.0003976326, 0.0004422982, 0.0005089536, 0.0005950109, 
    0.0006351805, 0.0005742777, 0.0005105246, 0.0002798535, 0.0002574496, 
    0.0002383988, 0.000332075, 0.0005313156, 0.0007357737, 0.00106312, 
    0.001224649, 0.001367589, 0.001619225, 0.002062282, 0.002553142, 
    0.003197307, 0.00427515, 0.00624533, 0.009317742, 0.01278567, 0.01715379, 
    0.02325564, 0.02834382, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0.0003113857, 0.0003914688, 0.0004731608, 0.0005486783, 0.0006372035, 
    0.0006257062, 0.0004300133, 0.0002280157, 1.114577e-05, 7.828446e-05, 
    0.0001513083, 0.0004297157, 0.0009020684, 0.001387971, 0.001724662, 
    0.001836161, 0.001914496, 0.001936912, 0.001699325, 0.001502143, 
    0.00140803, 0.001545498, 0.002019594, 0.00346276, 0.005782628, 
    0.008145876, 0.0102145, 0.01200862, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;

 u_west =
  -0.0005609904, -0.0006586229, -0.0005458365, -0.0006437502, -0.0008264347, 
    -0.001240726, -0.00149311, -0.001744555, -0.001678442, -0.0008124625, 
    0.0005376131, 0.002128962, 0.003299844, 0.003907657, 0.004644471, 
    0.005593318, 0.006545128, 0.00658676, 0.005705373, 0.004862352, 
    0.004670639, 0.004483731, 0.004248674, 0.00417891, 0.003957627, 
    0.003788455, 0.00343842, 0.002796349, 0.002020997, 0.001817432, 
    0.001872291, 0.001793962, 0.001584719, 0.001317679, 0.001034577, 
    0.0008378435, 0.0007899673, 0.0007547764, 0.0007001892, 0.0006668972, 
    0.000622046, 0.0005451408, 0.0003694768, 0.0002152439, 0.0001655161, 
    0.0002379938, 0.0002908029, 0.0003434924, 0.0004227406, 0.0005177781, 
    0.0006134532, 0.0006490806, 0.000697, 0.0007674557, 0.0007923699,
  -0.002268772, -0.002094491, -0.001611534, -0.001354993, -0.001175552, 
    -0.001368385, -0.001610406, -0.001851574, -0.001781641, -0.001253594, 
    -0.0007174448, 0.0003763504, 0.002029681, 0.003678013, 0.004649907, 
    0.005547764, 0.006448317, 0.006620186, 0.00605169, 0.005518108, 
    0.005198789, 0.004791704, 0.00438867, 0.004383859, 0.004212396, 
    0.00403359, 0.003467388, 0.002784749, 0.002153763, 0.001998808, 
    0.001926495, 0.001729654, 0.001412344, 0.001094642, 0.0007954929, 
    0.0006029038, 0.0005673631, 0.000545234, 0.0004974427, 0.0004782897, 
    0.0004431194, 0.0003561109, 0.0001346256, -8.568779e-05, -0.0001575737, 
    -5.108913e-05, 4.942787e-05, 0.0001604984, 0.0002917872, 0.0004293114, 
    0.0005633826, 0.0006173665, 0.0006707107, 0.0007303578, 0.0007577727,
  -0.002328006, -0.002171454, -0.001752818, -0.001550904, -0.001349886, 
    -0.001496769, -0.001727493, -0.001957161, -0.001882299, -0.00134894, 
    -0.0008056561, 0.0002824719, 0.001911416, 0.003534956, 0.004500508, 
    0.00538804, 0.006275302, 0.006465845, 0.005955997, 0.005435517, 
    0.005077124, 0.004675973, 0.004278526, 0.004258771, 0.004079238, 
    0.003886586, 0.003377917, 0.002835893, 0.002363923, 0.00215691, 
    0.001820477, 0.001505053, 0.001184593, 0.0008847495, 0.0006018737, 
    0.0004175736, 0.000379132, 0.0003529387, 0.0003017138, 0.0002800889, 
    0.0002438267, 0.0001586124, -4.188328e-05, -0.0002413121, -0.0002788378, 
    -0.0001663925, -5.939563e-05, 6.324895e-05, 0.0002103664, 0.0003631743, 
    0.0005001089, 0.0005680818, 0.0006408991, 0.0007096694, 0.0007347957,
  -0.002347663, -0.002209293, -0.001823008, -0.001643233, -0.001461604, 
    -0.001606534, -0.001824787, -0.00204209, -0.001964798, -0.001436079, 
    -0.0008926894, 0.0001798964, 0.001783664, 0.003383056, 0.004339593, 
    0.005211824, 0.006083891, 0.006277151, 0.005786889, 0.005281103, 
    0.004920261, 0.004508918, 0.004101517, 0.004065006, 0.003880949, 
    0.003684831, 0.003319896, 0.002903529, 0.002437221, 0.001981, 
    0.001615084, 0.00130108, 0.0009949032, 0.000714063, 0.0004472455, 
    0.0002664152, 0.0002193803, 0.0001837703, 0.0001260423, 0.0001018239, 
    6.339161e-05, -1.87828e-05, -0.0001955682, -0.0003721388, -0.0003894617, 
    -0.0002662928, -0.0001482906, -9.898846e-06, 0.0001564603, 0.0003272766, 
    0.0004763241, 0.0005596325, 0.0006459834, 0.0007139161, 0.0007271148,
  -0.002334728, -0.002214993, -0.001857813, -0.001696975, -0.001534417, 
    -0.001678089, -0.001884948, -0.00209093, -0.00200917, -0.001478042, 
    -0.0009431688, 0.000102344, 0.001669114, 0.003238554, 0.004182924, 
    0.005037158, 0.005891242, 0.006082993, 0.005608054, 0.005118767, 
    0.004763839, 0.00434789, 0.003934775, 0.003879439, 0.003687537, 
    0.003481106, 0.003133747, 0.002695761, 0.002242374, 0.001799194, 
    0.001442653, 0.001136452, 0.0008397907, 0.0005706583, 0.000314486, 
    0.0001353905, 8.090687e-05, 3.6975e-05, -2.732931e-05, -5.451778e-05, 
    -9.483544e-05, -0.0001737985, -0.0003292523, -0.0004845122, 
    -0.0004882062, -0.0003533076, -0.0002231768, -7.010202e-05, 0.0001129089, 
    0.0003000287, 0.0004611756, 0.0005543645, 0.0006503906, 0.0007191408, 
    0.0007247951,
  -0.002290677, -0.002188819, -0.001866934, -0.00173093, -0.001590352, 
    -0.00173374, -0.00192805, -0.002121489, -0.002038182, -0.001514891, 
    -0.0009781882, 5.219354e-05, 0.001586132, 0.003122317, 0.004049445, 
    0.004881086, 0.005713137, 0.00590025, 0.005437824, 0.004960473, 
    0.004603404, 0.004182656, 0.003764538, 0.003691498, 0.003494178, 
    0.003283374, 0.002941068, 0.002513314, 0.002070572, 0.001642105, 
    0.001293701, 0.0009918816, 0.0007035761, 0.0004390551, 0.0001888285, 
    1.087199e-05, -4.949865e-05, -9.912236e-05, -0.0001661529, -0.0001930607, 
    -0.00023265, -0.0003048755, -0.0004367981, -0.0005709155, -0.0005619577, 
    -0.000416542, -0.0002725599, -9.937987e-05, 0.0001036441, 0.0003060243, 
    0.0004764411, 0.0005828983, 0.0006971968, 0.0007659189, 0.000755029,
  -0.002218324, -0.002134041, -0.001841241, -0.00172362, -0.001601733, 
    -0.001743206, -0.001924139, -0.002104261, -0.002013213, -0.0014869, 
    -0.0009681297, 2.302508e-05, 0.001511885, 0.003018558, 0.003930364, 
    0.004741079, 0.005552178, 0.005733913, 0.005282, 0.004816199, 
    0.004459858, 0.004034956, 0.003612684, 0.003522752, 0.003318859, 
    0.003100974, 0.002761849, 0.002344494, 0.001915078, 0.001501669, 
    0.001156019, 0.0008464859, 0.0005603423, 0.0003076339, 6.928042e-05, 
    -0.0001048239, -0.0001699558, -0.0002250924, -0.0002941303, 
    -0.0003185297, -0.0003547241, -0.0004172979, -0.0005209745, 
    -0.0006266999, -0.0005987384, -0.0004373559, -0.0002772987, 
    -8.942426e-05, 0.0001268534, 0.000342519, 0.0005192112, 0.0006296774, 
    0.0007474681, 0.0008077754, 0.000782082,
  -0.00215193, -0.002083774, -0.001817663, -0.001716912, -0.001612177, 
    -0.001751892, -0.00192055, -0.002088453, -0.001990299, -0.001458698, 
    -0.0009341459, 4.442147e-05, 0.001498017, 0.002964074, 0.003854922, 
    0.004639465, 0.005425292, 0.005597801, 0.005153205, 0.004697826, 
    0.004341076, 0.003908341, 0.003475709, 0.003366345, 0.003153603, 
    0.002927823, 0.002594901, 0.002189259, 0.001772388, 0.001362732, 
    0.001008252, 0.0007043626, 0.000427864, 0.0001870305, -4.042752e-05, 
    -0.000210997, -0.0002804981, -0.0003406939, -0.0004115737, -0.000433671, 
    -0.00046675, -0.0005204666, -0.0005982222, -0.0006778924, -0.0006324916, 
    -0.0004564566, -0.0002816474, -8.028813e-05, 0.0001481524, 0.0003760098, 
    0.0005584608, 0.0006726062, 0.0007936017, 0.0008474921, 0.0008118179,
  -0.002030284, -0.001981432, -0.001754093, -0.001679795, -0.001598626, 
    -0.001737847, -0.001891068, -0.002043535, -0.001938759, -0.001411916, 
    -0.0009019699, 6.467958e-05, 0.00148754, 0.002922024, 0.003794889, 
    0.00455465, 0.005315608, 0.005478787, 0.005040661, 0.004592503, 
    0.004230996, 0.003788463, 0.003346022, 0.00321826, 0.002997138, 
    0.002763883, 0.002434252, 0.002033443, 0.001618899, 0.001213965, 
    0.0008683437, 0.0005697972, 0.0003024302, 6.416046e-05, -0.0001615532, 
    -0.000331709, -0.0004047033, -0.0004666702, -0.0005344649, -0.0005494762, 
    -0.0005766977, -0.000618607, -0.0006659441, -0.0007176045, -0.0006545471, 
    -0.000463584, -0.0002707437, -4.77431e-05, 0.0001993057, 0.0004406579, 
    0.0006293426, 0.0007528992, 0.0008893862, 0.0009377951, 0.0008796112,
  -0.001902002, -0.001872723, -0.001678169, -0.001624697, -0.001564844, 
    -0.001702971, -0.001840677, -0.001977682, -0.001861302, -0.001324312, 
    -0.0008040208, 0.0001273539, 0.001500283, 0.002894125, 0.003745104, 
    0.00447737, 0.005211705, 0.005363884, 0.004931121, 0.00449139, 
    0.004126448, 0.003672404, 0.00321556, 0.003064976, 0.00283007, 
    0.002581417, 0.002251109, 0.00186108, 0.001458324, 0.001068187, 
    0.0007232102, 0.000410881, 0.0001432958, -8.443975e-05, -0.0002969096, 
    -0.0004611454, -0.000536636, -0.0006019105, -0.0006680555, -0.0006732338, 
    -0.0006897234, -0.0007153222, -0.000723965, -0.0007366237, -0.0006463678, 
    -0.0004297037, -0.0002112875, 3.10191e-05, 0.0002915295, 0.0005467415, 
    0.0007416097, 0.0008627336, 0.0009958764, 0.001026284, 0.0009460427,
  -0.001771514, -0.001762306, -0.001601342, -0.001568943, -0.001530659, 
    -0.00166768, -0.001789685, -0.001911045, -0.001782922, -0.001235664, 
    -0.0007038121, 0.0002175489, 0.001556508, 0.002914752, 0.003743266, 
    0.004443873, 0.005146389, 0.005282436, 0.00484945, 0.004410057, 
    0.004030855, 0.003557042, 0.003080645, 0.00290531, 0.002655386, 
    0.002392809, 0.002065786, 0.001686665, 0.001295837, 0.0008928221, 
    0.0005316331, 0.000231713, -2.16874e-05, -0.0002348085, -0.0004338769, 
    -0.0005921222, -0.0006701387, -0.0007387603, -0.0008032359, 
    -0.0007984642, -0.0008040942, -0.0008131884, -0.0007826763, 
    -0.0007558693, -0.0006380911, -0.0003954202, -0.0001511238, 0.0001107186, 
    0.0003848509, 0.0006540875, 0.000855213, 0.000973875, 0.001103634, 
    0.001115826, 0.001013265,
  -0.001616665, -0.001636087, -0.001521385, -0.001518341, -0.001508764, 
    -0.001647347, -0.001751444, -0.001854759, -0.001709799, -0.001146311, 
    -0.0005990994, 0.0003114541, 0.00161476, 0.002936124, 0.003741361, 
    0.004409168, 0.005078717, 0.005198049, 0.004764832, 0.004325791, 
    0.003931814, 0.003437519, 0.002940681, 0.002734522, 0.002464724, 
    0.002178626, 0.001840277, 0.001461106, 0.001066201, 0.0006759962, 
    0.0003331479, 4.608481e-05, -0.000192619, -0.0004001572, -0.000595745, 
    -0.0007539634, -0.0008365957, -0.0009071641, -0.0009642619, 
    -0.0009419293, -0.0009325797, -0.0009196683, -0.0008392973, 
    -0.0007655679, -0.0006163759, -0.0003444397, -6.733509e-05, 0.0002263963, 
    0.0005233973, 0.0008093824, 0.001017828, 0.00113993, 0.001279362, 
    0.001274306, 0.001139275,
  -0.001454623, -0.001504006, -0.001437691, -0.00146682, -0.001490072, 
    -0.001631595, -0.001715689, -0.00179908, -0.001635892, -0.001054494, 
    -0.0004877436, 0.0004169277, 0.001684676, 0.002968474, 0.00374796, 
    0.004379689, 0.005013147, 0.005110699, 0.004670505, 0.004224211, 
    0.003801443, 0.003269111, 0.002732744, 0.002493433, 0.002199918, 
    0.001891776, 0.001557033, 0.001193173, 0.0008152019, 0.0004491001, 
    9.743118e-05, -0.0001883304, -0.0004183533, -0.0006134624, -0.0007957517, 
    -0.000949726, -0.001038151, -0.001115761, -0.001169119, -0.001122373, 
    -0.001087265, -0.001040339, -0.000889124, -0.0007438821, -0.0005417735, 
    -0.0002178391, 0.0001107521, 0.0004383618, 0.0007529692, 0.001057663, 
    0.001273868, 0.001380292, 0.001502314, 0.001457229, 0.001280457,
  -0.001365998, -0.001449996, -0.001427172, -0.001479477, -0.001529706, 
    -0.001671241, -0.001731587, -0.00179061, -0.001599559, -0.000984559, 
    -0.0003807193, 0.0005266579, 0.001758903, 0.003005338, 0.003758269, 
    0.004352202, 0.004947662, 0.005020383, 0.004568745, 0.004111746, 
    0.003658295, 0.003089137, 0.002516414, 0.002242614, 0.001924426, 
    0.001586485, 0.001240446, 0.0008809664, 0.0005044806, 0.0001351889, 
    -0.0001880911, -0.0004471796, -0.0006556243, -0.0008353718, -0.001003826, 
    -0.001153384, -0.001247837, -0.001332772, -0.001382239, -0.001310095, 
    -0.001248191, -0.001165877, -0.0009409605, -0.0007213216, -0.0004641617, 
    -8.613183e-05, 0.0002960228, 0.0006588772, 0.0009918011, 0.001315958, 
    0.001540236, 0.001630349, 0.001745445, 0.001679206, 0.001461133,
  -0.001323486, -0.001444766, -0.001476524, -0.001562293, -0.001646257, 
    -0.001787277, -0.001813984, -0.001839549, -0.001615784, -0.000967602, 
    -0.0003290979, 0.0005902399, 0.001806598, 0.00302976, 0.003761909, 
    0.004324637, 0.004888295, 0.004934577, 0.004462709, 0.003985769, 
    0.003483921, 0.002855322, 0.002221218, 0.001898111, 0.001539721, 
    0.001165766, 0.0008252628, 0.0004889703, 0.0001380169, -0.0001917705, 
    -0.0004651087, -0.0006783342, -0.0008547218, -0.00102085, -0.00118369, 
    -0.001343576, -0.001462841, -0.001573331, -0.001622386, -0.001507423, 
    -0.001401999, -0.00126121, -0.0009203348, -0.0005885084, -0.0002489499, 
    0.000209809, 0.0006780411, 0.001105612, 0.001471104, 0.001819712, 
    0.002051143, 0.002120037, 0.002211428, 0.002067174, 0.001772599,
  -0.00137204, -0.001516271, -0.001572816, -0.001666914, -0.001763403, 
    -0.001888003, -0.00186363, -0.001837532, -0.001569042, -0.0008875799, 
    -0.0002288186, 0.0006745068, 0.0018471, 0.003048748, 0.003762403, 
    0.004297663, 0.004833712, 0.004853586, 0.004356637, 0.003855431, 
    0.003301702, 0.002618823, 0.001932643, 0.001567094, 0.001170657, 
    0.000760795, 0.0004286149, 0.0001203936, -0.0001974072, -0.0004653252, 
    -0.0006865278, -0.000864394, -0.001021549, -0.001190879, -0.001357452, 
    -0.001530619, -0.001675015, -0.001812032, -0.001862542, -0.001703264, 
    -0.001552005, -0.001350393, -0.0008858237, -0.0004289091, 5.172678e-06, 
    0.000556903, 0.001116655, 0.001598562, 0.001984504, 0.002356157, 
    0.002593599, 0.002622873, 0.002689391, 0.002503257, 0.002143057,
  -0.001467527, -0.001625933, -0.001696076, -0.001785365, -0.001876613, 
    -0.001969687, -0.00188066, -0.001790212, -0.001462784, -0.0007238194, 
    -3.640682e-06, 0.0009378786, 0.002121171, 0.003316565, 0.004019664, 
    0.004541792, 0.00506498, 0.005054102, 0.00451117, 0.003974019, 
    0.003348545, 0.002570041, 0.001781027, 0.001343742, 0.0008840176, 
    0.0004132345, 8.000225e-05, -0.0002032694, -0.0004944089, -0.0006718964, 
    -0.0007428413, -0.0008236087, -0.000932758, -0.00110271, -0.001287356, 
    -0.001505911, -0.001721895, -0.001935332, -0.002010524, -0.001791251, 
    -0.001575237, -0.001282832, -0.0006375894, -4.794052e-06, 0.0005591321, 
    0.001235818, 0.001928063, 0.002501822, 0.00292524, 0.003323943, 
    0.00356773, 0.00355784, 0.003580779, 0.003278635, 0.002807974,
  -0.001152911, -0.001272433, -0.001304973, -0.001368077, -0.001428614, 
    -0.001462625, -0.001279406, -0.001095434, -0.0007064187, 5.156579e-05, 
    0.0007533177, 0.001640329, 0.002764046, 0.00393428, 0.00461961, 
    0.005129111, 0.005641858, 0.005590414, 0.004982981, 0.004409038, 
    0.003717976, 0.002846637, 0.001950802, 0.001433817, 0.0008957387, 
    0.0003555046, 3.952651e-05, -0.0001972736, -0.0004280784, -0.0005191588, 
    -0.0005713596, -0.0006316153, -0.0006937177, -0.0008663958, -0.001081842, 
    -0.001364898, -0.001674634, -0.001987819, -0.002095815, -0.001805539, 
    -0.001512004, -0.001112421, -0.0002642725, 0.0005631353, 0.001267534, 
    0.002074432, 0.002909142, 0.003583348, 0.004043823, 0.004463895, 
    0.004711568, 0.004661722, 0.004663704, 0.004284719, 0.003717132,
  -0.0002496155, -0.0003144749, -0.0003200094, -0.0003839788, -0.0004289189, 
    -0.0004053626, -0.000123569, 0.0001570409, 0.000598392, 0.00135044, 
    0.001986353, 0.002768578, 0.003838637, 0.005047556, 0.005744185, 
    0.006270904, 0.006800196, 0.006717917, 0.006030574, 0.005369791, 
    0.004523392, 0.003473839, 0.002446897, 0.001834932, 0.001201838, 
    0.0005798074, 0.0002876504, 0.0001079251, -4.452087e-05, 3.908102e-05, 
    0.0001496953, 0.0001846448, 7.716544e-05, -0.0002466761, -0.0006044185, 
    -0.001019005, -0.001466173, -0.001916118, -0.002063006, -0.00166295, 
    -0.001260264, -0.0007170737, 0.0004125765, 0.001525777, 0.002432846, 
    0.003407481, 0.00440417, 0.005151401, 0.005606976, 0.006030515, 
    0.006274218, 0.006133076, 0.006033052, 0.005511769, 0.004830108,
  0.001321838, 0.001321274, 0.001351437, 0.001299866, 0.001307298, 
    0.001393908, 0.001750587, 0.002106343, 0.002623079, 0.003483113, 
    0.004252637, 0.005170334, 0.006314926, 0.007538878, 0.008234731, 
    0.008779122, 0.00932899, 0.009175304, 0.008331983, 0.007548064, 
    0.006512971, 0.005219412, 0.00388949, 0.003051789, 0.002234581, 
    0.00142602, 0.00106284, 0.0008740572, 0.000706573, 0.0009470508, 
    0.001200267, 0.001314776, 0.001170433, 0.0006623816, 9.343854e-05, 
    -0.0005310017, -0.001182882, -0.001838087, -0.002011464, -0.001389401, 
    -0.000762313, 4.400044e-05, 0.001591989, 0.003112378, 0.00428457, 
    0.005429238, 0.006610722, 0.007449808, 0.007878872, 0.008258015, 
    0.00847512, 0.008235491, 0.008054051, 0.007397009, 0.006582706,
  0.004142272, 0.004160529, 0.004232593, 0.004165983, 0.00412806, 0.00424886, 
    0.004722301, 0.00519408, 0.005801763, 0.006758073, 0.007573293, 
    0.008502451, 0.009665754, 0.0109487, 0.0116618, 0.01223438, 0.01281563, 
    0.01256118, 0.01149322, 0.01051771, 0.009205991, 0.007565877, 
    0.005869613, 0.004765391, 0.003736621, 0.002724069, 0.002331398, 
    0.002195404, 0.002098525, 0.00231453, 0.0025717, 0.002732116, 
    0.002489561, 0.001700207, 0.0008252346, -7.627594e-05, -0.000961008, 
    -0.001845804, -0.002006773, -0.001044409, -7.684524e-05, 0.001099216, 
    0.003179441, 0.005219147, 0.006712892, 0.008018608, 0.009377514, 
    0.01027887, 0.01062798, 0.01090862, 0.0110766, 0.01070798, 0.0104131, 
    0.009591044, 0.008649814,
  0.00728587, 0.007242734, 0.007252094, 0.007122366, 0.007025502, 
    0.007192038, 0.00784178, 0.00849103, 0.009259471, 0.01041631, 0.01139692, 
    0.01244405, 0.01370897, 0.01511616, 0.01587251, 0.01648424, 0.01710692, 
    0.01672285, 0.01535935, 0.01410573, 0.01240227, 0.0102992, 0.008127203, 
    0.006701444, 0.005438393, 0.004194241, 0.00377776, 0.003718587, 
    0.003714273, 0.00405423, 0.004285428, 0.004391749, 0.003977995, 
    0.002796927, 0.001508747, 0.0002533307, -0.0008971574, -0.002039271, 
    -0.002134707, -0.000687312, 0.0007593111, 0.00243057, 0.00518406, 
    0.007885642, 0.009769142, 0.01122272, 0.01274148, 0.01365631, 0.0138522, 
    0.01396661, 0.01405872, 0.01352458, 0.01307321, 0.01204858, 0.01097025,
  0.01020649, 0.01003785, 0.009957976, 0.00979148, 0.009651395, 0.009896474, 
    0.0107928, 0.01169058, 0.01269258, 0.01414959, 0.01542616, 0.01671531, 
    0.01817504, 0.01977507, 0.02059676, 0.02124977, 0.02191434, 0.02136854, 
    0.01963926, 0.0180134, 0.01579716, 0.0131276, 0.01039058, 0.008628069, 
    0.007142528, 0.005676001, 0.005281454, 0.005347756, 0.00548277, 
    0.005939018, 0.006187861, 0.006286448, 0.005559165, 0.003845056, 
    0.002022345, 0.0003199265, -0.001145214, -0.002585124, -0.0025539, 
    -0.0004698407, 0.001596117, 0.003893804, 0.007480166, 0.01100758, 
    0.01335224, 0.01494109, 0.01659852, 0.01746977, 0.01743167, 0.01730723, 
    0.01729722, 0.01657681, 0.01594766, 0.01470294, 0.01348132,
  0.01250105, 0.01217014, 0.01199682, 0.01183295, 0.01168422, 0.01204612, 
    0.01323751, 0.01443154, 0.01571819, 0.0175534, 0.01923149, 0.02086195, 
    0.02257818, 0.02440598, 0.02528388, 0.02595507, 0.02663645, 0.02589241, 
    0.02374742, 0.02168683, 0.01889175, 0.01561994, 0.01228667, 0.01024521, 
    0.008600286, 0.006970521, 0.006689772, 0.00696466, 0.007323981, 
    0.007908966, 0.008153834, 0.008245395, 0.007125245, 0.004697222, 
    0.002156902, -0.0001250562, -0.00200074, -0.003844667, -0.003657511, 
    -0.000789775, 0.002053719, 0.005135786, 0.009744562, 0.01430435, 
    0.0172205, 0.01899058, 0.02081153, 0.02159579, 0.0212596, 0.02085169, 
    0.02073482, 0.01983328, 0.01901767, 0.0175424, 0.016164,
  0.0139251, 0.01338024, 0.01308656, 0.01293556, 0.01279095, 0.01327175, 
    0.01475495, 0.01624128, 0.01783451, 0.02010669, 0.02227465, 0.02436893, 
    0.02646143, 0.02860824, 0.0295417, 0.03023518, 0.03093398, 0.02995452, 
    0.02731892, 0.02474953, 0.02131039, 0.01740691, 0.0134467, 0.01125334, 
    0.009556008, 0.007869516, 0.007859452, 0.008485561, 0.009203814, 
    0.009937963, 0.01014474, 0.01020327, 0.008600861, 0.005269974, 
    0.001803413, -0.001104426, -0.003334397, -0.005520456, -0.005116249, 
    -0.001417532, 0.002243463, 0.00606982, 0.01157239, 0.01707955, 
    0.02049928, 0.02242673, 0.02434423, 0.02496122, 0.02428704, 0.02362803, 
    0.02341926, 0.02227944, 0.02106586, 0.01919905, 0.01761203,
  0.01404635, 0.01315614, 0.01257657, 0.01236138, 0.01214143, 0.01259898, 
    0.01420097, 0.01580456, 0.0175211, 0.02017459, 0.02288326, 0.02560681, 
    0.02830177, 0.03094049, 0.03209512, 0.03299864, 0.03389431, 0.03285298, 
    0.02987106, 0.02687916, 0.02277216, 0.01825693, 0.01373901, 0.01148097, 
    0.00976803, 0.008043184, 0.008276824, 0.00914788, 0.01002494, 0.01044426, 
    0.01001065, 0.009550859, 0.007416418, 0.003646055, -0.0001684608, 
    -0.003221247, -0.005294006, -0.007354315, -0.006681263, -0.002518085, 
    0.001644893, 0.005847202, 0.01138783, 0.01690653, 0.0202857, 0.02214491, 
    0.0240331, 0.0246135, 0.02385102, 0.02304977, 0.02259613, 0.02146223, 
    0.02042694, 0.01875647, 0.0172986,
  0.01379195, 0.01279314, 0.01198582, 0.01163403, 0.01128286, 0.01164273, 
    0.0133854, 0.01513041, 0.01688171, 0.01949868, 0.02210277, 0.02462176, 
    0.02708306, 0.02956112, 0.03067919, 0.03144636, 0.03222423, 0.03115426, 
    0.02822267, 0.02522484, 0.02104059, 0.01659639, 0.01219982, 0.01041749, 
    0.009230777, 0.008083146, 0.008874104, 0.01002608, 0.01123435, 
    0.01169802, 0.01073128, 0.009756887, 0.00742973, 0.003766917, 
    -6.983603e-05, -0.002935242, -0.004665328, -0.006491284, -0.005632279, 
    -0.001312173, 0.003121383, 0.007628303, 0.01350696, 0.01934572, 
    0.0231675, 0.02509544, 0.02711505, 0.02806406, 0.02779846, 0.0274161, 
    0.02703264, 0.0261087, 0.02540147, 0.02381076, 0.02241537,
  0.01453415, 0.01360906, 0.01285351, 0.01257156, 0.01229263, 0.01287913, 
    0.01506443, 0.01725256, 0.01947454, 0.02247662, 0.02534148, 0.02789548, 
    0.03025917, 0.03271591, 0.03367934, 0.03415971, 0.03464347, 0.03328348, 
    0.03010322, 0.02704125, 0.02340695, 0.01979369, 0.01616097, 0.01538034, 
    0.01501058, 0.01474931, 0.01628103, 0.01774745, 0.0193672, 0.02031484, 
    0.01982593, 0.01887635, 0.01589559, 0.01150473, 0.007183644, 0.003913653, 
    0.001770194, -0.0004950881, 0.0003368162, 0.004959586, 0.009720738, 
    0.01455745, 0.02056701, 0.02651589, 0.03057966, 0.03276336, 0.03506478, 
    0.03629345, 0.03626584, 0.03609388, 0.03578024, 0.03505584, 0.03455787, 
    0.0329119, 0.03162368,
  0.0164004, 0.01566935, 0.01525056, 0.0153594, 0.01547035, 0.01672835, 
    0.01979678, 0.02286844, 0.02599136, 0.02963259, 0.0331236, 0.0362963, 
    0.03926531, 0.04234382, 0.04398115, 0.04518144, 0.04638417, 0.04550292, 
    0.04256886, 0.03978091, 0.03632201, 0.03293354, 0.02950085, 0.02900481, 
    0.02863119, 0.0283529, 0.02995937, 0.03120062, 0.03257424, 0.03323869, 
    0.03275257, 0.03188267, 0.02868233, 0.02372653, 0.01888762, 0.01492724, 
    0.01198722, 0.008916623, 0.009530141, 0.01447424, 0.01956265, 0.0248985, 
    0.03156339, 0.03816751, 0.04268201, 0.04513545, 0.04767185, 0.04902775, 
    0.04904427, 0.04892318, 0.04859071, 0.0477416, 0.04711683, 0.04521457, 
    0.04402607,
  0.02181502, 0.0215111, 0.02187769, 0.02279733, 0.02372098, 0.02619654, 
    0.03069948, 0.03520325, 0.03971228, 0.04447234, 0.04913111, 0.05354426, 
    0.0577927, 0.06211736, 0.06493701, 0.06751858, 0.07009926, 0.07003749, 
    0.06735565, 0.06476105, 0.06099806, 0.05738649, 0.05375024, 0.05348985, 
    0.05266349, 0.05189368, 0.0531467, 0.0537358, 0.05440331, 0.05444378, 
    0.05379154, 0.05264886, 0.04869435, 0.04265955, 0.03662461, 0.03157401, 
    0.02731225, 0.02305028, 0.02329031, 0.0286999, 0.03410973, 0.03995356, 
    0.04762807, 0.05530252, 0.06040578, 0.06309547, 0.06578532, 0.06697825, 
    0.06667405, 0.06636968, 0.06616534, 0.06522677, 0.06428851, 0.06178953, 
    0.0604593,
  -0.0008747782, -0.000958401, -0.001023069, -0.001352619, -0.001745985, 
    -0.002247806, -0.002605177, -0.002961029, -0.002940941, -0.002099733, 
    -0.0007730495, 0.0007509969, 0.001861318, 0.00242334, 0.003007539, 
    0.00376294, 0.004515049, 0.004616299, 0.004059121, 0.003529087, 
    0.003442943, 0.003378175, 0.003318374, 0.003434847, 0.003454896, 
    0.003588392, 0.003556144, 0.003101567, 0.002467429, 0.002304113, 
    0.00238289, 0.002346527, 0.002226546, 0.00211534, 0.002014439, 
    0.001940233, 0.001949816, 0.001941845, 0.00181681, 0.001652266, 
    0.001508349, 0.001317319, 0.000964693, 0.0006396301, 0.0004636727, 
    0.0004320439, 0.000382011, 0.0003308196, 0.0003048193, 0.0002964148, 
    0.0003001092, 0.0002309096, 0.0001467993, 0.0001027739, 0.0001216497,
  -0.002029441, -0.001983996, -0.001837221, -0.001902707, -0.002026235, 
    -0.002362324, -0.002696123, -0.003028541, -0.003002571, -0.002517577, 
    -0.00202687, -0.001050044, 0.0004236917, 0.00189962, 0.002796439, 
    0.003582094, 0.004364755, 0.004603624, 0.004291816, 0.004004711, 
    0.003919337, 0.003834083, 0.003753289, 0.004003142, 0.004121314, 
    0.004231309, 0.003835696, 0.003208029, 0.002643467, 0.00253861, 
    0.002530539, 0.002414078, 0.002222104, 0.002061525, 0.001916385, 
    0.001821655, 0.001845278, 0.001882417, 0.001799038, 0.001644439, 
    0.001473706, 0.001238822, 0.0008154706, 0.0003928467, 0.0001724431, 
    0.0001574269, 0.0001367439, 0.0001279788, 0.0001400295, 0.0001582024, 
    0.0001759883, 0.0001220678, 6.506255e-05, 7.359863e-05, 0.0001197009,
  -0.002086224, -0.002060767, -0.001968637, -0.002074097, -0.002181033, 
    -0.002474428, -0.002782724, -0.003089344, -0.003056661, -0.002572981, 
    -0.002082037, -0.001125486, 0.0003029188, 0.001732699, 0.00261309, 
    0.003386124, 0.004158654, 0.004422017, 0.00417176, 0.003910342, 
    0.003803465, 0.003726399, 0.00365341, 0.003887828, 0.003992189, 
    0.004082579, 0.003744483, 0.003276254, 0.002885544, 0.002742372, 
    0.00246903, 0.002214062, 0.002009326, 0.00186126, 0.001727313, 
    0.001639183, 0.001657679, 0.001688307, 0.001602369, 0.00144501, 
    0.001272905, 0.001041483, 0.0006421325, 0.000243442, 5.848712e-05, 
    4.780958e-05, 3.195746e-05, 3.122866e-05, 5.374871e-05, 8.185738e-05, 
    8.890496e-05, 4.916552e-05, 1.053169e-05, 4.796045e-05, 0.000101238,
  -0.002103638, -0.002098243, -0.002038374, -0.0021618, -0.002284291, 
    -0.002566833, -0.002849022, -0.003129582, -0.003092888, -0.002621229, 
    -0.002134646, -0.001207021, 0.0001728053, 0.001556282, 0.002419324, 
    0.003177661, 0.003935519, 0.004208128, 0.003989881, 0.003755494, 
    0.003653313, 0.003569781, 0.003490873, 0.003707917, 0.003800898, 
    0.003881031, 0.003689445, 0.003358938, 0.002979894, 0.002578231, 
    0.002275371, 0.002025822, 0.001836342, 0.001705134, 0.001584397, 
    0.001498854, 0.001505576, 0.001523368, 0.001430987, 0.00126998, 
    0.001095116, 0.0008675136, 0.0004939771, 0.0001202475, -4.674084e-05, 
    -5.007811e-05, -5.852919e-05, -4.975221e-05, -1.637195e-05, 2.199606e-05, 
    3.676125e-05, 1.134707e-05, -1.413702e-05, 2.451369e-05, 6.866513e-05,
  -0.00208863, -0.002103438, -0.002071701, -0.002208277, -0.002343982, 
    -0.002615472, -0.002872643, -0.003128308, -0.003084622, -0.002616612, 
    -0.002147628, -0.001263725, 5.639076e-05, 0.001388749, 0.00223115, 
    0.002971895, 0.003712199, 0.003989489, 0.00379858, 0.003592753, 
    0.003503382, 0.003418748, 0.003338017, 0.003536227, 0.003615147, 
    0.003678793, 0.003503758, 0.003154235, 0.002791087, 0.002404042, 
    0.002118461, 0.001883651, 0.001701649, 0.001577304, 0.001462634, 
    0.001377216, 0.001373732, 0.001380474, 0.001282082, 0.001117424, 
    0.0009399655, 0.0007160015, 0.000365742, 1.529942e-05, -0.0001412018, 
    -0.0001368263, -0.0001371709, -0.0001192836, -7.635767e-05, 
    -2.883057e-05, -4.380547e-06, -1.992822e-05, -3.552001e-05, 5.311992e-06, 
    4.327691e-05,
  -0.002041423, -0.002075125, -0.002077405, -0.002233734, -0.002386539, 
    -0.002649173, -0.002881216, -0.003111803, -0.003065071, -0.002612557, 
    -0.002146865, -0.001291441, -2.649365e-05, 0.001249651, 0.002064708, 
    0.002783332, 0.003502056, 0.003781027, 0.003614706, 0.003432697, 
    0.003349083, 0.003264004, 0.003182549, 0.003363121, 0.003430259, 
    0.00348322, 0.003311028, 0.002974478, 0.002625869, 0.002258928, 
    0.001985499, 0.001758802, 0.001583366, 0.00146242, 0.001352879, 
    0.001269501, 0.001257996, 0.00125589, 0.001153709, 0.0009870795, 
    0.0008091902, 0.0005913576, 0.0002644586, -6.458382e-05, -0.0002121069, 
    -0.0002013809, -0.0001923686, -0.0001608751, -0.0001054809, 
    -4.951199e-05, -1.796085e-05, -2.157196e-05, -2.138333e-05, 1.913387e-05, 
    4.348567e-05,
  -0.001964902, -0.002016729, -0.002045312, -0.002212795, -0.002376992, 
    -0.002628744, -0.00283576, -0.00304142, -0.002984683, -0.002536645, 
    -0.002098956, -0.001298923, -0.0001006528, 0.001125378, 0.001915687, 
    0.002613553, 0.003311514, 0.003590701, 0.003445956, 0.003286609, 
    0.003211026, 0.003125705, 0.003044343, 0.003208735, 0.003263658, 
    0.003304028, 0.003133784, 0.002811495, 0.002479518, 0.002129455, 
    0.001863288, 0.001636829, 0.001465344, 0.001353293, 0.001252456, 
    0.001172715, 0.001154457, 0.00114494, 0.001041018, 0.0008748188, 
    0.0006981473, 0.0004879222, 0.0001876961, -0.0001145304, -0.0002483966, 
    -0.0002275866, -0.0002083637, -0.0001682491, -0.0001059343, 
    -4.309534e-05, -7.13207e-06, -6.495685e-06, -2.301512e-06, 3.150152e-05, 
    4.367244e-05,
  -0.001894681, -0.001963142, -0.002015861, -0.002193581, -0.00236823, 
    -0.002609997, -0.002794047, -0.002976833, -0.002910914, -0.002464, 
    -0.00202675, -0.00125268, -0.0001110826, 0.001052478, 0.001810999, 
    0.002482548, 0.00315513, 0.003430381, 0.003303573, 0.00316507, 
    0.003096734, 0.003008705, 0.002922117, 0.00306838, 0.003108554, 
    0.003135168, 0.002969385, 0.002661812, 0.002345219, 0.002002362, 
    0.001735379, 0.001519334, 0.001356447, 0.001253149, 0.001160298, 
    0.001083895, 0.001059439, 0.001043122, 0.0009376025, 0.0007717986, 
    0.0005962446, 0.0003930008, 0.0001172521, -0.0001603658, -0.0002816991, 
    -0.0002516352, -0.0002230422, -0.000175016, -0.0001063504, -3.720686e-05, 
    2.805371e-06, 7.339652e-06, 1.520974e-05, 4.384723e-05, 4.696667e-05,
  -0.001768961, -0.001856216, -0.00194337, -0.002139757, -0.002330518, 
    -0.002563652, -0.002721706, -0.002878584, -0.002804471, -0.002371482, 
    -0.001958386, -0.001208898, -0.0001181407, 0.0009930877, 0.00172268, 
    0.002369028, 0.003016338, 0.003287136, 0.003177022, 0.003056024, 
    0.002990805, 0.002897929, 0.002806393, 0.002935492, 0.002961702, 
    0.00297529, 0.002811472, 0.002512505, 0.00220259, 0.001867861, 
    0.001614272, 0.001408087, 0.001253341, 0.001152431, 0.001062991, 
    0.0009901779, 0.0009611555, 0.000940617, 0.000836315, 0.0006735108, 
    0.0005012159, 0.0003066739, 5.763123e-05, -0.0001951259, -0.0003045007, 
    -0.0002652722, -0.0002248694, -0.0001624778, -8.21572e-05, -5.478774e-06, 
    3.934098e-05, 5.233115e-05, 7.36963e-05, 9.580576e-05, 7.841572e-05,
  -0.001636619, -0.001742794, -0.001857595, -0.002065327, -0.002267835, 
    -0.00249113, -0.002623739, -0.002755259, -0.002667115, -0.002231453, 
    -0.001815412, -0.001117895, -9.939347e-05, 0.0009496092, 0.001645757, 
    0.002263881, 0.002883983, 0.003148474, 0.003053725, 0.002951062, 
    0.002890006, 0.002790949, 0.002690708, 0.002799598, 0.002806698, 
    0.002799806, 0.002634207, 0.00234931, 0.00205427, 0.001736062, 
    0.001488571, 0.001276936, 0.001124618, 0.001034572, 0.0009579312, 
    0.0008930301, 0.0008604933, 0.0008358142, 0.0007332656, 0.0005760684, 
    0.0004100809, 0.0002263213, 1.010691e-05, -0.000209558, -0.0003005684, 
    -0.0002445592, -0.0001874511, -0.0001130169, -2.503759e-05, 5.955091e-05, 
    0.0001095893, 0.0001214838, 0.0001411682, 0.0001467206, 0.0001092331,
  -0.00150219, -0.00162773, -0.001770798, -0.001990012, -0.002204405, 
    -0.002417744, -0.002524607, -0.002630465, -0.002528123, -0.002089757, 
    -0.001669484, -0.000995736, -3.209687e-05, 0.0009596591, 0.001619566, 
    0.002204207, 0.002790671, 0.003042679, 0.002956888, 0.002863818, 
    0.002797232, 0.002685006, 0.002571686, 0.002658919, 0.002645304, 
    0.002618809, 0.002454832, 0.002184173, 0.001904185, 0.001577074, 
    0.001322273, 0.001129201, 0.000991341, 0.0009153111, 0.0008516208, 
    0.0007947263, 0.0007586331, 0.0007297642, 0.0006289898, 0.0004774662, 
    0.0003178613, 0.0001450124, -3.7983e-05, -0.0002241619, -0.0002965894, 
    -0.0002235997, -0.0001495875, -6.296739e-05, 3.276179e-05, 0.0001253545, 
    0.0001806736, 0.0001914593, 0.0002094431, 0.0001982413, 0.0001404171,
  -0.001348134, -0.001500168, -0.001681117, -0.001916637, -0.002147083, 
    -0.002351868, -0.002430734, -0.002508547, -0.00238601, -0.001940225, 
    -0.001514249, -0.0008680261, 3.762735e-05, 0.0009700715, 0.001592429, 
    0.00214238, 0.002693993, 0.002933067, 0.002856557, 0.002773426, 
    0.00270111, 0.00257524, 0.002448196, 0.002508183, 0.00246911, 
    0.002413892, 0.002237886, 0.001971579, 0.001692181, 0.001380029, 
    0.001149979, 0.0009761386, 0.0008532585, 0.0007853258, 0.0007301314, 
    0.0006797602, 0.0006390163, 0.0006065992, 0.0005106158, 0.0003690941, 
    0.0002185515, 5.99128e-05, -8.22623e-05, -0.0002298687, -0.0002813549, 
    -0.0001891463, -9.295101e-05, 1.566315e-05, 0.0001266608, 0.0002295035, 
    0.0002915779, 0.0003062155, 0.0003334244, 0.0003031374, 0.000212209,
  -0.001186923, -0.00136668, -0.001587286, -0.001840785, -0.002089719, 
    -0.002286389, -0.002335082, -0.002382829, -0.002237907, -0.001781901, 
    -0.001343714, -0.0007163303, 0.0001323431, 0.001004756, 0.001584536, 
    0.002094571, 0.002606452, 0.002825601, 0.002749678, 0.002667208, 
    0.002574913, 0.00241876, 0.002259855, 0.00229246, 0.002224149, 
    0.002141346, 0.001966986, 0.001719597, 0.001460468, 0.001173833, 
    0.0009441361, 0.0007814978, 0.0006719502, 0.0006222339, 0.0005855961, 
    0.0005462046, 0.0005001456, 0.0004615476, 0.0003688184, 0.0002419508, 
    0.0001070012, -3.070126e-05, -0.0001161731, -0.0002065301, -0.0002215143, 
    -9.270055e-05, 3.97073e-05, 0.0001715134, 0.0002936834, 0.0004085115, 
    0.0004788821, 0.0004815938, 0.0004956262, 0.0004263026, 0.0002944881,
  -0.00110537, -0.001315831, -0.001568849, -0.001828996, -0.002088601, 
    -0.002273385, -0.002289338, -0.002303872, -0.002125835, -0.001642884, 
    -0.001174747, -0.0005585123, 0.0002345005, 0.001048484, 0.001584544, 
    0.002052693, 0.002522472, 0.002718029, 0.002637301, 0.002550816, 
    0.00243642, 0.002251383, 0.002063914, 0.00206803, 0.001969301, 
    0.00185154, 0.001664965, 0.001426311, 0.001172762, 0.0008852492, 
    0.0006932423, 0.0005661524, 0.0004814191, 0.0004525633, 0.0004352308, 
    0.0004072621, 0.0003556736, 0.0003106454, 0.0002213016, 0.000109679, 
    -9.04862e-06, -0.0001249703, -0.0001514517, -0.00018225, -0.0001592599, 
    7.635596e-06, 0.0001777167, 0.0003336502, 0.0004674431, 0.00059474, 
    0.0006737413, 0.000664046, 0.0006741998, 0.0005816796, 0.0004078671,
  -0.001073775, -0.001316581, -0.001612197, -0.001887815, -0.002162956, 
    -0.002334531, -0.002309754, -0.002283753, -0.002066782, -0.001555756, 
    -0.00105756, -0.0004368109, 0.0003269255, 0.001102552, 0.001601145, 
    0.002033058, 0.002466141, 0.00263384, 0.002535365, 0.002432397, 
    0.002275948, 0.002038485, 0.001796015, 0.001759383, 0.001615344, 
    0.00145619, 0.001271905, 0.00105873, 0.0008327138, 0.000584444, 
    0.0004520885, 0.000381476, 0.0003357347, 0.0003365833, 0.0003435398, 
    0.0003233875, 0.000251642, 0.0001842464, 9.104154e-05, 1.931109e-06, 
    -9.205595e-05, -0.0001739821, -0.0001111726, -5.570977e-05, 2.41429e-05, 
    0.0002495275, 0.0004827902, 0.0006868666, 0.0008445597, 0.0009887597, 
    0.001079431, 0.0010547, 0.001048148, 0.000879191, 0.0006296312,
  -0.001132379, -0.00139097, -0.001699527, -0.00196651, -0.002236859, 
    -0.002380858, -0.00230341, -0.00222442, -0.001955947, -0.001413051, 
    -0.0008956312, -0.0002944238, 0.0004159077, 0.001159593, 0.001625008, 
    0.002025213, 0.002426409, 0.002565757, 0.002442594, 0.002315659, 
    0.002110714, 0.001825058, 0.001536744, 0.001466891, 0.001279679, 
    0.001079755, 0.0009011077, 0.0007177189, 0.0005257639, 0.0003370323, 
    0.0002681973, 0.000244036, 0.0002256188, 0.0002403162, 0.0002601535, 
    0.0002426656, 0.00015023, 6.143944e-05, -3.467254e-05, -9.923884e-05, 
    -0.0001678913, -0.0002152911, -5.672246e-05, 9.563116e-05, 0.0002419427, 
    0.0005357962, 0.0008363226, 0.001079576, 0.001251001, 0.001411007, 
    0.001512911, 0.001457311, 0.001433637, 0.001221106, 0.0009056347,
  -0.001237005, -0.00150172, -0.001812249, -0.002058484, -0.002307485, 
    -0.0024107, -0.002272237, -0.002132503, -0.00179894, -0.001198928, 
    -0.0006199871, 2.519678e-05, 0.0007575736, 0.001503675, 0.001951341, 
    0.002337574, 0.002725088, 0.002829302, 0.002652762, 0.002483889, 
    0.002203372, 0.001822202, 0.001429997, 0.001297924, 0.001040158, 
    0.0007719219, 0.0005855674, 0.0004251624, 0.0002577217, 0.0001542451, 
    0.0002452305, 0.0003297599, 0.0003725617, 0.000420469, 0.0004593224, 
    0.0004307217, 0.000280226, 0.0001269118, 5.882982e-07, -3.926122e-05, 
    -7.667326e-05, -7.696007e-05, 0.0002158518, 0.000498471, 0.0007338383, 
    0.001119718, 0.001519127, 0.001831987, 0.002031576, 0.002210465, 
    0.002331886, 0.002250492, 0.002197828, 0.001873919, 0.00145169,
  -0.000919334, -0.001136646, -0.001404421, -0.001615221, -0.0018237, 
    -0.001864953, -0.00164845, -0.001431581, -0.001028476, -0.0004006574, 
    0.0001689707, 0.0007782184, 0.001475326, 0.00221723, 0.00264596, 
    0.003021535, 0.003400592, 0.003458796, 0.003205617, 0.002989668, 
    0.002634157, 0.002157348, 0.001654306, 0.001453561, 0.001108333, 
    0.0007615783, 0.0005833449, 0.0004629688, 0.0003481838, 0.0003204474, 
    0.0004437742, 0.0005617787, 0.0006663109, 0.0007524196, 0.0008070663, 
    0.0007576231, 0.000532936, 0.0002965512, 0.0001303367, 0.0001192358, 
    0.0001203227, 0.000175886, 0.000616666, 0.001040264, 0.001370212, 
    0.001850759, 0.002356186, 0.002745433, 0.002972537, 0.003164814, 
    0.003307171, 0.003201602, 0.003143277, 0.002745512, 0.002231383,
  -2.291061e-05, -0.0001795268, -0.0004189055, -0.0006224132, -0.0008073931, 
    -0.0007900362, -0.0004939965, -0.0001995022, 0.0002683997, 0.0009050889, 
    0.001422032, 0.001951804, 0.002632803, 0.00345297, 0.003902179, 
    0.004302825, 0.00470623, 0.004728222, 0.00437631, 0.004053918, 0.0035213, 
    0.002855882, 0.002212351, 0.001927414, 0.001475647, 0.001035138, 
    0.0008673567, 0.0007924154, 0.0007420994, 0.0008691779, 0.001166464, 
    0.001395747, 0.001484373, 0.001484902, 0.001460487, 0.001336062, 
    0.001003938, 0.0006625095, 0.0004571911, 0.000502454, 0.0005574143, 
    0.0006842415, 0.001331415, 0.001964962, 0.0024343, 0.003036292, 
    0.003658015, 0.004094967, 0.004310706, 0.004498831, 0.004663649, 
    0.004492472, 0.004358772, 0.00382852, 0.003208496,
  0.001525037, 0.001436299, 0.001230655, 0.001046041, 0.0009176478, 
    0.0009976442, 0.001349136, 0.001699423, 0.002261415, 0.003028741, 
    0.00370275, 0.004415838, 0.005242982, 0.006146433, 0.006614111, 
    0.007041146, 0.007474018, 0.007410021, 0.006864696, 0.00638312, 
    0.005621931, 0.004692207, 0.003723761, 0.003225922, 0.002571804, 
    0.001926483, 0.001668492, 0.001567532, 0.001485799, 0.001741903, 
    0.002195241, 0.002527567, 0.002628755, 0.002556725, 0.002440884, 
    0.002214692, 0.001735799, 0.001242198, 0.0009974522, 0.001168758, 
    0.001357373, 0.001629138, 0.002571482, 0.003491049, 0.00413191, 
    0.004842691, 0.005586603, 0.00607635, 0.006253155, 0.006386804, 
    0.00656784, 0.006332555, 0.006150424, 0.005499009, 0.004766233,
  0.0042406, 0.004177085, 0.004011566, 0.003834336, 0.003683899, 0.003813446, 
    0.004272072, 0.004728941, 0.005424833, 0.006325221, 0.00707855, 
    0.007858709, 0.008783529, 0.009825701, 0.01032892, 0.01078697, 
    0.01125451, 0.01106451, 0.01024131, 0.009515763, 0.008422479, 
    0.007120229, 0.005758964, 0.005014338, 0.004126241, 0.003253962, 
    0.002937105, 0.002859148, 0.002815537, 0.003029098, 0.003518167, 
    0.003930441, 0.004005434, 0.003800439, 0.003535258, 0.003171673, 
    0.002532451, 0.001876766, 0.001624405, 0.002008818, 0.002415702, 
    0.002903256, 0.004226491, 0.005515813, 0.006364668, 0.007167411, 
    0.008018356, 0.008525244, 0.008604435, 0.008623928, 0.008807389, 
    0.008480955, 0.008220238, 0.007420489, 0.006586552,
  0.007229995, 0.007126607, 0.006919661, 0.00672913, 0.00656784, 0.006776634, 
    0.007408408, 0.008039603, 0.00894756, 0.01007753, 0.01102213, 0.01197407, 
    0.01308409, 0.01433724, 0.01489548, 0.01538767, 0.01589213, 0.01553452, 
    0.0143447, 0.01327028, 0.01171428, 0.009918099, 0.00804986, 0.007011004, 
    0.005862986, 0.004732791, 0.004353742, 0.00431585, 0.004325455, 
    0.004628693, 0.005145509, 0.005559602, 0.005563377, 0.005149862, 
    0.00465798, 0.004106394, 0.003280204, 0.002443964, 0.002230242, 
    0.002941315, 0.003670127, 0.004461438, 0.00628954, 0.008072523, 
    0.009183863, 0.01006563, 0.01100733, 0.01148186, 0.01138352, 0.01121188, 
    0.01138065, 0.01092888, 0.0105507, 0.009569168, 0.008633406,
  0.009973269, 0.00977722, 0.009519014, 0.009358403, 0.009220025, 
    0.009557841, 0.01044362, 0.01133092, 0.01253544, 0.01399397, 0.01525828, 
    0.01650699, 0.01789993, 0.01943734, 0.02006149, 0.02058365, 0.02111877, 
    0.02054507, 0.01889357, 0.01735378, 0.0151944, 0.012787, 0.01030495, 
    0.008959375, 0.007556121, 0.006168297, 0.005760864, 0.005812223, 
    0.005924282, 0.006314286, 0.006921509, 0.00741327, 0.007234548, 
    0.00648649, 0.005667619, 0.004858931, 0.003792727, 0.00272991, 
    0.002597561, 0.003754888, 0.004915166, 0.006109907, 0.008605597, 
    0.01105032, 0.01250121, 0.01347292, 0.014507, 0.01489584, 0.01452516, 
    0.01407653, 0.0142168, 0.01360999, 0.01308356, 0.01189753, 0.01086282,
  0.01205063, 0.01172218, 0.01140368, 0.01130874, 0.01122512, 0.01174365, 
    0.01295933, 0.0141787, 0.01575889, 0.01763711, 0.01934293, 0.02100635, 
    0.02276577, 0.02464188, 0.02532443, 0.02587039, 0.02642664, 0.02558718, 
    0.02338249, 0.02127434, 0.01839772, 0.01529925, 0.01212672, 0.01052578, 
    0.008919428, 0.007322521, 0.006971515, 0.007203452, 0.007508769, 
    0.008003585, 0.008702289, 0.009296217, 0.008903379, 0.00769264, 
    0.006406181, 0.00525111, 0.003858199, 0.002471273, 0.002420077, 
    0.004117155, 0.00581567, 0.007517316, 0.01084442, 0.0141318, 0.01601945, 
    0.0171516, 0.01833003, 0.01859984, 0.01788158, 0.0171001, 0.01723147, 
    0.0164644, 0.01576878, 0.0143615, 0.01322623,
  0.01345591, 0.01294224, 0.01248266, 0.01240688, 0.01234011, 0.0130236, 
    0.01457256, 0.01612431, 0.01810879, 0.02043766, 0.02265884, 0.02485322, 
    0.02709551, 0.0293996, 0.03016086, 0.03080569, 0.03145534, 0.03034578, 
    0.02750138, 0.02472473, 0.02099284, 0.01710915, 0.01316612, 0.01142688, 
    0.009716362, 0.008012655, 0.007856665, 0.008397037, 0.009010128, 
    0.009622645, 0.01038011, 0.01104476, 0.0103972, 0.008567251, 0.00660155, 
    0.005067086, 0.003459182, 0.001894827, 0.002048908, 0.004358276, 
    0.006640008, 0.008831471, 0.01285132, 0.01685303, 0.01907484, 0.02029971, 
    0.0215434, 0.02165803, 0.02061289, 0.01954831, 0.01967437, 0.01875855, 
    0.01784445, 0.01619051, 0.01493266,
  0.01391646, 0.0132233, 0.01260038, 0.01254972, 0.01249417, 0.01325725, 
    0.01501822, 0.0167814, 0.01900474, 0.02159309, 0.02417855, 0.02680224, 
    0.02948579, 0.03218198, 0.03304147, 0.03386221, 0.03468334, 0.03342063, 
    0.03007271, 0.02669885, 0.0221214, 0.0175191, 0.01291672, 0.01115, 
    0.009423192, 0.007671441, 0.007603738, 0.008268602, 0.008902404, 
    0.009013633, 0.009045871, 0.009163631, 0.008190008, 0.006231445, 
    0.004204394, 0.002733631, 0.001400375, 8.16645e-05, 0.0006503663, 
    0.003557468, 0.00645091, 0.009104371, 0.01340764, 0.01771816, 0.02006816, 
    0.02124547, 0.02241275, 0.02239352, 0.0212124, 0.02004406, 0.01998114, 
    0.01887535, 0.01772195, 0.01577492, 0.01435783,
  0.01324217, 0.01253056, 0.01186536, 0.01190323, 0.0119322, 0.01281801, 
    0.01481697, 0.01681903, 0.01918786, 0.02182096, 0.02443787, 0.02698769, 
    0.02949308, 0.03201253, 0.03274358, 0.03341462, 0.0340893, 0.03263874, 
    0.02905965, 0.02546728, 0.02074809, 0.01609458, 0.0114472, 0.009992127, 
    0.008486266, 0.006995468, 0.007230654, 0.008095498, 0.00898851, 
    0.00931275, 0.009473083, 0.009728922, 0.008908855, 0.006990836, 
    0.004982901, 0.003579447, 0.002369519, 0.001044169, 0.001422409, 
    0.004135411, 0.006968383, 0.009600878, 0.01371285, 0.01780634, 
    0.02019113, 0.0213176, 0.02250485, 0.02273344, 0.02190413, 0.02099258, 
    0.02071456, 0.01950276, 0.01844066, 0.01639404, 0.01500691,
  0.01220439, 0.01161129, 0.01110567, 0.01135847, 0.01160115, 0.01273892, 
    0.01520889, 0.01768293, 0.02039899, 0.0233813, 0.02628017, 0.02891181, 
    0.0313586, 0.03385947, 0.03455448, 0.03503923, 0.0355294, 0.0339636, 
    0.03034941, 0.02678692, 0.02254777, 0.01856535, 0.01460401, 0.01404969, 
    0.01326833, 0.01259123, 0.01344175, 0.01453585, 0.01575885, 0.01669, 
    0.0175093, 0.01794601, 0.01689999, 0.01503383, 0.01336678, 0.01209221, 
    0.0103154, 0.008368464, 0.008282518, 0.01034402, 0.01258019, 0.01475742, 
    0.01861663, 0.02246069, 0.02495366, 0.0264365, 0.02798743, 0.02853613, 
    0.02797164, 0.02731897, 0.02696744, 0.02584479, 0.02490449, 0.02289038, 
    0.02157488,
  0.009916167, 0.00967037, 0.009550197, 0.01028154, 0.01099718, 0.01280946, 
    0.0161443, 0.01948401, 0.02297753, 0.02666576, 0.03026134, 0.0333347, 
    0.03597517, 0.03867721, 0.03957919, 0.04008781, 0.04060065, 0.03951, 
    0.03681967, 0.03421682, 0.03104926, 0.02833304, 0.02561843, 0.02629349, 
    0.02626343, 0.02634804, 0.02770955, 0.02899104, 0.03045368, 0.03157023, 
    0.0326299, 0.03321163, 0.03210004, 0.0302047, 0.02849692, 0.02710788, 
    0.02441344, 0.02155017, 0.02069015, 0.02137288, 0.02222811, 0.02334817, 
    0.0265144, 0.02963901, 0.03177918, 0.03365539, 0.03556878, 0.03635602, 
    0.03593184, 0.03540234, 0.03514111, 0.03450263, 0.03406414, 0.03224974, 
    0.03098602,
  0.00380238, 0.004210137, 0.004880434, 0.006493942, 0.008094986, 0.01125195, 
    0.01620719, 0.02116502, 0.02649345, 0.03172525, 0.0368993, 0.04172726, 
    0.04623675, 0.05076254, 0.05332414, 0.0559882, 0.05864365, 0.05928016, 
    0.05792007, 0.05664122, 0.05406717, 0.05193437, 0.04978117, 0.0514449, 
    0.05132802, 0.05127217, 0.0526129, 0.05383951, 0.05516314, 0.0557094, 
    0.05688639, 0.05751052, 0.05618534, 0.05381096, 0.05143647, 0.04930354, 
    0.04460103, 0.03989835, 0.03784312, 0.03742092, 0.03699894, 0.03752737, 
    0.04088951, 0.0442516, 0.0462772, 0.04798315, 0.04968924, 0.05019393, 
    0.04949702, 0.04879995, 0.04869959, 0.04856013, 0.04842094, 0.04638703, 
    0.04497231 ;

 u_east =
  0.001466074, -2.602085e-18, 8.673617e-19, -1.734723e-18, 3.469447e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 8.673617e-19, 0, 0, 
    2.602085e-18, 0, 0, 1.734723e-18, -8.673617e-19, -8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.001642626, -2.602085e-18, 8.673617e-19, -1.734723e-18, 3.469447e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 8.673617e-19, 0, 0, 
    2.602085e-18, 0, 0, 1.734723e-18, -8.673617e-19, -8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.001936389, -2.602085e-18, 8.673617e-19, -1.734723e-18, 3.469447e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 8.673617e-19, 0, 0, 
    2.602085e-18, 0, 0, 1.734723e-18, -8.673617e-19, -8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.00219953, -2.602085e-18, 8.673617e-19, -1.734723e-18, 3.469447e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 8.673617e-19, 0, 0, 
    2.602085e-18, 0, 0, 1.734723e-18, -8.673617e-19, -8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.002428095, -2.602085e-18, 8.673617e-19, -1.734723e-18, 3.469447e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 8.673617e-19, 0, 0, 
    2.602085e-18, 0, 0, 1.734723e-18, -8.673617e-19, -8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.002629247, -2.602085e-18, 8.673617e-19, -1.734723e-18, 3.469447e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 8.673617e-19, 0, 0, 
    2.602085e-18, 0, 0, 1.734723e-18, -8.673617e-19, -8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.003040971, -2.602085e-18, 8.673617e-19, -1.734723e-18, 3.469447e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 8.673617e-19, 0, 0, 
    2.602085e-18, 0, 0, 1.734723e-18, -8.673617e-19, -8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.003508306, -2.602085e-18, 8.673617e-19, -1.734723e-18, 3.469447e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 8.673617e-19, 0, 0, 
    2.602085e-18, 0, 0, 1.734723e-18, -8.673617e-19, -8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.003951326, -2.602085e-18, 8.673617e-19, -1.734723e-18, 3.469447e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 8.673617e-19, 0, 0, 
    2.602085e-18, 0, 0, 1.734723e-18, -8.673617e-19, -8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.004385646, -2.602085e-18, 8.673617e-19, -1.734723e-18, 3.469447e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 8.673617e-19, 0, 0, 
    2.602085e-18, 0, 0, 1.734723e-18, -8.673617e-19, -8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.004857041, -2.602085e-18, 8.673617e-19, -1.734723e-18, 3.469447e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 8.673617e-19, 0, 0, 
    2.602085e-18, 0, 0, 1.734723e-18, -8.673617e-19, -8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.005512151, -2.602085e-18, 8.673617e-19, -1.734723e-18, 3.469447e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 8.673617e-19, 0, 0, 
    2.602085e-18, 0, 0, 1.734723e-18, -8.673617e-19, -8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.006197008, -2.602085e-18, 8.673617e-19, -1.734723e-18, 3.469447e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 8.673617e-19, 0, 0, 
    2.602085e-18, 0, 0, 1.734723e-18, -8.673617e-19, -8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.006998337, -2.602085e-18, 8.673617e-19, -1.734723e-18, 3.469447e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 8.673617e-19, 0, 0, 
    2.602085e-18, 0, 0, 1.734723e-18, -8.673617e-19, -8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.008224713, -2.602085e-18, 8.673617e-19, -1.734723e-18, 3.469447e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 8.673617e-19, 0, 0, 
    2.602085e-18, 0, 0, 1.734723e-18, -8.673617e-19, -8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.009505251, -2.602085e-18, 8.673617e-19, -1.734723e-18, 3.469447e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 8.673617e-19, 0, 0, 
    2.602085e-18, 0, 0, 1.734723e-18, -8.673617e-19, -8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.01099717, -2.602085e-18, 8.673617e-19, -1.734723e-18, 3.469447e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 8.673617e-19, 0, 0, 
    2.602085e-18, 0, 0, 1.734723e-18, -8.673617e-19, -8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.01161294, -2.602085e-18, 8.673617e-19, -1.734723e-18, 3.469447e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 8.673617e-19, 0, 0, 
    2.602085e-18, 0, 0, 1.734723e-18, -8.673617e-19, -8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.0116982, -2.602085e-18, 8.673617e-19, -1.734723e-18, 3.469447e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 8.673617e-19, 0, 0, 
    2.602085e-18, 0, 0, 1.734723e-18, -8.673617e-19, -8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.01002061, -2.602085e-18, 8.673617e-19, -1.734723e-18, 3.469447e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 8.673617e-19, 0, 0, 
    2.602085e-18, 0, 0, 1.734723e-18, -8.673617e-19, -8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.008479221, -2.602085e-18, 8.673617e-19, -1.734723e-18, 3.469447e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 8.673617e-19, 0, 0, 
    2.602085e-18, 0, 0, 1.734723e-18, -8.673617e-19, -8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.007479208, -2.602085e-18, 8.673617e-19, -1.734723e-18, 3.469447e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 8.673617e-19, 0, 0, 
    2.602085e-18, 0, 0, 1.734723e-18, -8.673617e-19, -8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.006713503, -2.602085e-18, 8.673617e-19, -1.734723e-18, 3.469447e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 8.673617e-19, 0, 0, 
    2.602085e-18, 0, 0, 1.734723e-18, -8.673617e-19, -8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.006404259, -2.602085e-18, 8.673617e-19, -1.734723e-18, 3.469447e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 8.673617e-19, 0, 0, 
    2.602085e-18, 0, 0, 1.734723e-18, -8.673617e-19, -8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.006360231, -2.602085e-18, 8.673617e-19, -1.734723e-18, 3.469447e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 8.673617e-19, 0, 0, 
    2.602085e-18, 0, 0, 1.734723e-18, -8.673617e-19, -8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.0063251, -2.602085e-18, 8.673617e-19, -1.734723e-18, 3.469447e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 8.673617e-19, 0, 0, 
    2.602085e-18, 0, 0, 1.734723e-18, -8.673617e-19, -8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.006296711, -2.602085e-18, 8.673617e-19, -1.734723e-18, 3.469447e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 8.673617e-19, 0, 0, 
    2.602085e-18, 0, 0, 1.734723e-18, -8.673617e-19, -8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.006296711, -2.602085e-18, 8.673617e-19, -1.734723e-18, 3.469447e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 8.673617e-19, 0, 0, 
    2.602085e-18, 0, 0, 1.734723e-18, -8.673617e-19, -8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.006296711, -2.602085e-18, 8.673617e-19, -1.734723e-18, 3.469447e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 8.673617e-19, 0, 0, 
    2.602085e-18, 0, 0, 1.734723e-18, -8.673617e-19, -8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.006296711, -2.602085e-18, 8.673617e-19, -1.734723e-18, 3.469447e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 8.673617e-19, 0, 0, 
    2.602085e-18, 0, 0, 1.734723e-18, -8.673617e-19, -8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.000486705, 8.673617e-19, 1.734723e-18, -8.673617e-19, 2.602085e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 0, 0, 0, 0, -8.673617e-19, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.0006085275, 8.673617e-19, 1.734723e-18, -8.673617e-19, 2.602085e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 0, 0, 0, 0, -8.673617e-19, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.0008568077, 8.673617e-19, 1.734723e-18, -8.673617e-19, 2.602085e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 0, 0, 0, 0, -8.673617e-19, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.001080886, 8.673617e-19, 1.734723e-18, -8.673617e-19, 2.602085e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 0, 0, 0, 0, -8.673617e-19, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.00127552, 8.673617e-19, 1.734723e-18, -8.673617e-19, 2.602085e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 0, 0, 0, 0, -8.673617e-19, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.001446811, 8.673617e-19, 1.734723e-18, -8.673617e-19, 2.602085e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 0, 0, 0, 0, -8.673617e-19, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.001860361, 8.673617e-19, 1.734723e-18, -8.673617e-19, 2.602085e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 0, 0, 0, 0, -8.673617e-19, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.002340313, 8.673617e-19, 1.734723e-18, -8.673617e-19, 2.602085e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 0, 0, 0, 0, -8.673617e-19, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.002795293, 8.673617e-19, 1.734723e-18, -8.673617e-19, 2.602085e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 0, 0, 0, 0, -8.673617e-19, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.003241339, 8.673617e-19, 1.734723e-18, -8.673617e-19, 2.602085e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 0, 0, 0, 0, -8.673617e-19, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.00371393, 8.673617e-19, 1.734723e-18, -8.673617e-19, 2.602085e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 0, 0, 0, 0, -8.673617e-19, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.004314506, 8.673617e-19, 1.734723e-18, -8.673617e-19, 2.602085e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 0, 0, 0, 0, -8.673617e-19, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.004942353, 8.673617e-19, 1.734723e-18, -8.673617e-19, 2.602085e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 0, 0, 0, 0, -8.673617e-19, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.005689062, 8.673617e-19, 1.734723e-18, -8.673617e-19, 2.602085e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 0, 0, 0, 0, -8.673617e-19, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.006880624, 8.673617e-19, 1.734723e-18, -8.673617e-19, 2.602085e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 0, 0, 0, 0, -8.673617e-19, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.008087293, 8.673617e-19, 1.734723e-18, -8.673617e-19, 2.602085e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 0, 0, 0, 0, -8.673617e-19, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.00935362, 8.673617e-19, 1.734723e-18, -8.673617e-19, 2.602085e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 0, 0, 0, 0, -8.673617e-19, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.009337617, 8.673617e-19, 1.734723e-18, -8.673617e-19, 2.602085e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 0, 0, 0, 0, -8.673617e-19, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.008609463, 8.673617e-19, 1.734723e-18, -8.673617e-19, 2.602085e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 0, 0, 0, 0, -8.673617e-19, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.007013762, 8.673617e-19, 1.734723e-18, -8.673617e-19, 2.602085e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 0, 0, 0, 0, -8.673617e-19, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.005610432, 8.673617e-19, 1.734723e-18, -8.673617e-19, 2.602085e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 0, 0, 0, 0, -8.673617e-19, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.004935597, 8.673617e-19, 1.734723e-18, -8.673617e-19, 2.602085e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 0, 0, 0, 0, -8.673617e-19, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.004455573, 8.673617e-19, 1.734723e-18, -8.673617e-19, 2.602085e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 0, 0, 0, 0, -8.673617e-19, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.00454212, 8.673617e-19, 1.734723e-18, -8.673617e-19, 2.602085e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 0, 0, 0, 0, -8.673617e-19, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.004925412, 8.673617e-19, 1.734723e-18, -8.673617e-19, 2.602085e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 0, 0, 0, 0, -8.673617e-19, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.005231262, 8.673617e-19, 1.734723e-18, -8.673617e-19, 2.602085e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 0, 0, 0, 0, -8.673617e-19, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.005477995, 8.673617e-19, 1.734723e-18, -8.673617e-19, 2.602085e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 0, 0, 0, 0, -8.673617e-19, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.005477995, 8.673617e-19, 1.734723e-18, -8.673617e-19, 2.602085e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 0, 0, 0, 0, -8.673617e-19, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.005477995, 8.673617e-19, 1.734723e-18, -8.673617e-19, 2.602085e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 0, 0, 0, 0, -8.673617e-19, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.005477995, 8.673617e-19, 1.734723e-18, -8.673617e-19, 2.602085e-18, 
    -8.673617e-19, -1.734723e-18, 2.602085e-18, 0, 0, 0, 0, -8.673617e-19, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18 ;

 u_south =
  -0.0005609904, -0.0004633578, 1.162663e-05, 0.0005948897, 0.001179608, 
    0.001657261, 0.001836214, 0.002005413, 0.002272355, 0.002689276, 
    0.003101133, 0.002987586, 0.002993569, 0.00317264, 0.003139157, 
    0.003041232, 0.002928466, 0.0029508, 0.002911107, 0.00279286, 
    0.002690305, 0.002589567, 0.002495976, 0.002277859, 0.00211237, 
    0.002032376, 0.001713253, 0.001479352, 0.001329385, 0.001299939, 
    0.001258944, 0.001218875, 0.001127945, 0.001036676, 0.0009479147, 
    0.0008874572, 0.0008641996, 0.000875823, 0.0009494195, 0.0009785173, 
    0.0009441052, 0.0007935585, 0.0007650956, 0.0008775667, 0.0006746348, 
    -7.825776e-05, 0.000163365, -0.0005870005, -0.0002031225, 0.0001744701, 
    0.0003674711, 0.00101575, 0.001964191, 0.002932148, 0.001466074,
  -0.002268772, -0.002443053, -0.002096892, -0.001697105, -0.001384857, 
    -0.000980037, -0.0007235377, -0.0003525313, 0.0003151879, 0.001256253, 
    0.002377359, 0.002541743, 0.002839819, 0.003282851, 0.003223781, 
    0.003199628, 0.003196689, 0.003100005, 0.002975176, 0.002830121, 
    0.002727602, 0.002625069, 0.002517379, 0.002220651, 0.002025961, 
    0.001945773, 0.001629549, 0.001398384, 0.001247963, 0.001231376, 
    0.001206051, 0.001170577, 0.001084143, 0.00099747, 0.0009139245, 
    0.0008536613, 0.0008299606, 0.0008411143, 0.0009226274, 0.0009302553, 
    0.0008650015, 0.0007072914, 0.0006101782, 0.0004767018, -1.491226e-05, 
    -5.13328e-05, -4.163486e-06, -0.0004005873, -1.78054e-05, 0.0003015892, 
    0.0005955662, 0.001289678, 0.002427111, 0.003285252, 0.001642626,
  -0.002328006, -0.002484559, -0.002137073, -0.001914675, -0.00182397, 
    -0.00144061, -0.0009623311, -0.0003925743, 0.0002732899, 0.00113673, 
    0.002198387, 0.002386991, 0.002692005, 0.003117773, 0.003069481, 
    0.003053809, 0.003058221, 0.00296597, 0.002849339, 0.002711845, 
    0.002605155, 0.002502822, 0.002400564, 0.002116057, 0.001931145, 
    0.001856146, 0.00155931, 0.001340749, 0.001196383, 0.001180067, 
    0.001154796, 0.001118985, 0.00103162, 0.0009492885, 0.0008771659, 
    0.0008250083, 0.0008030116, 0.0008096132, 0.0008860969, 0.0008937848, 
    0.000833595, 0.000682816, 0.000510936, 0.000313219, 1.874009e-06, 
    -2.832456e-05, -0.0001899812, -0.0002412741, 0.0001405885, 0.0004102571, 
    0.0007905944, 0.001523961, 0.002835459, 0.003872778, 0.001936389,
  -0.002347663, -0.002486032, -0.002141843, -0.001914262, -0.00180517, 
    -0.001422703, -0.0009487876, -0.0003940882, 0.0002580782, 0.001082147, 
    0.002082382, 0.002274879, 0.002575345, 0.002985617, 0.002948761, 
    0.002941546, 0.002954033, 0.002867944, 0.002755223, 0.002621762, 
    0.002511214, 0.002407529, 0.002306769, 0.00203061, 0.001851328, 
    0.001778416, 0.001496657, 0.001287032, 0.001145786, 0.001128332, 
    0.001103476, 0.00106976, 0.000985016, 0.0009147748, 0.0008549241, 
    0.0008092581, 0.0007872768, 0.000789549, 0.0008627375, 0.0008715946, 
    0.0008162474, 0.000673835, 0.0005050034, 0.0003088998, 1.629891e-05, 
    -2.907024e-05, -0.0002232389, -8.256143e-05, 0.0002774135, 0.0005460483, 
    0.0009583008, 0.001725488, 0.003186862, 0.00439906, 0.00219953,
  -0.002334728, -0.002454463, -0.002112257, -0.001874168, -0.001741938, 
    -0.001362302, -0.0009009902, -0.0003678681, 0.0002681995, 0.001054897, 
    0.00199617, 0.002191636, 0.002484887, 0.002877625, 0.002850712, 
    0.002850381, 0.002867437, 0.002783981, 0.00267742, 0.002547723, 
    0.002432612, 0.002326469, 0.002226746, 0.001960429, 0.001791116, 
    0.001723526, 0.001456609, 0.001255025, 0.001116693, 0.001098904, 
    0.001076623, 0.001049762, 0.0009723502, 0.000906456, 0.000853758, 
    0.0008136799, 0.0007916421, 0.0007881706, 0.000855637, 0.0008612784, 
    0.000805212, 0.0006662834, 0.0004998609, 0.0003297987, 9.098804e-05, 
    -2.980596e-05, -6.169462e-05, 0.0001011471, 0.0003969629, 0.0007516395, 
    0.001208193, 0.002013253, 0.003491938, 0.004856189, 0.002428095,
  -0.002290677, -0.002392535, -0.002056978, -0.001818619, -0.001673999, 
    -0.001297845, -0.0008418993, -0.0003232881, 0.000296631, 0.001045156, 
    0.001929799, 0.002127903, 0.002416011, 0.002793361, 0.002777183, 
    0.002783835, 0.002806571, 0.002729278, 0.002625742, 0.002499281, 
    0.002382215, 0.002275253, 0.002176029, 0.001917764, 0.001752963, 
    0.00168601, 0.001431664, 0.001237627, 0.001101968, 0.001083437, 
    0.001061943, 0.001037405, 0.0009612276, 0.0008991507, 0.0008527339, 
    0.0008175631, 0.0007954756, 0.0007869601, 0.0008494016, 0.0008612309, 
    0.0008294277, 0.0007253581, 0.0005849897, 0.0004017482, 0.0001656695, 
    1.502854e-05, 8.018337e-05, 0.0002625053, 0.0005019825, 0.0009322794, 
    0.001429847, 0.002359041, 0.004138018, 0.005258494, 0.002629247,
  -0.002218324, -0.002302608, -0.0019719, -0.001726926, -0.001564461, 
    -0.001193949, -0.0007523349, -0.0002555699, 0.0003455387, 0.001057386, 
    0.001886969, 0.002086273, 0.002365905, 0.002725157, 0.002718232, 
    0.002730385, 0.002755333, 0.002680332, 0.002579504, 0.002455937, 
    0.002337122, 0.002229428, 0.00213065, 0.00187959, 0.001718826, 
    0.001652443, 0.001412303, 0.001224545, 0.001091429, 0.001074236, 
    0.001060148, 0.001053799, 0.001002927, 0.0009675453, 0.0009392067, 
    0.0009112222, 0.0008873104, 0.0008766842, 0.0009437537, 0.0009580194, 
    0.0009215424, 0.0008126894, 0.0006629257, 0.0004661281, 0.0002324946, 
    0.0001803672, 0.0002125274, 0.0004069114, 0.0005959817, 0.001093994, 
    0.001628331, 0.00266879, 0.004736474, 0.006081942, 0.003040971,
  -0.00215193, -0.002220085, -0.001893829, -0.001642783, -0.001463943, 
    -0.001098608, -0.0006701456, -0.0001934277, 0.0003904192, 0.00106861, 
    0.001847666, 0.00204807, 0.002319925, 0.002662569, 0.002665484, 
    0.002685205, 0.002720322, 0.002661326, 0.002573719, 0.002454672, 
    0.002331721, 0.002220187, 0.002121374, 0.001886154, 0.001745705, 
    0.00169246, 0.001464855, 0.001285253, 0.001156449, 0.001140799, 
    0.001130404, 0.001129586, 0.001081178, 0.001050138, 0.00102859, 
    0.001008887, 0.0009878413, 0.0009740422, 0.001036804, 0.001046841, 
    0.001006075, 0.0008928324, 0.000734447, 0.0005609992, 0.0003985725, 
    0.0003321027, 0.0003852868, 0.0005305612, 0.000702819, 0.001242462, 
    0.001810596, 0.002953313, 0.005286407, 0.007016613, 0.003508306,
  -0.002030284, -0.002079136, -0.001762238, -0.001515437, -0.001330241, 
    -0.0009713275, -0.0005487985, -8.468976e-05, 0.0004807513, 0.001121388, 
    0.001847872, 0.002050792, 0.00232004, 0.002651293, 0.002666883, 
    0.002692818, 0.002729258, 0.002674852, 0.00259158, 0.002476805, 
    0.0023554, 0.002245152, 0.002147276, 0.001920642, 0.001784247, 
    0.001731044, 0.001514611, 0.001342733, 0.001218011, 0.001203823, 
    0.001196924, 0.001201342, 0.001155268, 0.001128339, 0.001113221, 
    0.001101359, 0.001083026, 0.001066223, 0.001124906, 0.001135078, 
    0.001121554, 0.001046974, 0.0009188656, 0.0007263228, 0.0005614426, 
    0.0004757743, 0.0005488695, 0.0006373483, 0.0009089472, 0.001479606, 
    0.00204583, 0.003222882, 0.005807576, 0.007902651, 0.003951326,
  -0.001902002, -0.001931281, -0.001620403, -0.001369106, -0.001169511, 
    -0.0008174929, -0.0004094436, 3.419229e-05, 0.0005797353, 0.001185832, 
    0.001862364, 0.002066995, 0.002328141, 0.002641792, 0.002668254, 
    0.002700279, 0.002738015, 0.002688106, 0.002609081, 0.002498494, 
    0.002378603, 0.002269615, 0.002172657, 0.001954437, 0.001822015, 
    0.001768852, 0.001566473, 0.001401703, 0.001281123, 0.001270304, 
    0.00127338, 0.001299, 0.001278715, 0.001278334, 0.001281575, 0.00128344, 
    0.001270347, 0.001258909, 0.001326299, 0.001348807, 0.001331919, 
    0.001248167, 0.001103676, 0.0008883259, 0.0007210418, 0.0006620043, 
    0.0007091695, 0.0007419945, 0.001110949, 0.001732452, 0.002417312, 
    0.00381728, 0.006502984, 0.008771292, 0.004385646,
  -0.001771514, -0.001780723, -0.001476879, -0.001221032, -0.001006867, 
    -0.0006618267, -0.0002684296, 0.0001544897, 0.0006798978, 0.001251043, 
    0.001877029, 0.00208339, 0.002337161, 0.002638, 0.002678463, 0.00271919, 
    0.002765417, 0.002733435, 0.002669533, 0.002565887, 0.002446355, 
    0.002336424, 0.002240343, 0.00203974, 0.001927331, 0.001886499, 
    0.001696513, 0.00154106, 0.001426577, 0.001420459, 0.001431797, 
    0.00146856, 0.001451676, 0.001456417, 0.001467788, 0.001486263, 
    0.001484856, 0.001478872, 0.001544792, 0.001565079, 0.001544787, 
    0.001451754, 0.001290685, 0.001054173, 0.0009171017, 0.000864178, 
    0.0008611705, 0.0008478835, 0.001315346, 0.001988289, 0.002793178, 
    0.004502844, 0.007685104, 0.009714082, 0.004857041,
  -0.001616665, -0.001597243, -0.00129853, -0.001040659, -0.0008149596, 
    -0.0004767347, -9.416488e-05, 0.0003132249, 0.0008188137, 0.001355204, 
    0.001932456, 0.002144016, 0.002394539, 0.002678554, 0.002734909, 
    0.002784861, 0.002833182, 0.0028108, 0.002755126, 0.002659031, 
    0.002545812, 0.0024403, 0.00234637, 0.002157266, 0.002049794, 
    0.002008811, 0.001831243, 0.001685443, 0.001577277, 0.001576029, 
    0.001595927, 0.001644234, 0.001630872, 0.001640922, 0.001660714, 
    0.001696399, 0.0017071, 0.001706766, 0.001771163, 0.001789314, 
    0.001767279, 0.001670903, 0.001510629, 0.00128482, 0.001148136, 
    0.001073637, 0.0009820892, 0.001022407, 0.001530921, 0.002253298, 
    0.003182481, 0.00521282, 0.008909103, 0.0110243, 0.005512151,
  -0.001454623, -0.00140524, -0.001111729, -0.0008485165, -0.0006078162, 
    -0.0002764602, 9.198351e-05, 0.0004799759, 0.0009642898, 0.001465988, 
    0.001994106, 0.002210649, 0.002454582, 0.002720992, 0.002793977, 
    0.002853582, 0.002904095, 0.002891757, 0.002844414, 0.002756335, 
    0.002649988, 0.002549001, 0.002457321, 0.002280572, 0.002178973, 
    0.002137343, 0.001972338, 0.00183596, 0.001733529, 0.001736568, 
    0.001764839, 0.001824827, 0.001811096, 0.001820954, 0.001843418, 
    0.001901494, 0.001931736, 0.001946108, 0.002008932, 0.002027499, 
    0.002007208, 0.001909457, 0.001749602, 0.001526173, 0.001389895, 
    0.00126226, 0.001108616, 0.001306385, 0.001938903, 0.00276581, 
    0.003801713, 0.006010512, 0.01018898, 0.01239402, 0.006197008,
  -0.001365998, -0.001282, -0.000987932, -0.0007094695, -0.0004448007, 
    -0.0001185882, 0.0002312771, 0.0005973931, 0.001063258, 0.001538132, 
    0.002025852, 0.002250914, 0.002490132, 0.002741654, 0.002835872, 
    0.002909268, 0.002964474, 0.002967258, 0.002933086, 0.002855325, 
    0.002761743, 0.00266752, 0.002576213, 0.002414644, 0.002317799, 
    0.00227233, 0.002119345, 0.001991366, 0.001893085, 0.001899211, 
    0.0019361, 0.002009473, 0.001994991, 0.002005582, 0.002031559, 
    0.002113208, 0.002164244, 0.002195223, 0.002256349, 0.002275292, 
    0.002256815, 0.002157633, 0.001982453, 0.001740565, 0.001584381, 
    0.001426293, 0.001280828, 0.001601796, 0.002363288, 0.003405209, 
    0.00487301, 0.007680174, 0.01226911, 0.01399667, 0.006998337,
  -0.001323486, -0.001202206, -0.000909235, -0.000622924, -0.0003417069, 
    -1.900601e-05, 0.0003230011, 0.0006779199, 0.001129134, 0.001579085, 
    0.00203109, 0.002268621, 0.002509424, 0.002751899, 0.002870861, 
    0.002960559, 0.003023268, 0.003043892, 0.003023445, 0.002956199, 
    0.002875625, 0.00278834, 0.00269742, 0.002551268, 0.002455054, 
    0.002397178, 0.002253862, 0.002133981, 0.002038753, 0.002044504, 
    0.002083094, 0.00215554, 0.002117984, 0.002105678, 0.00211894, 
    0.002221532, 0.002296865, 0.002346419, 0.002397146, 0.00240773, 
    0.002382329, 0.002282423, 0.002117713, 0.001881658, 0.001755037, 
    0.001604402, 0.001598808, 0.002058098, 0.002935742, 0.004091869, 
    0.005964538, 0.009381256, 0.01465619, 0.01644943, 0.008224713,
  -0.00137204, -0.001227809, -0.0009337882, -0.0006322073, -0.0003270797, 
    -8.83234e-06, 0.000317888, 0.0006564975, 0.001096754, 0.001533042, 
    0.001962946, 0.00221584, 0.002459827, 0.00269743, 0.002843163, 
    0.002952829, 0.003025164, 0.003059744, 0.003047512, 0.002985158, 
    0.002925956, 0.002844789, 0.002743472, 0.002611481, 0.002511277, 
    0.002436068, 0.002302256, 0.002185573, 0.002087048, 0.002081607, 
    0.002115487, 0.002189546, 0.002141158, 0.002119124, 0.002123715, 
    0.002242456, 0.002337059, 0.002408772, 0.002456492, 0.00247527, 
    0.002468618, 0.002398577, 0.00225204, 0.002038048, 0.001975637, 
    0.001915826, 0.00193826, 0.002620749, 0.003883411, 0.005635579, 
    0.008036318, 0.01197637, 0.01781008, 0.0190105, 0.009505251,
  -0.001467527, -0.001309121, -0.001018084, -0.0007118228, -0.0003936494, 
    -8.121141e-05, 0.0002404865, 0.0005742642, 0.001008234, 0.001433035, 
    0.001846674, 0.002117839, 0.002373829, 0.002616727, 0.002791908, 
    0.002926889, 0.00303097, 0.003108539, 0.003121383, 0.003060016, 
    0.003013915, 0.002928515, 0.002809637, 0.002702269, 0.002611733, 
    0.002519057, 0.002394164, 0.002276974, 0.002171304, 0.002145353, 
    0.002165622, 0.002231645, 0.002164797, 0.002121926, 0.0021048, 
    0.002224901, 0.002330932, 0.00242182, 0.002459953, 0.002484906, 
    0.00250067, 0.002474955, 0.002386835, 0.002238367, 0.002235475, 
    0.002282159, 0.002540766, 0.003533981, 0.005151809, 0.007347585, 
    0.0101895, 0.01491282, 0.02146652, 0.02199434, 0.01099717,
  -0.001152911, -0.00103339, -0.0007629328, -0.0004812057, -0.0001812323, 
    0.0001104057, 0.0004270997, 0.000759305, 0.001180978, 0.001589613, 
    0.001989879, 0.002279605, 0.002558447, 0.002822913, 0.003030453, 
    0.003189405, 0.003308812, 0.003392189, 0.003397578, 0.003317321, 
    0.003290694, 0.003193743, 0.003031171, 0.002935428, 0.002824226, 
    0.002682244, 0.002558701, 0.002435677, 0.002316255, 0.002252229, 
    0.002240775, 0.002281518, 0.002187643, 0.00213805, 0.002118194, 
    0.002226742, 0.002327797, 0.002435919, 0.002476506, 0.002530055, 
    0.002602066, 0.002660483, 0.002663715, 0.002616814, 0.002728894, 
    0.002867915, 0.003388438, 0.004662008, 0.007116578, 0.01017572, 
    0.01389345, 0.01925079, 0.02556915, 0.02322588, 0.01161294,
  -0.0002496155, -0.000184756, 5.284074e-05, 0.0002690607, 0.0005030173, 
    0.0007665514, 0.001104421, 0.001463415, 0.001868568, 0.002244948, 
    0.002623153, 0.00293827, 0.003267864, 0.003586544, 0.003842722, 
    0.004040945, 0.004227984, 0.004390157, 0.004428547, 0.004311674, 
    0.004279039, 0.004133984, 0.003895355, 0.003835519, 0.003747144, 
    0.003569687, 0.003448825, 0.003305828, 0.003159705, 0.00303187, 
    0.002972274, 0.002987415, 0.00289089, 0.002807005, 0.002719808, 
    0.002773694, 0.002834255, 0.002913024, 0.002906502, 0.002932747, 
    0.002996118, 0.003063881, 0.003097561, 0.003155428, 0.003477651, 
    0.003952529, 0.004615336, 0.00694835, 0.01025073, 0.01394989, 0.01828144, 
    0.02384645, 0.02739459, 0.02339641, 0.0116982,
  0.001321838, 0.001322403, 0.00152731, 0.001661284, 0.00184941, 0.002081041, 
    0.002395265, 0.002791442, 0.003172183, 0.003507434, 0.003861035, 
    0.004207878, 0.004605454, 0.004999626, 0.005319322, 0.005569581, 
    0.005853396, 0.006134808, 0.006231084, 0.006069926, 0.006022012, 
    0.005808669, 0.005472917, 0.005469225, 0.005441986, 0.005252949, 
    0.005145276, 0.004980891, 0.004808696, 0.004613554, 0.004512285, 
    0.004529563, 0.004485127, 0.004430096, 0.004305494, 0.004267982, 
    0.004230785, 0.004238373, 0.004186268, 0.004200043, 0.004288823, 
    0.004408537, 0.004510108, 0.004595018, 0.004830789, 0.005606846, 
    0.007077972, 0.01016005, 0.01428911, 0.01863522, 0.0232661, 0.02713679, 
    0.02729297, 0.02004121, 0.01002061,
  0.004142272, 0.004124016, 0.004362497, 0.004498768, 0.004591932, 
    0.004809035, 0.005149115, 0.005530977, 0.005864007, 0.006194165, 
    0.006570472, 0.006980777, 0.007417384, 0.00783872, 0.008226863, 
    0.008534863, 0.008841802, 0.009103904, 0.009154129, 0.008936959, 
    0.008934719, 0.008695263, 0.008251631, 0.00823086, 0.008150209, 
    0.007937326, 0.007849379, 0.007671904, 0.007482848, 0.007222373, 
    0.00708237, 0.007113371, 0.007150874, 0.007153392, 0.007003759, 
    0.006868464, 0.006708881, 0.006617651, 0.006524834, 0.006537095, 
    0.006675545, 0.006872735, 0.007057701, 0.007218823, 0.00761079, 
    0.008295927, 0.0106949, 0.01447465, 0.01957505, 0.02412349, 0.02770485, 
    0.0274502, 0.02419884, 0.01695844, 0.008479221,
  0.00728587, 0.007329006, 0.007629429, 0.007745986, 0.007751046, 
    0.007988757, 0.008382455, 0.008832127, 0.00913059, 0.009451579, 
    0.009857967, 0.01038856, 0.01095251, 0.01149556, 0.01203871, 0.01248323, 
    0.01293931, 0.01334487, 0.01346541, 0.01321885, 0.01328177, 0.01301369, 
    0.0124636, 0.01252184, 0.01246028, 0.01212184, 0.01206272, 0.01192902, 
    0.01177986, 0.01148972, 0.01130123, 0.01125271, 0.01120025, 0.01123908, 
    0.01107484, 0.01087754, 0.01061453, 0.01042135, 0.01030362, 0.01032426, 
    0.01052452, 0.01079898, 0.01105709, 0.01126195, 0.01186853, 0.01299908, 
    0.01560237, 0.02026902, 0.0260642, 0.02922312, 0.02832133, 0.02420738, 
    0.02154736, 0.01495842, 0.007479208,
  0.01020649, 0.01037513, 0.01077426, 0.01092051, 0.01087896, 0.01116546, 
    0.01161374, 0.01213332, 0.01240975, 0.01275423, 0.01322567, 0.01391596, 
    0.01462096, 0.0152885, 0.0160258, 0.01664103, 0.01724787, 0.01778612, 
    0.01797164, 0.01771418, 0.01789046, 0.01763181, 0.01699167, 0.01713047, 
    0.01711128, 0.01676447, 0.0168086, 0.01678783, 0.01676856, 0.01656139, 
    0.01648071, 0.01658079, 0.01668086, 0.01670788, 0.0165409, 0.01643229, 
    0.01622615, 0.01602415, 0.0159048, 0.01587752, 0.016063, 0.01637913, 
    0.01665739, 0.01683451, 0.0176682, 0.01920019, 0.02197757, 0.02740013, 
    0.03227586, 0.02997698, 0.02541068, 0.02106143, 0.0198624, 0.01342701, 
    0.006713503,
  0.01250105, 0.01283195, 0.01335147, 0.01356559, 0.01351962, 0.0138704, 
    0.01437111, 0.01495762, 0.0152346, 0.01563565, 0.01620401, 0.01707906, 
    0.01793205, 0.01872298, 0.01967983, 0.02048282, 0.02122683, 0.02187783, 
    0.02210825, 0.02183809, 0.02214364, 0.0219046, 0.02116689, 0.02135151, 
    0.02132108, 0.02093396, 0.0210807, 0.02121202, 0.02138399, 0.02132919, 
    0.0214382, 0.02176842, 0.0220338, 0.02222626, 0.02222389, 0.02240506, 
    0.02245108, 0.02247252, 0.02257363, 0.0227744, 0.0231216, 0.02348554, 
    0.02377216, 0.0238858, 0.02494276, 0.02666754, 0.02914213, 0.03388106, 
    0.0328516, 0.02765563, 0.02223456, 0.01947177, 0.01853365, 0.01280852, 
    0.006404259,
  0.0139251, 0.01446996, 0.01515033, 0.01547439, 0.01546986, 0.01591671, 
    0.01647353, 0.01708984, 0.01735142, 0.01779559, 0.01845134, 0.01950623, 
    0.02049637, 0.02139639, 0.02258512, 0.02357362, 0.02442648, 0.02517879, 
    0.02543824, 0.02514488, 0.02557009, 0.02532996, 0.02445737, 0.02464057, 
    0.02453969, 0.02405805, 0.02426852, 0.0245433, 0.0249189, 0.02503918, 
    0.02538334, 0.02599838, 0.02641552, 0.02677841, 0.02699355, 0.02762904, 
    0.02813929, 0.02861769, 0.02906256, 0.02962598, 0.03035482, 0.03089929, 
    0.03123098, 0.03130468, 0.03239815, 0.03372826, 0.03397351, 0.03429864, 
    0.03104703, 0.02502943, 0.02079542, 0.01822434, 0.01788121, 0.01272046, 
    0.006360231,
  0.01404635, 0.01493656, 0.01578319, 0.01626174, 0.01637142, 0.01698733, 
    0.01769586, 0.01850071, 0.01890764, 0.01942298, 0.02006968, 0.02118701, 
    0.02216429, 0.02297593, 0.02421312, 0.02518588, 0.02590892, 0.02652868, 
    0.02664917, 0.02627084, 0.026713, 0.0264702, 0.02554333, 0.02571487, 
    0.02559915, 0.0251957, 0.02555518, 0.0260789, 0.02677558, 0.02722423, 
    0.02789824, 0.02882866, 0.0294263, 0.02986073, 0.03021028, 0.03129591, 
    0.03230593, 0.03325197, 0.03383839, 0.03446613, 0.03513316, 0.0355907, 
    0.03572532, 0.03552882, 0.03595291, 0.03557082, 0.03406942, 0.03271885, 
    0.02909391, 0.02380942, 0.01984302, 0.0184158, 0.01744717, 0.0126502, 
    0.0063251,
  0.01379195, 0.01479076, 0.01555596, 0.01597813, 0.01605329, 0.01661227, 
    0.01724857, 0.01797288, 0.01835593, 0.01888016, 0.01952656, 0.0206439, 
    0.02146034, 0.02198528, 0.02305584, 0.02377977, 0.02410828, 0.02437645, 
    0.02420552, 0.02364497, 0.02382652, 0.02350351, 0.02264187, 0.02280985, 
    0.02270105, 0.02241017, 0.02316607, 0.02411543, 0.02522821, 0.02613939, 
    0.02726339, 0.0286106, 0.02947387, 0.03012549, 0.03056051, 0.03176763, 
    0.03282762, 0.03373497, 0.03416819, 0.03466852, 0.03524066, 0.03577631, 
    0.03592939, 0.03569081, 0.03601653, 0.03512777, 0.03261835, 0.03135275, 
    0.02799957, 0.02368888, 0.02087135, 0.01864683, 0.01709867, 0.01259342, 
    0.006296711,
  0.01453415, 0.01545924, 0.01611431, 0.01639954, 0.01632632, 0.01675198, 
    0.01728412, 0.01791287, 0.01822691, 0.01862866, 0.01912301, 0.02024987, 
    0.02103134, 0.02146515, 0.02245723, 0.02303169, 0.0231803, 0.02330003, 
    0.02290096, 0.0220004, 0.02187447, 0.02129626, 0.02025187, 0.02026688, 
    0.02021305, 0.02015004, 0.02104437, 0.02227693, 0.02383055, 0.02511041, 
    0.02654592, 0.02813851, 0.02918708, 0.02990131, 0.03027369, 0.03145394, 
    0.03249533, 0.03339436, 0.03386976, 0.03444541, 0.03519313, 0.03582549, 
    0.03596774, 0.03562515, 0.03584863, 0.03464885, 0.03196511, 0.03050924, 
    0.02857028, 0.02535811, 0.02170031, 0.01883426, 0.01695137, 0.01259342, 
    0.006296711,
  0.0164004, 0.01713146, 0.01768159, 0.0178555, 0.01766733, 0.01798559, 
    0.01846103, 0.01907679, 0.01948098, 0.01993984, 0.02046395, 0.02160259, 
    0.0222415, 0.02236279, 0.02330067, 0.02360971, 0.02329099, 0.02316211, 
    0.02241647, 0.02106266, 0.02039719, 0.01941274, 0.01809734, 0.01784214, 
    0.01778838, 0.01798008, 0.01918623, 0.02092523, 0.0231858, 0.02517864, 
    0.02741817, 0.02992526, 0.03189907, 0.03337025, 0.03428831, 0.03571502, 
    0.03671911, 0.03733315, 0.037824, 0.03820718, 0.0385747, 0.03867368, 
    0.03833074, 0.03748034, 0.03713941, 0.03590681, 0.0338391, 0.03252438, 
    0.02995479, 0.02664274, 0.02207021, 0.01883975, 0.01695137, 0.01259342, 
    0.006296711,
  0.02181502, 0.02211894, 0.02257652, 0.02253128, 0.02200015, 0.0220748, 
    0.022321, 0.02271881, 0.0230113, 0.0234561, 0.02406269, 0.02526185, 
    0.02578332, 0.02561697, 0.026701, 0.02684277, 0.02605265, 0.02566681, 
    0.02454301, 0.0226775, 0.02139609, 0.01997352, 0.01840935, 0.01811234, 
    0.01826023, 0.01884916, 0.02081704, 0.0235764, 0.02712725, 0.03012065, 
    0.03349457, 0.03724903, 0.04028115, 0.04243103, 0.04369867, 0.04567214, 
    0.04698727, 0.04764403, 0.0484382, 0.04871991, 0.04848917, 0.04772552, 
    0.04608527, 0.04356841, 0.0417806, 0.03934333, 0.03625658, 0.03350467, 
    0.03030006, 0.02664274, 0.02207021, 0.01883975, 0.01695137, 0.01259342, 
    0.006296711,
  -0.0008747782, -0.0007911554, -0.0004619039, -6.275935e-05, 0.0003473594, 
    0.0007082514, 0.0008512459, 0.0009699367, 0.00112668, 0.001358047, 
    0.001553163, 0.001489344, 0.001502652, 0.001628678, 0.001583004, 
    0.001506884, 0.001416319, 0.001360187, 0.001281413, 0.001189368, 
    0.001142005, 0.001102707, 0.001062829, 0.0009234047, 0.0008145094, 
    0.0007982749, 0.0006302141, 0.0005476022, 0.0005402043, 0.0005996764, 
    0.000642806, 0.0006847489, 0.0007282568, 0.0007608937, 0.0007844177, 
    0.0007905756, 0.0007927371, 0.0007880151, 0.0009304385, 0.00102355, 
    0.001035924, 0.0008214139, 0.0008473934, 0.001093907, 0.0007403736, 
    -0.0004342074, -0.0001426325, -0.002096713, -0.001929009, -0.001306232, 
    -0.0006309382, -8.834258e-05, 0.0004121025, 0.0009734099, 0.000486705,
  -0.002029441, -0.002074885, -0.00181563, -0.001556724, -0.001380261, 
    -0.001069695, -0.0008794503, -0.0006334311, -0.0002745381, 0.000281125, 
    0.0009668351, 0.001094582, 0.001291199, 0.001568742, 0.001521553, 
    0.001488837, 0.001455097, 0.001320961, 0.001188851, 0.001067096, 
    0.001000904, 0.0009512462, 0.000912519, 0.0007433097, 0.0006616664, 
    0.0006808475, 0.000530262, 0.0004568268, 0.0004560332, 0.0005307366, 
    0.0005925377, 0.0006401176, 0.000689611, 0.000727316, 0.0007558733, 
    0.0007555297, 0.0007510119, 0.0007407928, 0.0009582148, 0.001036725, 
    0.0009746879, 0.0006999883, 0.0005496773, 0.0003552479, -0.0004222489, 
    -0.0005282257, -0.0007010479, -0.00197203, -0.001905731, -0.001159078, 
    -0.0004991502, 1.377273e-05, 0.0006967039, 0.001217055, 0.0006085275,
  -0.002086224, -0.00211168, -0.001851727, -0.001703615, -0.001673558, 
    -0.001378372, -0.001039911, -0.0006608869, -0.0003057625, 0.0001869534, 
    0.0008181509, 0.0009610003, 0.001158052, 0.001411938, 0.001366999, 
    0.001333164, 0.00129625, 0.001169254, 0.001048499, 0.0009372587, 
    0.0008667523, 0.0008179325, 0.0007860629, 0.0006315989, 0.0005621808, 
    0.0005888288, 0.0004587643, 0.0003994376, 0.0004067942, 0.0004844247, 
    0.0005481356, 0.0005966692, 0.0006492394, 0.0006940019, 0.0007342506, 
    0.000735409, 0.0007267643, 0.0007069189, 0.00090356, 0.0009682525, 
    0.0008994992, 0.0006320894, 0.0003330202, 2.171799e-06, -0.0005149915, 
    -0.0006085675, -0.00128781, -0.001865472, -0.001885835, -0.001033283, 
    -0.0003864676, 0.0001011093, 0.0009492578, 0.001713615, 0.0008568077,
  -0.002103638, -0.002109033, -0.001852992, -0.001700699, -0.001653532, 
    -0.001359962, -0.001023561, -0.0006538487, -0.0003100646, 0.0001484727, 
    0.0007263173, 0.0008697795, 0.001058452, 0.001291962, 0.001250485, 
    0.001215914, 0.00117715, 0.001058976, 0.0009445221, 0.0008399312, 
    0.0007646915, 0.0007150126, 0.0006865356, 0.0005420937, 0.0004802534, 
    0.0005111568, 0.0003970817, 0.0003482756, 0.0003610071, 0.0004403117, 
    0.0005059675, 0.0005568171, 0.000614348, 0.0006730349, 0.0007257637, 
    0.0007270747, 0.0007126086, 0.0006829289, 0.0008613289, 0.0009114117, 
    0.0008285392, 0.0005558608, 0.0002503701, -8.973942e-05, -0.0005946877, 
    -0.0008716928, -0.001572693, -0.001809365, -0.001809014, -0.0009128714, 
    -0.0002895709, 0.0001762349, 0.001166592, 0.002161772, 0.001080886,
  -0.00208863, -0.002073823, -0.001820371, -0.001658795, -0.001590371, 
    -0.001300094, -0.0009734196, -0.0006191499, -0.0002885386, 0.0001388122, 
    0.0006671148, 0.0008103097, 0.0009873719, 0.001197958, 0.001158537, 
    0.001122067, 0.001078282, 0.0009645167, 0.0008584298, 0.0007598759, 
    0.0006790336, 0.0006273053, 0.0006015589, 0.0004683181, 0.0004181139, 
    0.0004567668, 0.0003583748, 0.0003191933, 0.0003372131, 0.0004192746, 
    0.0004892662, 0.0005474038, 0.0006151858, 0.0006788759, 0.0007379714, 
    0.0007380956, 0.0007165427, 0.0006738341, 0.0008324726, 0.0008640897, 
    0.0007643955, 0.0004894396, 0.0001787283, -0.0001641468, -0.0006751457, 
    -0.001100627, -0.00148932, -0.001835788, -0.001661888, -0.0007830228, 
    -0.0001819778, 0.0003240316, 0.001355275, 0.00255104, 0.00127552,
  -0.002041423, -0.002007721, -0.001761543, -0.001601174, -0.001522386, 
    -0.001235943, -0.0009117225, -0.0005657235, -0.0002477698, 0.0001476511, 
    0.0006284882, 0.0007712209, 0.0009398501, 0.001131026, 0.001094581, 
    0.001056283, 0.001008732, 0.0009023341, 0.0008006092, 0.0007072297, 
    0.0006223216, 0.0005697842, 0.0005467086, 0.0004221207, 0.0003781079, 
    0.000420076, 0.0003349666, 0.0003048866, 0.0003279701, 0.0004123752, 
    0.0004846209, 0.0005449073, 0.0006159215, 0.0006840054, 0.0007486917, 
    0.0007477736, 0.0007199974, 0.0006658473, 0.0008071319, 0.0008297515, 
    0.0007325038, 0.0004710552, 0.0001564494, -0.0002180442, -0.0007474665, 
    -0.001239111, -0.001416096, -0.001858997, -0.001532644, -0.0006689331, 
    -8.695957e-05, 0.0005218615, 0.001874108, 0.002893623, 0.001446811,
  -0.001964902, -0.001913074, -0.001672215, -0.001506632, -0.001412384, 
    -0.001131653, -0.0008186516, -0.0004882808, -0.000185034, 0.0001811342, 
    0.0006176273, 0.0007578325, 0.0009135848, 0.001081764, 0.001046489, 
    0.001004922, 0.0009501702, 0.0008466959, 0.0007488739, 0.0006601242, 
    0.0005715782, 0.0005183169, 0.000497631, 0.0003807853, 0.0003423122, 
    0.0003872466, 0.0003170115, 0.0002945932, 0.0003223738, 0.0004109796, 
    0.0004922053, 0.0005709918, 0.0006699862, 0.0007656805, 0.0008471232, 
    0.0008454782, 0.0008064482, 0.0007388297, 0.000869796, 0.0008765932, 
    0.0007547429, 0.000475563, 0.0001373145, -0.0002662712, -0.0008121794, 
    -0.001190738, -0.001359434, -0.001879767, -0.001416962, -0.0005667962, 
    -1.874158e-06, 0.0006990731, 0.002357223, 0.003720722, 0.001860361,
  -0.001894681, -0.00182622, -0.001590243, -0.001419874, -0.00131144, 
    -0.00103595, -0.0007332443, -0.0004172147, -0.000127464, 0.0002118602, 
    0.0006076609, 0.0007455466, 0.0008894823, 0.001036559, 0.001003926, 
    0.0009621972, 0.0009099143, 0.0008239473, 0.0007406767, 0.0006576618, 
    0.0005620315, 0.0005045087, 0.0004857923, 0.0003846185, 0.0003677747, 
    0.0004291752, 0.0003715666, 0.0003585364, 0.0003930028, 0.0004869564, 
    0.0005736183, 0.0006575953, 0.000760943, 0.0008610307, 0.0009476474, 
    0.0009467077, 0.0009011108, 0.0008190584, 0.0009328228, 0.0009195791, 
    0.0007751515, 0.0004796997, 0.0001197545, -0.0002783266, -0.0007757718, 
    -0.001146345, -0.001391931, -0.001823762, -0.001300492, -0.0004730257, 
    7.625856e-05, 0.0008618524, 0.002801167, 0.004680627, 0.002340313,
  -0.001768961, -0.001681707, -0.001455469, -0.001290691, -0.0011782, 
    -0.0009088196, -0.0006086849, -0.00029857, -2.16876e-05, 0.0002885048, 
    0.000643142, 0.0007801151, 0.0009184954, 0.001051314, 0.001023399, 
    0.0009791788, 0.000919061, 0.0008368474, 0.0007579279, 0.0006800292, 
    0.0005826175, 0.0005257772, 0.000510159, 0.0004166368, 0.0004050003, 
    0.0004695817, 0.0004232203, 0.000419079, 0.0004598755, 0.0005588926, 
    0.0006507017, 0.0007395932, 0.0008470629, 0.0009513106, 0.001042826, 
    0.001042554, 0.0009907397, 0.0008950208, 0.0009924981, 0.0009640955, 
    0.0008267846, 0.0005485651, 0.0001991301, -0.0002218056, -0.0007361575, 
    -0.001104311, -0.001422702, -0.001683744, -0.001137684, -0.000331451, 
    0.0002001476, 0.001016076, 0.003221891, 0.005590586, 0.002795293,
  -0.001636619, -0.001530443, -0.001310629, -0.001142848, -0.001018591, 
    -0.0007555188, -0.0004661037, -0.0001696196, 9.31813e-05, 0.0003779661, 
    0.0006950655, 0.0008300675, 0.0009564108, 0.00106763, 0.00104248, 
    0.0009958191, 0.0009280238, 0.0008494883, 0.0007748325, 0.0007019471, 
    0.0006027899, 0.0005466182, 0.0005340361, 0.0004480117, 0.0004414779, 
    0.0005091762, 0.0004770628, 0.0004811242, 0.0005282537, 0.0006342923, 
    0.0007380652, 0.0008487672, 0.0009850765, 0.001117093, 0.001225955, 
    0.001230803, 0.001171631, 0.001064739, 0.001157831, 0.001125083, 
    0.0009660034, 0.000657669, 0.0002802828, -0.0001664199, -0.0006973389, 
    -0.001100641, -0.001452855, -0.001546533, -0.0009781349, -0.0001815319, 
    0.0004338781, 0.001472348, 0.003825742, 0.006482678, 0.003241339,
  -0.00150219, -0.001376651, -0.001164063, -0.0009932443, -0.0008570821, 
    -0.0006003928, -0.0003218249, -3.91339e-05, 0.0002094178, 0.0004684925, 
    0.0007476073, 0.0008806146, 0.0009957294, 0.001091056, 0.001072244, 
    0.001026208, 0.0009595214, 0.0008996617, 0.0008407673, 0.000775016, 
    0.0006717104, 0.0006132945, 0.0006036771, 0.000533667, 0.0005486158, 
    0.0006331076, 0.0006121671, 0.0006258393, 0.0006808726, 0.000796706, 
    0.0009115287, 0.001033811, 0.001175401, 0.00131257, 0.001427941, 
    0.001440449, 0.001379375, 0.001259734, 0.001338788, 0.001287987, 
    0.001106879, 0.0007680713, 0.0003624012, -0.0001122608, -0.0006777538, 
    -0.001108264, -0.001439095, -0.001407692, -0.0008166941, -2.983876e-05, 
    0.0006703664, 0.002011733, 0.004932803, 0.007427861, 0.00371393,
  -0.001348134, -0.001196101, -0.0009896056, -0.0008178478, -0.0006721253, 
    -0.0004208501, -0.0001484777, 0.0001272327, 0.0003646303, 0.0006010237, 
    0.0008467246, 0.0009823838, 0.00109208, 0.001168174, 0.001157449, 
    0.001112656, 0.001039786, 0.0009872506, 0.0009353101, 0.0008768349, 
    0.0007751788, 0.0007199469, 0.0007147016, 0.0006531553, 0.0006735901, 
    0.0007619559, 0.0007521432, 0.0007757727, 0.0008389949, 0.0009649762, 
    0.001091247, 0.001225528, 0.001372588, 0.001515095, 0.00163721, 
    0.001657654, 0.001594609, 0.001461759, 0.001526268, 0.001458106, 
    0.001261786, 0.0009046935, 0.0004563815, -0.0001140706, -0.0006733683, 
    -0.001116162, -0.001266205, -0.001221924, -0.000646774, 0.0001272926, 
    0.0009153087, 0.002570325, 0.006079084, 0.008629013, 0.004314506,
  -0.001186923, -0.001007166, -0.0008069158, -0.0006317384, -0.0004738158, 
    -0.0002277622, 3.613223e-05, 0.0003019148, 0.0005271592, 0.0007415992, 
    0.0009544977, 0.001092493, 0.001192906, 0.001248874, 0.00124661, 
    0.001203118, 0.001123778, 0.001078907, 0.001034914, 0.0009842059, 
    0.0008839669, 0.0008315526, 0.0008308825, 0.0007790981, 0.0008072421, 
    0.0009002351, 0.0009010902, 0.000933737, 0.001004087, 0.001140691, 
    0.00127986, 0.001429266, 0.001580281, 0.001725663, 0.001851809, 
    0.001887354, 0.00182896, 0.001689453, 0.001743451, 0.001664976, 
    0.001456536, 0.001072631, 0.0005577221, -0.0001159644, -0.0006687794, 
    -0.0010214, -0.001085296, -0.0009619673, -0.0003413867, 0.0005060448, 
    0.001372295, 0.003210666, 0.007277695, 0.009884707, 0.004942353,
  -0.00110537, -0.0008949084, -0.000696377, -0.0005073059, -0.000326776, 
    -8.398494e-05, 0.0001667976, 0.0004206894, 0.0006385098, 0.0008408241, 
    0.001031269, 0.001177013, 0.001272007, 0.00131296, 0.001326205, 
    0.001290801, 0.001211267, 0.001180976, 0.00114864, 0.001106972, 
    0.00101449, 0.0009670859, 0.0009684312, 0.0009263949, 0.0009586803, 
    0.001052202, 0.001061079, 0.001100295, 0.001175065, 0.001322778, 
    0.001476946, 0.001644337, 0.001797019, 0.001944448, 0.002074623, 
    0.00212659, 0.002074132, 0.001928565, 0.001970736, 0.001880191, 
    0.001659141, 0.001247341, 0.0006678001, -5.976134e-05, -0.0005297969, 
    -0.0008142433, -0.0008651181, -0.0006915446, -2.372097e-05, 0.0009968756, 
    0.002252159, 0.004730303, 0.009250022, 0.01137812, 0.005689062,
  -0.001073775, -0.0008309688, -0.0006372326, -0.0004432116, -0.0002481119, 
    -6.803091e-06, 0.0002432357, 0.0004977868, 0.0007134227, 0.0009064168, 
    0.001079911, 0.001239033, 0.001336384, 0.001369121, 0.001402127, 
    0.001377934, 0.001300443, 0.001285222, 0.001264531, 0.001232074, 
    0.001147497, 0.001105365, 0.001108849, 0.001076495, 0.00110943, 
    0.001195757, 0.001209755, 0.001254547, 0.001332063, 0.001487836, 
    0.001651123, 0.001824717, 0.001958383, 0.00208701, 0.002208644, 
    0.002280126, 0.002241737, 0.002097202, 0.002125463, 0.002023048, 
    0.001793474, 0.001370021, 0.0008100793, 0.0001201952, -0.0003233666, 
    -0.00059027, -0.0005284505, -0.0002882284, 0.0004346537, 0.001532182, 
    0.003148638, 0.006278537, 0.01151873, 0.01376125, 0.006880624,
  -0.001132379, -0.0008737884, -0.0006859732, -0.0004800673, -0.0002613944, 
    -2.323341e-05, 0.0002180848, 0.000468364, 0.0006875228, 0.0008836321, 
    0.001054005, 0.001231786, 0.001335185, 0.001365658, 0.001423995, 
    0.001417751, 0.001347818, 0.001346754, 0.001333943, 0.001304782, 
    0.001236107, 0.001197179, 0.001190287, 0.001164522, 0.001191037, 
    0.001262406, 0.001277242, 0.001319156, 0.001389781, 0.001544185, 
    0.001713883, 0.001901236, 0.002026889, 0.002149781, 0.002268262, 
    0.002359393, 0.002335634, 0.002200134, 0.002223169, 0.002123798, 
    0.001904991, 0.00148805, 0.0009616128, 0.0003339484, -3.270161e-05, 
    -0.0002097188, -0.0001720361, 0.0002022309, 0.00125522, 0.002927518, 
    0.005042572, 0.008724133, 0.01456835, 0.01617459, 0.008087293,
  -0.001237005, -0.0009722908, -0.0007961357, -0.0005898924, -0.0003579554, 
    -0.0001250433, 0.0001179136, 0.000375706, 0.0006036986, 0.0008049969, 
    0.0009773837, 0.00117821, 0.001297314, 0.001335898, 0.001423437, 
    0.001441687, 0.001402896, 0.00144635, 0.001459166, 0.001429492, 
    0.001368118, 0.00132148, 0.001296314, 0.001287181, 0.001320849, 
    0.001376438, 0.00138907, 0.001421691, 0.001478848, 0.001621495, 
    0.001788896, 0.001982257, 0.002091268, 0.00219853, 0.002304899, 
    0.002410877, 0.002405277, 0.002289659, 0.002310409, 0.002223786, 
    0.002034805, 0.001664044, 0.00119962, 0.0006462359, 0.0003272909, 
    0.0002307879, 0.000430638, 0.001046959, 0.002409097, 0.004507108, 
    0.007029708, 0.01151915, 0.01813574, 0.01870724, 0.00935362,
  -0.000919334, -0.0007020218, -0.0005617154, -0.0003852486, -0.0001670008, 
    4.418507e-05, 0.0002890368, 0.0005596039, 0.0007954292, 0.0009992233, 
    0.001175845, 0.001404497, 0.001552668, 0.001615471, 0.001740576, 
    0.001783975, 0.001757149, 0.001806697, 0.001811171, 0.001760998, 
    0.001713341, 0.001650691, 0.001578491, 0.001568549, 0.001573617, 
    0.001576831, 0.001574915, 0.001588362, 0.001620845, 0.001732683, 
    0.001880705, 0.002065885, 0.002149343, 0.002255589, 0.00237004, 
    0.002482526, 0.00248496, 0.002394611, 0.002428003, 0.002378823, 
    0.002254913, 0.001972501, 0.001609033, 0.001165888, 0.0009657956, 
    0.0009147286, 0.001287111, 0.002112702, 0.004283091, 0.007257819, 
    0.0106227, 0.01569496, 0.0215774, 0.01867523, 0.009337617,
  -2.291061e-05, 0.0001337056, 0.0002232324, 0.0003308523, 0.0004929426, 
    0.0006747385, 0.0009475438, 0.001260576, 0.001503698, 0.001695822, 
    0.00186781, 0.002135134, 0.002341492, 0.002459415, 0.002642378, 
    0.00272776, 0.002765292, 0.002899603, 0.002940237, 0.00285269, 
    0.002791947, 0.002674359, 0.002519932, 0.002533291, 0.002552143, 
    0.002513055, 0.002490595, 0.002462469, 0.002448435, 0.002500944, 
    0.002612533, 0.002790937, 0.002868995, 0.002947329, 0.003010486, 
    0.003096456, 0.003084557, 0.002988465, 0.00299237, 0.002930979, 
    0.002810503, 0.0025425, 0.002206787, 0.001862209, 0.001877001, 
    0.002125136, 0.002535872, 0.004374673, 0.007384795, 0.01100877, 
    0.01486728, 0.01974851, 0.02203229, 0.01721893, 0.008609463,
  0.001525037, 0.001613775, 0.001650095, 0.001676176, 0.00180754, 
    0.001955889, 0.002213047, 0.002578461, 0.002825206, 0.003000255, 
    0.003165949, 0.003482792, 0.003764559, 0.003955231, 0.004215383, 
    0.004356632, 0.004483921, 0.004745268, 0.004848449, 0.004716865, 
    0.004634322, 0.004440506, 0.004179748, 0.004235786, 0.004303121, 
    0.004240062, 0.004202759, 0.004126547, 0.004060736, 0.004049834, 
    0.004132322, 0.004334128, 0.004459915, 0.004574649, 0.004621266, 
    0.004649409, 0.004570927, 0.004432376, 0.004414596, 0.004363596, 
    0.004290968, 0.004094449, 0.003831839, 0.003499255, 0.003425152, 
    0.003919193, 0.005049448, 0.007604063, 0.01144977, 0.01566713, 
    0.01941046, 0.02178398, 0.0201121, 0.01402752, 0.007013762,
  0.0042406, 0.004304115, 0.004336556, 0.004359812, 0.00442779, 0.004554686, 
    0.004845382, 0.005223786, 0.005469663, 0.005675935, 0.005890472, 
    0.006304897, 0.006639846, 0.006852302, 0.007209828, 0.00741714, 
    0.007554823, 0.007813073, 0.007878774, 0.007693108, 0.007650611, 
    0.007420655, 0.007037286, 0.007063033, 0.007061321, 0.006955535, 
    0.006904439, 0.006782543, 0.006667385, 0.006594906, 0.006652744, 
    0.006892472, 0.007092851, 0.007273855, 0.007322833, 0.007292658, 
    0.007127478, 0.006921462, 0.006893298, 0.00686856, 0.006870956, 
    0.006767666, 0.006587035, 0.006311919, 0.006409517, 0.006760887, 
    0.00874937, 0.01199416, 0.01680782, 0.02086304, 0.02264492, 0.01996762, 
    0.01691298, 0.01122086, 0.005610432,
  0.007229995, 0.007333384, 0.007376099, 0.007374124, 0.007391734, 
    0.00751858, 0.007858753, 0.008320915, 0.00859053, 0.008837112, 
    0.009119868, 0.009694045, 0.01017295, 0.01050224, 0.01106171, 0.01142077, 
    0.01168923, 0.01213182, 0.01229645, 0.01209588, 0.01211143, 0.01183592, 
    0.01131945, 0.01141037, 0.01140234, 0.01113504, 0.01106829, 0.01094481, 
    0.01082342, 0.01072266, 0.01075201, 0.01095058, 0.01105998, 0.01128979, 
    0.01136159, 0.01131676, 0.01108873, 0.01081316, 0.01080122, 0.01082098, 
    0.01091711, 0.01090423, 0.01079269, 0.01053968, 0.01087861, 0.01165328, 
    0.01379676, 0.01793509, 0.02319375, 0.02464772, 0.02080274, 0.01648192, 
    0.01425813, 0.009871193, 0.004935597,
  0.009973269, 0.01016932, 0.01025406, 0.01027068, 0.0102757, 0.01041663, 
    0.0107945, 0.01132856, 0.01163741, 0.01196308, 0.01235872, 0.01312782, 
    0.01376601, 0.01422324, 0.01503889, 0.01559346, 0.01599886, 0.01664954, 
    0.01693929, 0.01676901, 0.01689465, 0.01660962, 0.01596951, 0.01612656, 
    0.01612394, 0.01578466, 0.01575722, 0.01568011, 0.0156195, 0.01558246, 
    0.01572765, 0.01610945, 0.01635516, 0.01659803, 0.01672393, 0.01682548, 
    0.01670238, 0.0164564, 0.01650799, 0.0165345, 0.01666236, 0.01670725, 
    0.01661543, 0.01631758, 0.01693535, 0.01812373, 0.02033529, 0.02502611, 
    0.02800366, 0.02261273, 0.01741166, 0.01339587, 0.01278232, 0.008911146, 
    0.004455573,
  0.01205063, 0.01237908, 0.01252763, 0.01259952, 0.01263075, 0.01279566, 
    0.01320047, 0.01379176, 0.01416002, 0.01459792, 0.0151418, 0.01611879, 
    0.01692211, 0.01751594, 0.01862188, 0.01939889, 0.01993888, 0.02081543, 
    0.02125085, 0.02115286, 0.02142021, 0.02114795, 0.02038603, 0.02058288, 
    0.02053031, 0.02007158, 0.02006952, 0.02005801, 0.02009478, 0.0201681, 
    0.0204963, 0.02113668, 0.0215195, 0.02194195, 0.02229094, 0.02274146, 
    0.02292035, 0.02293807, 0.02329311, 0.02362584, 0.02398693, 0.02408233, 
    0.02397978, 0.02358413, 0.02444851, 0.02576036, 0.02709389, 0.02989145, 
    0.02552739, 0.01955462, 0.01426704, 0.01207616, 0.0116185, 0.00908424, 
    0.00454212,
  0.01345591, 0.01396959, 0.01418254, 0.01431364, 0.01438918, 0.014592, 
    0.01504741, 0.01571199, 0.016159, 0.01671124, 0.01739936, 0.01856648, 
    0.0195273, 0.02025133, 0.02162021, 0.02258639, 0.02321919, 0.02428665, 
    0.02484875, 0.02483899, 0.02522817, 0.0249709, 0.02410379, 0.02428963, 
    0.02413905, 0.02353831, 0.02350171, 0.02353433, 0.02367759, 0.02388621, 
    0.02443745, 0.02537917, 0.02587878, 0.0264755, 0.02708091, 0.02801087, 
    0.02866401, 0.0291349, 0.02987521, 0.03060959, 0.0312787, 0.03133333, 
    0.03107636, 0.03050426, 0.03110855, 0.03145166, 0.02968984, 0.0270404, 
    0.02256152, 0.01684555, 0.01312805, 0.01104056, 0.01184454, 0.009850824, 
    0.004925412,
  0.01391646, 0.01460963, 0.01481633, 0.01500469, 0.01517004, 0.01541229, 
    0.01587976, 0.01657637, 0.01711552, 0.01778105, 0.01857506, 0.01988991, 
    0.02088771, 0.02155761, 0.02310759, 0.02411851, 0.0245946, 0.02575976, 
    0.02640085, 0.02649249, 0.02689028, 0.02662704, 0.0257085, 0.02602875, 
    0.02583658, 0.02508613, 0.02526516, 0.02548069, 0.02574672, 0.02603999, 
    0.02671831, 0.02780405, 0.02832744, 0.02851899, 0.02891721, 0.03006859, 
    0.03107272, 0.03179844, 0.03238302, 0.03285451, 0.03318296, 0.03286161, 
    0.03229239, 0.03151215, 0.03129372, 0.029703, 0.02669277, 0.02405907, 
    0.02014961, 0.01591932, 0.01246452, 0.01213877, 0.01226381, 0.01046252, 
    0.005231262,
  0.01324217, 0.01395377, 0.01402448, 0.01413021, 0.01425608, 0.0144273, 
    0.01478434, 0.01535481, 0.01590069, 0.0165484, 0.01727566, 0.01849833, 
    0.01930226, 0.01970706, 0.02112064, 0.02192885, 0.02206841, 0.02294313, 
    0.02322809, 0.02298205, 0.02299317, 0.0223977, 0.02114929, 0.02088742, 
    0.02009976, 0.01896209, 0.01894186, 0.0191502, 0.01951698, 0.0197135, 
    0.02027602, 0.02115907, 0.02135633, 0.02157856, 0.02200862, 0.0231403, 
    0.02421982, 0.02515709, 0.02592252, 0.02664044, 0.0273109, 0.02755992, 
    0.02755469, 0.02726903, 0.02766238, 0.0265469, 0.023751, 0.021886, 
    0.01897426, 0.01611016, 0.0142495, 0.01314069, 0.01260045, 0.01095599, 
    0.005477995,
  0.01220439, 0.0127975, 0.01273553, 0.01268674, 0.01263938, 0.0126763, 
    0.01286857, 0.01324313, 0.01360265, 0.01404259, 0.01453967, 0.01543478, 
    0.01596513, 0.01615811, 0.01719342, 0.01765632, 0.01747756, 0.01800779, 
    0.0179182, 0.01727519, 0.01687995, 0.01598083, 0.01453429, 0.0140091, 
    0.01311806, 0.01200434, 0.01191627, 0.01212117, 0.01256326, 0.01272503, 
    0.01327508, 0.01417594, 0.01451641, 0.01504589, 0.01585, 0.01732974, 
    0.01874555, 0.02003984, 0.02109702, 0.02222229, 0.02342933, 0.02415786, 
    0.02443594, 0.02424473, 0.02498777, 0.02422079, 0.02190466, 0.0205316, 
    0.01956356, 0.01819685, 0.01568841, 0.0139535, 0.01274214, 0.01095599, 
    0.005477995,
  0.009916167, 0.01016196, 0.009694543, 0.009409444, 0.00927501, 0.009050101, 
    0.009100439, 0.009478839, 0.009967448, 0.01057953, 0.01128467, 
    0.01227903, 0.01283086, 0.01295574, 0.01405224, 0.0142856, 0.0136162, 
    0.01368473, 0.0130423, 0.01173431, 0.01061521, 0.009164579, 0.00734896, 
    0.006323426, 0.005145693, 0.003929531, 0.003827904, 0.004116658, 
    0.004750577, 0.005088976, 0.005950906, 0.007318707, 0.008147624, 
    0.009088684, 0.01018193, 0.0119862, 0.01389515, 0.01587345, 0.01761157, 
    0.01930581, 0.02099949, 0.02221997, 0.02281038, 0.02275205, 0.0237027, 
    0.02338121, 0.0218955, 0.02173654, 0.02101775, 0.01980311, 0.01632995, 
    0.01397629, 0.01274214, 0.01095599, 0.005477995,
  0.00380238, 0.003394623, 0.002320348, 0.001682671, 0.001457854, 
    0.0009705022, 0.0009730479, 0.001502685, 0.002657045, 0.003910207, 
    0.005241344, 0.006914776, 0.007782926, 0.007856324, 0.009362484, 
    0.00969774, 0.008843089, 0.008901197, 0.008120545, 0.006512391, 
    0.004923839, 0.003097245, 0.00102271, -0.0002167651, -0.001130232, 
    -0.001675119, -0.001194192, -0.0001685533, 0.001401795, 0.002889352, 
    0.004829013, 0.007220779, 0.009016003, 0.01067656, 0.01220246, 
    0.01416237, 0.01593751, 0.01752785, 0.01931088, 0.02100157, 0.02259992, 
    0.0238352, 0.02429009, 0.02396456, 0.0246055, 0.02416566, 0.02264506, 
    0.02232842, 0.0213811, 0.01980311, 0.01632995, 0.01397629, 0.01274214, 
    0.01095599, 0.005477995 ;

 u_north =
  0.0007923699, 0.000817284, 0.0008270862, 0.0007784893, 0.0006235225, 
    0.0005948534, 0.0005526033, 0.0004868061, 0.000472589, 0.0004239023, 
    0.0003354909, 0.0001829801, 7.403502e-05, 3.400862e-05, 5.058293e-05, 
    0.0001491776, 0.0003020245, 0.0004128614, 0.0004074894, 0.0002523101, 
    0.0001017511, -4.95348e-05, -0.0006617901, -0.001697982, -0.002800554, 
    -0.00371915, -0.004399224, 1.734723e-18, -1.734723e-18, -8.673617e-19, 
    -1.734723e-18, -1.734723e-18, -8.673617e-19, 0, 8.673617e-19, 
    -8.673617e-19, -1.734723e-18, 1.734723e-18, -8.673617e-19, 8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.0007577727, 0.0007851875, 0.0008083834, 0.000732062, 0.0005713456, 
    0.000534724, 0.000476676, 0.00039199, 0.0003234863, 0.00023209, 
    0.0001285757, -4.099279e-05, -0.0001171951, -0.000104304, -9.427591e-05, 
    -1.540274e-05, 0.0001411811, 0.0002655799, 0.0002678712, 0.0001436882, 
    7.507227e-05, -0.0001641513, -0.0009015528, -0.00198876, -0.00306848, 
    -0.003837887, -0.004584889, 1.734723e-18, -1.734723e-18, -8.673617e-19, 
    -1.734723e-18, -1.734723e-18, -8.673617e-19, 0, 8.673617e-19, 
    -8.673617e-19, -1.734723e-18, 1.734723e-18, -8.673617e-19, 8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.0007347957, 0.000759922, 0.0007745048, 0.0006917988, 0.0005303793, 
    0.0004857077, 0.0004188395, 0.0003260413, 0.0002450331, 0.0001657006, 
    9.124844e-05, -7.685324e-05, -0.0001578879, -0.0001557657, -0.0001953209, 
    -0.0001490266, -8.769965e-06, 9.940141e-05, 0.0001206112, 5.0863e-05, 
    -6.395997e-05, -0.0003428875, -0.001218685, -0.002305605, -0.003300061, 
    -0.003939493, -0.004903315, 1.734723e-18, -1.734723e-18, -8.673617e-19, 
    -1.734723e-18, -1.734723e-18, -8.673617e-19, 0, 8.673617e-19, 
    -8.673617e-19, -1.734723e-18, 1.734723e-18, -8.673617e-19, 8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.0007271148, 0.0007403136, 0.0007446103, 0.0006684425, 0.0005131828, 
    0.0004594173, 0.0003818912, 0.0002792635, 0.0001919071, 0.0001175598, 
    5.91706e-05, -0.0001076707, -0.0001928584, -0.0002194646, -0.0003038275, 
    -0.0002840881, -0.0001578483, -5.590045e-05, -2.476515e-05, 
    -9.217853e-05, -0.0001849339, -0.0005603491, -0.001531979, -0.00257803, 
    -0.003499252, -0.004038735, -0.005238381, 1.734723e-18, -1.734723e-18, 
    -8.673617e-19, -1.734723e-18, -1.734723e-18, -8.673617e-19, 0, 
    8.673617e-19, -8.673617e-19, -1.734723e-18, 1.734723e-18, -8.673617e-19, 
    8.673617e-19, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18,
  0.0007247951, 0.0007304493, 0.0007406196, 0.0006621311, 0.0005002494, 
    0.0004366276, 0.0003498625, 0.0002387139, 0.0001474097, 7.285636e-05, 
    1.096149e-05, -0.0001712332, -0.0002842081, -0.0003334954, -0.0004287961, 
    -0.0004297041, -0.0003340015, -0.0002374431, -0.0001960901, 
    -0.0002355974, -0.0002907356, -0.0007488872, -0.001803645, -0.002814319, 
    -0.003672092, -0.004188772, -0.005529669, 1.734723e-18, -1.734723e-18, 
    -8.673617e-19, -1.734723e-18, -1.734723e-18, -8.673617e-19, 0, 
    8.673617e-19, -8.673617e-19, -1.734723e-18, 1.734723e-18, -8.673617e-19, 
    8.673617e-19, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18,
  0.000755029, 0.0007441391, 0.0007433011, 0.0006565884, 0.0004924946, 
    0.0004264668, 0.0003360343, 0.0002201832, 0.0001161303, 2.803257e-05, 
    -4.705206e-05, -0.0002373126, -0.000364464, -0.0004336439, -0.0005385512, 
    -0.000557593, -0.0004887096, -0.0003968841, -0.0003465577, -0.0003615579, 
    -0.000481445, -0.000914495, -0.002042309, -0.003026623, -0.003784398, 
    -0.00432077, -0.005786249, 1.734723e-18, -1.734723e-18, -8.673617e-19, 
    -1.734723e-18, -1.734723e-18, -8.673617e-19, 0, 8.673617e-19, 
    -8.673617e-19, -1.734723e-18, 1.734723e-18, -8.673617e-19, 8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.000782082, 0.0007563885, 0.0007457006, 0.0006684189, 0.0005068356, 
    0.0004311332, 0.0003306456, 0.0002044287, 8.814029e-05, -1.207766e-05, 
    -9.896532e-05, -0.0002964439, -0.0004362814, -0.0005232629, 
    -0.0006489232, -0.0006860312, -0.0006271522, -0.0005395616, 
    -0.0004812056, -0.0005107815, -0.000652112, -0.00123331, -0.002308901, 
    -0.003236853, -0.003881967, -0.004439086, -0.006762284, 1.734723e-18, 
    -1.734723e-18, -8.673617e-19, -1.734723e-18, -1.734723e-18, 
    -8.673617e-19, 0, 8.673617e-19, -8.673617e-19, -1.734723e-18, 
    1.734723e-18, -8.673617e-19, 8.673617e-19, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.0008118179, 0.0007761438, 0.000774015, 0.0006902638, 0.0005199967, 
    0.0004354156, 0.0003257002, 0.0001899701, 6.245272e-05, -4.888854e-05, 
    -0.0001529142, -0.0003745096, -0.0005528391, -0.0006938612, 
    -0.0008483311, -0.0009133227, -0.0008866079, -0.0007813445, -0.00070517, 
    -0.0006792739, -0.00080875, -0.001535065, -0.002569652, -0.003429884, 
    -0.003971586, -0.004547825, -0.00859932, 1.734723e-18, -1.734723e-18, 
    -8.673617e-19, -1.734723e-18, -1.734723e-18, -8.673617e-19, 0, 
    8.673617e-19, -8.673617e-19, -1.734723e-18, 1.734723e-18, -8.673617e-19, 
    8.673617e-19, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18,
  0.0008796112, 0.0008214272, 0.0008057513, 0.0007109475, 0.0005324584, 
    0.0004394704, 0.0003229334, 0.000177677, 3.103473e-05, -0.0001070467, 
    -0.0002424808, -0.0004853714, -0.0006903268, -0.0008628963, -0.001037147, 
    -0.001128541, -0.001135003, -0.001025495, -0.0009201878, -0.000838817, 
    -0.0009603202, -0.001820813, -0.002816593, -0.003612719, -0.00405649, 
    -0.004742833, -0.01034163, 1.734723e-18, -1.734723e-18, -8.673617e-19, 
    -1.734723e-18, -1.734723e-18, -8.673617e-19, 0, 8.673617e-19, 
    -8.673617e-19, -1.734723e-18, 1.734723e-18, -8.673617e-19, 8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.0009460427, 0.000865801, 0.0008368502, 0.0007350745, 0.0005580416, 
    0.0004585772, 0.0003289147, 0.0001671105, -2.697324e-06, -0.0001666552, 
    -0.0003302497, -0.0005940081, -0.0008250551, -0.001028539, -0.001222173, 
    -0.00133944, -0.001378413, -0.001264746, -0.00113089, -0.0009951588, 
    -0.00131935, -0.002100835, -0.003058594, -0.003791906, -0.004159981, 
    -0.005007484, -0.01205005, 1.734723e-18, -1.734723e-18, -8.673617e-19, 
    -1.734723e-18, -1.734723e-18, -8.673617e-19, 0, 8.673617e-19, 
    -8.673617e-19, -1.734723e-18, 1.734723e-18, -8.673617e-19, 8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.001013265, 0.0009107029, 0.0008858715, 0.0007841222, 0.0005911103, 
    0.0004792677, 0.0003349672, 0.0001564183, -3.683052e-05, -0.0002269725, 
    -0.0004190622, -0.0007039366, -0.0009613853, -0.001203985, -0.001435997, 
    -0.001582818, -0.001642296, -0.001515428, -0.001371324, -0.001291929, 
    -0.001682646, -0.002432317, -0.003311391, -0.00395242, -0.004358868, 
    -0.005275222, -0.01355297, 1.734723e-18, -1.734723e-18, -8.673617e-19, 
    -1.734723e-18, -1.734723e-18, -8.673617e-19, 0, 8.673617e-19, 
    -8.673617e-19, -1.734723e-18, 1.734723e-18, -8.673617e-19, 8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.001139275, 0.001004245, 0.0009573225, 0.0008349374, 0.0006253707, 
    0.0005007038, 0.0003412378, 0.0001453409, -7.184017e-05, -0.0002950015, 
    -0.0005310008, -0.0008589207, -0.001172726, -0.001477188, -0.001746517, 
    -0.001933832, -0.002037173, -0.00195951, -0.001821036, -0.001696441, 
    -0.002059018, -0.002807996, -0.003596774, -0.004097546, -0.004564842, 
    -0.005552428, -0.01388821, 1.734723e-18, -1.734723e-18, -8.673617e-19, 
    -1.734723e-18, -1.734723e-18, -8.673617e-19, 0, 8.673617e-19, 
    -8.673617e-19, -1.734723e-18, 1.734723e-18, -8.673617e-19, 8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.001280457, 0.001103685, 0.00103209, 0.0008930531, 0.0006862176, 
    0.0005523817, 0.0003760105, 0.000155645, -0.0001064108, -0.0003800821, 
    -0.0006713304, -0.001043018, -0.0014055, -0.001763063, -0.002071439, 
    -0.002301127, -0.002450366, -0.00242419, -0.002291608, -0.002119713, 
    -0.002483399, -0.003201077, -0.003895353, -0.004249365, -0.004780272, 
    -0.008019906, -0.01423852, 1.734723e-18, -1.734723e-18, -8.673617e-19, 
    -1.734723e-18, -1.734723e-18, -8.673617e-19, 0, 8.673617e-19, 
    -8.673617e-19, -1.734723e-18, 1.734723e-18, -8.673617e-19, 8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.001461133, 0.00124306, 0.00117415, 0.001030465, 0.0007859547, 
    0.0006265747, 0.0004205502, 0.0001665943, -0.000142375, -0.000468592, 
    -0.0008173161, -0.001234536, -0.001647656, -0.002052275, -0.002399136, 
    -0.002678257, -0.002881602, -0.002904269, -0.002777569, -0.002574345, 
    -0.002974335, -0.003635918, -0.004203479, -0.004453904, -0.005201587, 
    -0.01231416, -0.01664259, 1.734723e-18, -1.734723e-18, -8.673617e-19, 
    -1.734723e-18, -1.734723e-18, -8.673617e-19, 0, 8.673617e-19, 
    -8.673617e-19, -1.734723e-18, 1.734723e-18, -8.673617e-19, 8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.001772599, 0.001478025, 0.0013598, 0.00117049, 0.0008922124, 
    0.0007363827, 0.0005251405, 0.0002615471, -8.325063e-05, -0.0004571292, 
    -0.0008590419, -0.00132669, -0.00180298, -0.002292246, -0.002698345, 
    -0.003046004, -0.00332828, -0.003365824, -0.003253537, -0.003054349, 
    -0.003474599, -0.004127888, -0.004473847, -0.004854445, -0.005728836, 
    -0.01630226, -0.02470552, 1.734723e-18, -1.734723e-18, -8.673617e-19, 
    -1.734723e-18, -1.734723e-18, -8.673617e-19, 0, 8.673617e-19, 
    -8.673617e-19, -1.734723e-18, 1.734723e-18, -8.673617e-19, 8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.002143057, 0.001782857, 0.001684341, 0.0015238, 0.001243885, 0.001046448, 
    0.0007885303, 0.0004727186, 6.235077e-05, -0.0003826601, -0.0008614304, 
    -0.001400484, -0.001955127, -0.002525231, -0.002974105, -0.003392901, 
    -0.003763629, -0.003821226, -0.003721268, -0.003531003, -0.004036615, 
    -0.00461812, -0.004740621, -0.005263472, -0.009078053, -0.01733181, 
    -0.0306591, 1.734723e-18, -1.734723e-18, -8.673617e-19, -1.734723e-18, 
    -1.734723e-18, -8.673617e-19, 0, 8.673617e-19, -8.673617e-19, 
    -1.734723e-18, 1.734723e-18, -8.673617e-19, 8.673617e-19, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.002807974, 0.002337314, 0.00215689, 0.001919389, 0.001665109, 
    0.001476247, 0.001216934, 0.0008962456, 0.0004504924, -4.724534e-05, 
    -0.0005868798, -0.00118686, -0.001816874, -0.002480911, -0.003037012, 
    -0.003561597, -0.004039816, -0.004146595, -0.004111782, -0.003991753, 
    -0.004578627, -0.005118464, -0.00531142, -0.006056207, -0.01681793, 
    -0.0200562, -0.02978524, 1.734723e-18, -1.734723e-18, -8.673617e-19, 
    -1.734723e-18, -1.734723e-18, -8.673617e-19, 0, 8.673617e-19, 
    -8.673617e-19, -1.734723e-18, 1.734723e-18, -8.673617e-19, 8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.003717132, 0.003149544, 0.002987836, 0.002791354, 0.00246554, 
    0.002224908, 0.001906078, 0.001516378, 0.0009929048, 0.000406944, 
    -0.0001963982, -0.000851398, -0.001552971, -0.002305179, -0.002973383, 
    -0.003619655, -0.004216559, -0.004404328, -0.004450208, -0.004411738, 
    -0.0051369, -0.005796185, -0.005984565, -0.009702701, -0.01997573, 
    -0.02526997, -0.02770307, 1.734723e-18, -1.734723e-18, -8.673617e-19, 
    -1.734723e-18, -1.734723e-18, -8.673617e-19, 0, 8.673617e-19, 
    -8.673617e-19, -1.734723e-18, 1.734723e-18, -8.673617e-19, 8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.004830108, 0.004148448, 0.004030267, 0.003911112, 0.003631681, 
    0.003409915, 0.003092373, 0.002692365, 0.002123805, 0.001453137, 
    0.0006967676, -0.0001015505, -0.0009555044, -0.001868312, -0.002724808, 
    -0.003518688, -0.004228224, -0.004544693, -0.004713247, -0.004784698, 
    -0.005918164, -0.006717572, -0.006942309, -0.0180254, -0.02415873, 
    -0.02459628, -0.02245573, 1.734723e-18, -1.734723e-18, -8.673617e-19, 
    -1.734723e-18, -1.734723e-18, -8.673617e-19, 0, 8.673617e-19, 
    -8.673617e-19, -1.734723e-18, 1.734723e-18, -8.673617e-19, 8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.006582706, 0.005768403, 0.005526529, 0.005318936, 0.005092982, 
    0.00490366, 0.00459774, 0.004194317, 0.003580973, 0.002804746, 
    0.001887501, 0.0009690775, -2.584135e-05, -0.001101366, -0.002335465, 
    -0.003396103, -0.004244076, -0.004956171, -0.005374456, -0.005577446, 
    -0.007036692, -0.008544928, -0.01183997, -0.01960102, -0.03122979, 
    -0.0219474, -0.0180191, 1.734723e-18, -1.734723e-18, -8.673617e-19, 
    -1.734723e-18, -1.734723e-18, -8.673617e-19, 0, 8.673617e-19, 
    -8.673617e-19, -1.734723e-18, 1.734723e-18, -8.673617e-19, 8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.008649814, 0.007708583, 0.007502823, 0.007322053, 0.00699451, 
    0.006775029, 0.006472251, 0.006060074, 0.005389749, 0.004465453, 
    0.00330592, 0.002241496, 0.001075861, -0.0001976394, -0.00210019, 
    -0.003582054, -0.004575902, -0.006041064, -0.006831541, -0.007086141, 
    -0.009182456, -0.011725, -0.01460237, -0.02797914, -0.02953572, 
    -0.0164191, -0.01473739, 1.734723e-18, -1.734723e-18, -8.673617e-19, 
    -1.734723e-18, -1.734723e-18, -8.673617e-19, 0, 8.673617e-19, 
    -8.673617e-19, -1.734723e-18, 1.734723e-18, -8.673617e-19, 8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.01097025, 0.009891913, 0.009702652, 0.009559275, 0.009264504, 
    0.009117412, 0.008794631, 0.008314564, 0.007519744, 0.006382752, 
    0.004878038, 0.003660603, 0.002312554, 0.0008244152, -0.002046866, 
    -0.004113833, -0.005284836, -0.00789717, -0.009117732, -0.009089692, 
    -0.0118186, -0.01469178, -0.01960233, -0.02981065, -0.02435168, 
    -0.01187208, -0.01207916, 1.734723e-18, -1.734723e-18, -8.673617e-19, 
    -1.734723e-18, -1.734723e-18, -8.673617e-19, 0, 8.673617e-19, 
    -8.673617e-19, -1.734723e-18, 1.734723e-18, -8.673617e-19, 8.673617e-19, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.01348132, 0.01225971, 0.01207692, 0.01195273, 0.0116751, 0.01163371, 
    0.0113932, 0.01097651, 0.01008885, 0.008624393, 0.00659745, 0.005235378, 
    0.003712758, 0.002025406, -0.002035989, -0.004811064, -0.006210077, 
    -0.01027168, -0.01188782, -0.01116273, -0.01427396, -0.02027029, 
    -0.02418665, -0.02604485, -0.01858695, -0.008095913, -0.009767345, 
    1.734723e-18, -1.734723e-18, -8.673617e-19, -1.734723e-18, -1.734723e-18, 
    -8.673617e-19, 0, 8.673617e-19, -8.673617e-19, -1.734723e-18, 
    1.734723e-18, -8.673617e-19, 8.673617e-19, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.016164, 0.01478561, 0.01453576, 0.01434542, 0.01402466, 0.01409778, 
    0.01396358, 0.01364716, 0.01264543, 0.01086765, 0.008295567, 0.006699102, 
    0.004975987, 0.003161492, -0.001927144, -0.005196725, -0.006654313, 
    -0.01200454, -0.01466833, -0.01601175, -0.02267131, -0.02541151, 
    -0.02098996, -0.01917402, -0.01409907, -0.005040115, -0.007806812, 
    1.734723e-18, -1.734723e-18, -8.673617e-19, -1.734723e-18, -1.734723e-18, 
    -8.673617e-19, 0, 8.673617e-19, -8.673617e-19, -1.734723e-18, 
    1.734723e-18, -8.673617e-19, 8.673617e-19, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.01761203, 0.01602501, 0.01511892, 0.01421, 0.0134849, 0.01344967, 
    0.01323451, 0.01282945, 0.01177323, 0.009929067, 0.007515062, 
    0.006398823, 0.005266316, 0.004043475, -0.001142381, -0.004435841, 
    -0.005769091, -0.01189872, -0.01710721, -0.02108076, -0.02320697, 
    -0.0214313, -0.01333039, -0.01385473, -0.01058535, -0.001987682, 
    -0.006241117, 1.734723e-18, -1.734723e-18, -8.673617e-19, -1.734723e-18, 
    -1.734723e-18, -8.673617e-19, 0, 8.673617e-19, -8.673617e-19, 
    -1.734723e-18, 1.734723e-18, -8.673617e-19, 8.673617e-19, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.0172986, 0.01584073, 0.015683, 0.01565781, 0.01548363, 0.01566052, 
    0.01566791, 0.01554025, 0.01460173, 0.01302335, 0.0108669, 0.0101677, 
    0.009413297, 0.008243903, 0.003221271, -0.0003937466, -0.002452062, 
    -0.009053649, -0.01377161, -0.01590957, -0.01635998, -0.01302242, 
    -0.007219801, -0.009713696, -0.007470636, 0.0004386415, -0.004979648, 
    1.734723e-18, -1.734723e-18, -8.673617e-19, -1.734723e-18, -1.734723e-18, 
    -8.673617e-19, 0, 8.673617e-19, -8.673617e-19, -1.734723e-18, 
    1.734723e-18, -8.673617e-19, 8.673617e-19, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.02241537, 0.02101998, 0.02173685, 0.0226208, 0.02300152, 0.02361992, 
    0.0241075, 0.0245438, 0.02407481, 0.02289972, 0.02113479, 0.02069732, 
    0.01975361, 0.01830086, 0.01250535, 0.008443368, 0.006217245, 
    -0.0008391172, -0.005141106, -0.00620944, -0.007936591, -0.006333036, 
    -0.002295462, -0.006174934, -0.004908859, 0.002391743, -0.004625074, 
    1.734723e-18, -1.734723e-18, -8.673617e-19, -1.734723e-18, -1.734723e-18, 
    -8.673617e-19, 0, 8.673617e-19, -8.673617e-19, -1.734723e-18, 
    1.734723e-18, -8.673617e-19, 8.673617e-19, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.03162368, 0.03033546, 0.0316451, 0.03289506, 0.033356, 0.03428645, 
    0.03500626, 0.03557833, 0.03519425, 0.03405667, 0.03228532, 0.031621, 
    0.03044583, 0.02876497, 0.02217277, 0.01759446, 0.01512472, 0.007326108, 
    0.002687077, 0.001433556, -0.001226424, -0.0007498109, 0.002149783, 
    -0.003233554, -0.002832841, 0.002923594, -0.004625074, 1.734723e-18, 
    -1.734723e-18, -8.673617e-19, -1.734723e-18, -1.734723e-18, 
    -8.673617e-19, 0, 8.673617e-19, -8.673617e-19, -1.734723e-18, 
    1.734723e-18, -8.673617e-19, 8.673617e-19, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.04402607, 0.04283758, 0.04468332, 0.04609592, 0.04638866, 0.04757839, 
    0.04840134, 0.04891919, 0.04845141, 0.04724553, 0.0454129, 0.04437114, 
    0.04283102, 0.04079298, 0.03314729, 0.02785552, 0.02500861, 0.01624787, 
    0.01077858, 0.008726324, 0.005448233, 0.004680289, 0.005881156, 
    -0.001426912, -0.002613442, 0.002923594, -0.004625074, 1.734723e-18, 
    -1.734723e-18, -8.673617e-19, -1.734723e-18, -1.734723e-18, 
    -8.673617e-19, 0, 8.673617e-19, -8.673617e-19, -1.734723e-18, 
    1.734723e-18, -8.673617e-19, 8.673617e-19, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.0604593, 0.05912908, 0.06056419, 0.06087698, 0.06006747, 0.06105214, 
    0.06155799, 0.06158503, 0.06072105, 0.05919665, 0.05701184, 0.05531149, 
    0.05312408, 0.05044961, 0.04172389, 0.03582297, 0.03274684, 0.02327293, 
    0.01695393, 0.01378983, 0.009391731, 0.006956183, 0.006483187, 
    -0.001426912, -0.002613442, 0.002923594, -0.004625074, 1.734723e-18, 
    -1.734723e-18, -8.673617e-19, -1.734723e-18, -1.734723e-18, 
    -8.673617e-19, 0, 8.673617e-19, -8.673617e-19, -1.734723e-18, 
    1.734723e-18, -8.673617e-19, 8.673617e-19, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 3.469447e-18, 
    3.469447e-18, 3.469447e-18, 3.469447e-18,
  0.0001216497, 0.0001405254, 0.0001967185, 0.0002656978, 0.0003831011, 
    0.0004159177, 0.0004504895, 0.0005010087, 0.0005183161, 0.0005437832, 
    0.0005412099, 0.0006022652, 0.0006673236, 0.000737133, 0.0006469135, 
    0.00059919, 0.0006073394, 0.0005936912, 0.0005905931, 0.0006045277, 
    0.0006863389, 0.0008403345, 0.0009095875, 0.000390181, -0.0007514646, 
    -0.001652375, -0.002211781, 1.734723e-18, 8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -2.602085e-18, 0, 0, -8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -8.673617e-19, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.0001197009, 0.0001658031, 0.0002150354, 0.0002507666, 0.0003256972, 
    0.0003404797, 0.0003769687, 0.0004377062, 0.0005824295, 0.000650466, 
    0.0006016846, 0.000660751, 0.0007144849, 0.0007635298, 0.0006970453, 
    0.0006772856, 0.0006914221, 0.0006591171, 0.0006454094, 0.000652048, 
    0.0008063577, 0.000827739, 0.0009488039, 0.0001383949, -0.001011, 
    -0.001728506, -0.002312623, 1.734723e-18, 8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -2.602085e-18, 0, 0, -8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -8.673617e-19, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.000101238, 0.0001545156, 0.0001611085, 0.0001906173, 0.0002669042, 
    0.0002782265, 0.0003179414, 0.0003811619, 0.0005472942, 0.0006137916, 
    0.0005887611, 0.0006441128, 0.0006954033, 0.0007432215, 0.0007364203, 
    0.0007521337, 0.0007786221, 0.0007318552, 0.0007026668, 0.0006926576, 
    0.000784751, 0.000866247, 0.0007545815, -0.0001984692, -0.001233461, 
    -0.001793654, -0.002555619, 1.734723e-18, 8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -2.602085e-18, 0, 0, -8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -8.673617e-19, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  6.866513e-05, 0.0001128166, 0.0001117275, 0.0001467592, 0.0002301533, 
    0.0002395245, 0.0002740924, 0.0003309621, 0.0004908477, 0.0005705917, 
    0.000577655, 0.0006298144, 0.0006790051, 0.0007075765, 0.0007192778, 
    0.0007560782, 0.0008118741, 0.0007728125, 0.0007286884, 0.0006753518, 
    0.0007645948, 0.0009382825, 0.0005050459, -0.0004881081, -0.001424808, 
    -0.00185253, -0.002824656, 1.734723e-18, 8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -2.602085e-18, 0, 0, -8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -8.673617e-19, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  4.327691e-05, 8.124183e-05, 8.341987e-05, 0.0001184467, 0.0001998055, 
    0.0002059758, 0.0002360819, 0.0002874462, 0.0004416521, 0.0005267928, 
    0.0005415331, 0.0005730983, 0.0005994575, 0.0006217287, 0.0006317056, 
    0.0006743241, 0.0007439386, 0.0007273816, 0.0006954581, 0.0006443296, 
    0.0007477165, 0.001000737, 0.0002886663, -0.0007393273, -0.001590842, 
    -0.001918864, -0.003058541, 1.734723e-18, 8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -2.602085e-18, 0, 0, -8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -8.673617e-19, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  4.348567e-05, 6.783746e-05, 6.265133e-05, 9.358254e-05, 0.0001748018, 
    0.0001806477, 0.0002075981, 0.0002525739, 0.0003971202, 0.000476437, 
    0.0004894523, 0.0005109497, 0.0005295636, 0.0005463322, 0.0005547943, 
    0.0006025225, 0.0006842738, 0.0006874816, 0.0006662733, 0.0006170837, 
    0.000795432, 0.001055595, 9.857253e-05, -0.0009609148, -0.001664796, 
    -0.001977223, -0.003264559, 1.734723e-18, 8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -2.602085e-18, 0, 0, -8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -8.673617e-19, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  4.367244e-05, 5.584336e-05, 4.406764e-05, 8.040923e-05, 0.0001621638, 
    0.0001637576, 0.0001845026, 0.0002215311, 0.0003572714, 0.0004313764, 
    0.0004428478, 0.000455336, 0.0004670187, 0.0004788628, 0.0004756214, 
    0.0005263413, 0.0006308819, 0.0006517767, 0.0006401569, 0.0005935249, 
    0.0008381329, 0.0008687362, -0.0001748793, -0.001162887, -0.001725534, 
    -0.002029533, -0.003689348, 1.734723e-18, 8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -2.602085e-18, 0, 0, -8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -8.673617e-19, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  4.696667e-05, 5.008612e-05, 4.243934e-05, 7.425967e-05, 0.0001505657, 
    0.0001482571, 0.0001633072, 0.0001930419, 0.0003207005, 0.0003900224, 
    0.0003952379, 0.0003851558, 0.0003671053, 0.0003398704, 0.0003194188, 
    0.0003631588, 0.000466841, 0.000516502, 0.0005416174, 0.0005726141, 
    0.0008773237, 0.0006846192, -0.000457145, -0.001348334, -0.001781321, 
    -0.002077609, -0.004382601, 1.734723e-18, 8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -2.602085e-18, 0, 0, -8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -8.673617e-19, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  7.841572e-05, 6.102568e-05, 4.380893e-05, 6.843697e-05, 0.0001395839, 
    0.0001335804, 0.0001419425, 0.000158526, 0.0002704966, 0.0003254199, 
    0.0003206114, 0.0002889834, 0.0002497291, 0.000201716, 0.0001715134, 
    0.0002086443, 0.0003091508, 0.0003743506, 0.0004461254, 0.0005528139, 
    0.000911003, 0.0005102691, -0.0007244613, -0.001523987, -0.001834175, 
    -0.002207317, -0.005040107, 1.734723e-18, 8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -2.602085e-18, 0, 0, -8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -8.673617e-19, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.0001092331, 7.174551e-05, 4.515102e-05, 6.430291e-05, 0.0001313936, 
    0.0001185907, 0.0001151257, 0.0001167145, 0.0002148342, 0.000259254, 
    0.0002474828, 0.0001947413, 0.0001347086, 6.633406e-05, 2.657611e-05, 
    5.723051e-05, 0.0001546253, 0.0002350521, 0.0003525499, 0.000533411, 
    0.0007231027, 0.0003394128, -0.00098643, -0.001696136, -0.001892908, 
    -0.002401823, -0.005684824, 1.734723e-18, 8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -2.602085e-18, 0, 0, -8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -8.673617e-19, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.0001404171, 8.259289e-05, 5.565808e-05, 7.015742e-05, 0.0001244869, 
    0.0001033682, 8.799005e-05, 7.440565e-05, 0.00015851, 0.0001923012, 
    0.0001734846, 9.937862e-05, 1.832057e-05, -7.905555e-05, -0.0001502088, 
    -0.0001329002, -2.580445e-05, 8.813163e-05, 0.0002420339, 0.0004082877, 
    0.0005329698, 4.675077e-05, -0.001252837, -0.001828872, -0.001984576, 
    -0.002598599, -0.006285734, 1.734723e-18, 8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -2.602085e-18, 0, 0, -8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -8.673617e-19, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.000212209, 0.0001212806, 7.731599e-05, 7.622292e-05, 0.0001173314, 
    8.759725e-05, 5.987669e-05, 3.057258e-05, 9.962269e-05, 0.0001177066, 
    8.027384e-05, -3.631056e-05, -0.0001710839, -0.0003277783, -0.0004341773, 
    -0.0004516639, -0.00037903, -0.0001919995, 1.10022e-05, 0.0002048059, 
    0.000335993, -0.000336711, -0.001532761, -0.001924227, -0.002079511, 
    -0.002802332, -0.00662903, 1.734723e-18, 8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -2.602085e-18, 0, 0, -8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -8.673617e-19, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.0002944881, 0.0001626736, 9.997922e-05, 8.636821e-05, 0.0001282321, 
    9.149461e-05, 4.757687e-05, -7.446233e-06, 3.488271e-05, 2.652676e-05, 
    -3.653029e-05, -0.0001979815, -0.0003806999, -0.0005880378, 
    -0.0007313169, -0.0007852124, -0.0007486393, -0.0004851242, 
    -0.0002307455, -8.112764e-06, 2.519316e-05, -0.000737934, -0.001825629, 
    -0.002023979, -0.002178804, -0.003768042, -0.006987771, 1.734723e-18, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -2.602085e-18, 0, 0, 
    -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -8.673617e-19, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18,
  0.0004078671, 0.0002340546, 0.0001739439, 0.0001561153, 0.0001663819, 
    0.0001098034, 3.985872e-05, -4.691475e-05, -3.246688e-05, -6.832833e-05, 
    -0.0001580423, -0.0003661682, -0.0005987636, -0.0008539372, -0.00103749, 
    -0.001138083, -0.00114589, -0.0008087151, -0.000519628, -0.0003519964, 
    -0.0004674963, -0.001160206, -0.002124159, -0.002147533, -0.002479491, 
    -0.005370804, -0.007790792, 1.734723e-18, 8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -2.602085e-18, 0, 0, -8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -8.673617e-19, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.0006296312, 0.0003800715, 0.000281375, 0.0002271889, 0.0002096261, 
    0.0001613829, 8.944495e-05, -5.896446e-06, -4.961849e-06, -6.099244e-05, 
    -0.0001724142, -0.0004360098, -0.0007408672, -0.001092443, -0.001339588, 
    -0.001517266, -0.001616989, -0.001293396, -0.001015104, -0.000845496, 
    -0.0009695465, -0.001599726, -0.002320026, -0.002355021, -0.002884041, 
    -0.006927922, -0.009795765, 1.734723e-18, 8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -2.602085e-18, 0, 0, -8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -8.673617e-19, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.0009056347, 0.0005901636, 0.0005178381, 0.0004990619, 0.0004862326, 
    0.0004065297, 0.0002938715, 0.0001485041, 0.0001097973, 1.08787e-05, 
    -0.0001469223, -0.0004880225, -0.0008801023, -0.001324434, -0.001619455, 
    -0.001876305, -0.002077076, -0.001771615, -0.001500257, -0.001319869, 
    -0.001464122, -0.002021197, -0.002513289, -0.002574765, -0.004061291, 
    -0.007893029, -0.01148459, 1.734723e-18, 8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -2.602085e-18, 0, 0, -8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -8.673617e-19, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.00145169, 0.001029461, 0.0008941709, 0.0008136525, 0.0008341572, 
    0.0007736271, 0.0006662837, 0.0005181044, 0.0004700458, 0.000345472, 
    0.0001543778, -0.0002598975, -0.0007460011, -0.001309486, -0.001698958, 
    -0.002065117, -0.002393183, -0.002091879, -0.001856315, -0.00173449, 
    -0.001930369, -0.002331706, -0.00285971, -0.003223648, -0.006434824, 
    -0.009072081, -0.01214086, 1.734723e-18, 8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -2.602085e-18, 0, 0, -8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -8.673617e-19, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.002231383, 0.001717253, 0.001620685, 0.0015974, 0.001558135, 0.001462416, 
    0.001304487, 0.001089175, 0.0009881805, 0.0007998971, 0.000570061, 
    8.785608e-05, -0.0004895027, -0.001168272, -0.001649519, -0.002135741, 
    -0.00260159, -0.002320186, -0.002122517, -0.002042739, -0.002256301, 
    -0.002752124, -0.003332893, -0.004480902, -0.008071853, -0.01055839, 
    -0.01296773, 1.734723e-18, 8.673617e-19, 8.673617e-19, 8.673617e-19, 0, 
    -2.602085e-18, 0, 0, -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, 
    -8.673617e-19, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18,
  0.003208496, 0.002588471, 0.002555653, 0.002625219, 0.002641107, 
    0.002587388, 0.002444879, 0.002223433, 0.002103947, 0.001856382, 
    0.001497013, 0.0008514259, 9.481997e-05, -0.0007777613, -0.001411841, 
    -0.002036625, -0.002632038, -0.002379652, -0.00224319, -0.002253495, 
    -0.002737245, -0.003323366, -0.004182424, -0.006750575, -0.009714451, 
    -0.0116891, -0.01430304, 1.734723e-18, 8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -2.602085e-18, 0, 0, -8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -8.673617e-19, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.004766233, 0.004033457, 0.003924808, 0.003934833, 0.004010188, 
    0.004017084, 0.003903602, 0.003684052, 0.00354442, 0.003209097, 
    0.002697755, 0.001905911, 0.0009692768, -0.0001192484, -0.001109538, 
    -0.001999615, -0.002751903, -0.002730132, -0.002721742, -0.002770122, 
    -0.003478486, -0.004748261, -0.005461288, -0.008157383, -0.01169798, 
    -0.01278353, -0.0153251, 1.734723e-18, 8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -2.602085e-18, 0, 0, -8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -8.673617e-19, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.006586552, 0.005752615, 0.005725742, 0.005794666, 0.005791214, 
    0.005811342, 0.005730339, 0.005517283, 0.00534617, 0.004870344, 
    0.004103633, 0.003133142, 0.001971298, 0.0006052646, -0.001051069, 
    -0.002381838, -0.003319368, -0.003795015, -0.003975259, -0.003945874, 
    -0.005134926, -0.006582864, -0.00659153, -0.01027504, -0.01293342, 
    -0.01400537, -0.01352196, 1.734723e-18, 8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -2.602085e-18, 0, 0, -8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -8.673617e-19, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.008633406, 0.007697643, 0.007757423, 0.007913687, 0.007965744, 
    0.008123433, 0.008061406, 0.007793605, 0.007508815, 0.006806816, 
    0.005652702, 0.004494547, 0.0030807, 0.001389171, -0.001226486, 
    -0.003183647, -0.004388244, -0.005640329, -0.006012441, -0.005599465, 
    -0.007316356, -0.008444028, -0.008017086, -0.01201829, -0.01417199, 
    -0.0139047, -0.01206139, 1.734723e-18, 8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -2.602085e-18, 0, 0, -8.673617e-19, 8.673617e-19, 
    8.673617e-19, 0, -8.673617e-19, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18,
  0.01086282, 0.009828099, 0.009984443, 0.01022506, 0.01032589, 0.01067664, 
    0.01075657, 0.010584, 0.01022389, 0.009163, 0.007412568, 0.006071981, 
    0.004386617, 0.002330512, -0.001423546, -0.004144398, -0.005740343, 
    -0.007930553, -0.008434178, -0.007315984, -0.0092641, -0.01028544, 
    -0.009873249, -0.01323392, -0.01525981, -0.01190971, -0.008459027, 
    1.734723e-18, 8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -2.602085e-18, 
    0, 0, -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -8.673617e-19, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18,
  0.01322623, 0.01209097, 0.01227868, 0.01251553, 0.01260978, 0.01315519, 
    0.01339615, 0.01335436, 0.01293775, 0.01157947, 0.009272804, 0.007738994, 
    0.005759692, 0.003321366, -0.001408633, -0.00475145, -0.006677908, 
    -0.009582207, -0.01026178, -0.008912238, -0.01127583, -0.01230159, 
    -0.0113752, -0.01405884, -0.01332307, -0.01002285, -0.004008415, 
    1.734723e-18, 8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -2.602085e-18, 
    0, 0, -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -8.673617e-19, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18,
  0.01493266, 0.01367481, 0.01357636, 0.01344964, 0.01332436, 0.01382942, 
    0.01405116, 0.01400025, 0.01359595, 0.01212949, 0.009432256, 0.007765642, 
    0.005581478, 0.002875935, -0.002262801, -0.005814572, -0.007804323, 
    -0.01094001, -0.01194366, -0.01089343, -0.01332483, -0.01388795, 
    -0.01147532, -0.01256442, -0.01138569, -0.005739278, -0.0004541221, 
    1.734723e-18, 8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -2.602085e-18, 
    0, 0, -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -8.673617e-19, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18,
  0.01435783, 0.01294075, 0.01269243, 0.01233148, 0.01187868, 0.01225575, 
    0.01225617, 0.01184392, 0.01110531, 0.009473911, 0.006935346, 
    0.005290614, 0.003492943, 0.001197792, -0.003451834, -0.007108262, 
    -0.009681559, -0.01300822, -0.01380179, -0.01209396, -0.01411556, 
    -0.01417295, -0.009519524, -0.01008835, -0.007082656, -0.002334345, 
    0.002409544, 1.734723e-18, 8.673617e-19, 8.673617e-19, 8.673617e-19, 0, 
    -2.602085e-18, 0, 0, -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, 
    -8.673617e-19, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18,
  0.01500691, 0.01361977, 0.01458739, 0.01536914, 0.01549227, 0.01618991, 
    0.01649099, 0.01644643, 0.01583415, 0.01443072, 0.01231792, 0.01096243, 
    0.008944365, 0.00624883, 0.001263245, -0.002800374, -0.005880474, 
    -0.01032474, -0.01201672, -0.01097807, -0.01323056, -0.01125193, 
    -0.006264102, -0.005268745, -0.00299966, 0.0004064999, 0.003226432, 
    1.734723e-18, 8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -2.602085e-18, 
    0, 0, -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -8.673617e-19, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18,
  0.02157488, 0.02025939, 0.02153402, 0.0224119, 0.02236979, 0.02305521, 
    0.02334202, 0.02327902, 0.02262836, 0.02136482, 0.01958451, 0.01821643, 
    0.01621024, 0.01357534, 0.008272826, 0.003954748, 0.0006824987, 
    -0.004732701, -0.006942522, -0.005777734, -0.008420462, -0.006582231, 
    0.0002074631, -0.0003475662, 0.0003091274, 0.001167735, 0.003226432, 
    1.734723e-18, 8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -2.602085e-18, 
    0, 0, -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -8.673617e-19, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18,
  0.03098602, 0.0297223, 0.03128592, 0.03222966, 0.0319822, 0.03274052, 
    0.03305401, 0.0329761, 0.0324276, 0.03149695, 0.03029714, 0.02891356, 
    0.02694781, 0.02440435, 0.01854596, 0.0139393, 0.01065576, 0.004047906, 
    0.001338356, 0.002772226, 3.523609e-05, 0.001321273, 0.006223608, 
    0.002676297, 0.0006724431, 0.001167735, 0.003226432, 1.734723e-18, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -2.602085e-18, 0, 0, 
    -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -8.673617e-19, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18,
  0.04497231, 0.04355758, 0.04468865, 0.04465833, 0.04346661, 0.04399176, 
    0.04400197, 0.04349723, 0.0427901, 0.04195892, 0.04100368, 0.03923925, 
    0.03691877, 0.03404224, 0.02742193, 0.02256103, 0.01945955, 0.01192869, 
    0.0087241, 0.009845764, 0.005503885, 0.004615062, 0.007179296, 
    0.002676297, 0.0006724431, 0.001167735, 0.003226432, 1.734723e-18, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -2.602085e-18, 0, 0, 
    -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -8.673617e-19, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18, 
    5.20417e-18, 5.20417e-18, 5.20417e-18, 5.20417e-18 ;

 v_west =
  -0.002053349, -0.001874023, -0.00175441, -0.001997134, -0.002672717, 
    -0.003350866, -0.003727, -0.003803608, -0.004125544, -0.003854587, 
    -0.003266465, -0.002910377, -0.002717788, -0.002576548, -0.002740991, 
    -0.002422532, -0.001577531, -0.001358396, -0.001024024, -0.0006485867, 
    -0.0001815921, -0.0002251074, -0.0006975927, -0.0006425674, 
    -0.0006679801, -0.0008541886, -0.0006999351, -0.0007226765, 
    -0.0008734977, -0.0006703213, -0.0005366738, -0.0007473875, 
    -0.0009139795, -0.001141787, -0.001363133, -0.001419942, -0.001344198, 
    -0.00116813, -0.0009668108, -0.000841494, -0.0007702512, -0.0007671276, 
    -0.0006575207, -0.0005202217, -0.0004828128, -0.0004292648, 
    -0.0003778311, -0.000418978, -0.0004157454, -0.0003784097, -0.0003333698, 
    -0.0003838494, -0.0004871148, -0.0004091309,
  -0.0009936204, -0.00103249, -0.001419314, -0.00192139, -0.002602797, 
    -0.003292903, -0.003683416, -0.003776603, -0.004152802, -0.004305172, 
    -0.004231582, -0.00409421, -0.003869103, -0.003557478, -0.003071493, 
    -0.002437913, -0.001627909, -0.001422252, -0.001346798, -0.001469014, 
    -0.001023773, -0.0009056919, -0.00110972, -0.001033878, -0.001081232, 
    -0.001255337, -0.0009348248, -0.0008280439, -0.0009326728, -0.0008788148, 
    -0.001092318, -0.001449868, -0.001535855, -0.001635761, -0.001752503, 
    -0.001780557, -0.001773544, -0.00172817, -0.001656839, -0.001550093, 
    -0.001410272, -0.001427105, -0.001377226, -0.001262702, -0.001256553, 
    -0.001159609, -0.0009720937, -0.0009347546, -0.0008862521, -0.0008219389, 
    -0.0007588322, -0.0007339813, -0.0007287709, -0.0007257851,
  -0.0009881345, -0.001027194, -0.001389176, -0.001902448, -0.002568727, 
    -0.003250935, -0.003644431, -0.003751604, -0.004123044, -0.004276602, 
    -0.004209354, -0.004078384, -0.003856024, -0.003546601, -0.003088379, 
    -0.002470571, -0.001692789, -0.001490292, -0.001434623, -0.001526658, 
    -0.001098108, -0.0009827273, -0.0011738, -0.001107522, -0.001159485, 
    -0.001333217, -0.00104743, -0.000968023, -0.001133011, -0.00113807, 
    -0.001211092, -0.001416294, -0.00149989, -0.001597442, -0.00171162, 
    -0.001747391, -0.001750902, -0.001718878, -0.001664905, -0.001574314, 
    -0.001449248, -0.001466182, -0.001416578, -0.001302325, -0.001286535, 
    -0.001185801, -0.001000328, -0.001004566, -0.0009734288, -0.0009026651, 
    -0.0009102552, -0.0009096924, -0.0008666518, -0.0009088299,
  -0.0009793601, -0.001018364, -0.001383555, -0.001890683, -0.002540746, 
    -0.003209501, -0.003601124, -0.00372029, -0.004089337, -0.004244771, 
    -0.004177459, -0.004051209, -0.003834495, -0.003528668, -0.00308909, 
    -0.002496823, -0.001751455, -0.001551147, -0.001491446, -0.001572836, 
    -0.001163033, -0.001050772, -0.001228742, -0.001171811, -0.001228652, 
    -0.00140251, -0.001148669, -0.001082868, -0.001193363, -0.001127597, 
    -0.001196709, -0.001377236, -0.001452847, -0.001547716, -0.001662924, 
    -0.001713071, -0.001732336, -0.001716516, -0.001682901, -0.001610469, 
    -0.00150193, -0.001523351, -0.001476016, -0.00136302, -0.001339557, 
    -0.001237255, -0.001057799, -0.001062763, -0.001026128, -0.000949708, 
    -0.0009522158, -0.0009286713, -0.0008758684, -0.0009050265,
  -0.0009674193, -0.00100572, -0.001370369, -0.001866718, -0.002495689, 
    -0.003147065, -0.003534602, -0.003662624, -0.004020893, -0.004175738, 
    -0.004122703, -0.004014094, -0.00381012, -0.00350884, -0.003085958, 
    -0.002517476, -0.001803011, -0.001604561, -0.00154078, -0.001612118, 
    -0.001214338, -0.001094939, -0.001251022, -0.00119456, -0.001243608, 
    -0.001392883, -0.00114085, -0.001073325, -0.00117753, -0.001100665, 
    -0.001141557, -0.001313057, -0.001398196, -0.001500204, -0.001620079, 
    -0.001683323, -0.001716252, -0.001714982, -0.001700565, -0.001645089, 
    -0.001551058, -0.001577554, -0.001534991, -0.001426232, -0.001398563, 
    -0.001296083, -0.001120347, -0.001112761, -0.001067562, -0.0009864267, 
    -0.0009783235, -0.0009451222, -0.0008838573, -0.000901702,
  -0.0009430419, -0.0009810082, -0.001347644, -0.001837105, -0.002448591, 
    -0.003083196, -0.003464396, -0.003600325, -0.003956825, -0.004109266, 
    -0.004053272, -0.003944885, -0.003741161, -0.003442945, -0.003038485, 
    -0.002494484, -0.001810991, -0.001614, -0.001542908, -0.001595452, 
    -0.001208385, -0.00108745, -0.00122611, -0.001173551, -0.001218684, 
    -0.001356602, -0.001125315, -0.001057367, -0.001125744, -0.001040612, 
    -0.001088216, -0.001256697, -0.001343072, -0.001435239, -0.001550603, 
    -0.001625692, -0.001676119, -0.001695062, -0.001704113, -0.001667578, 
    -0.001589465, -0.001624439, -0.001588879, -0.001485213, -0.001454508, 
    -0.001352265, -0.001180664, -0.001163894, -0.00111103, -0.00102355, 
    -0.001005721, -0.0009625822, -0.0008890388, -0.0008971078,
  -0.0009055574, -0.0009418062, -0.001304057, -0.001779473, -0.002367308, 
    -0.002981525, -0.003354868, -0.003494915, -0.003837929, -0.003995667, 
    -0.003960864, -0.003875985, -0.003679461, -0.003381435, -0.002991119, 
    -0.002467457, -0.001810493, -0.001613132, -0.001535949, -0.001576837, 
    -0.001203059, -0.001074025, -0.001186797, -0.001130589, -0.001164056, 
    -0.001277179, -0.001050381, -0.0009835291, -0.001056485, -0.0009868797, 
    -0.001013786, -0.001155752, -0.001242644, -0.00134599, -0.001469298, 
    -0.001560246, -0.001627153, -0.001663665, -0.001694769, -0.00167863, 
    -0.001618982, -0.001665616, -0.001640157, -0.001544868, -0.00151475, 
    -0.001414084, -0.001244899, -0.001218952, -0.001157457, -0.00106179, 
    -0.001033856, -0.0009793567, -0.0008935464, -0.0008929326,
  -0.0008711594, -0.0009058322, -0.00126406, -0.001726586, -0.002292718, 
    -0.002888226, -0.00325436, -0.003398185, -0.003728824, -0.003877336, 
    -0.003836947, -0.003748994, -0.003559373, -0.003268244, -0.002895602, 
    -0.002394635, -0.001766029, -0.001569752, -0.00148402, -0.001503488, 
    -0.001129355, -0.0009931189, -0.00108995, -0.001037426, -0.001068656, 
    -0.001174299, -0.0009699694, -0.0009157715, -0.0009929275, -0.0008852822, 
    -0.0009071119, -0.001050601, -0.001150483, -0.001264088, -0.001394685, 
    -0.001500187, -0.001582218, -0.001634852, -0.001686194, -0.001688773, 
    -0.001646069, -0.001703404, -0.001687215, -0.001599613, -0.001570034, 
    -0.001470814, -0.001303847, -0.001269477, -0.001200062, -0.001096882, 
    -0.001059675, -0.0009947504, -0.0008976831, -0.0008880975,
  -0.0007742649, -0.0008101587, -0.001172227, -0.001629136, -0.002176935, 
    -0.00275196, -0.003106734, -0.003254099, -0.003583907, -0.003749969, 
    -0.003719622, -0.003628758, -0.003437165, -0.00314499, -0.002785433, 
    -0.002303498, -0.001699825, -0.001501916, -0.001409045, -0.001416234, 
    -0.001054344, -0.0009165169, -0.0009982563, -0.0009492195, -0.0009783314, 
    -0.001076892, -0.0008763671, -0.0008130232, -0.000858687, -0.0007728627, 
    -0.0008061104, -0.0009510408, -0.001060225, -0.001171795, -0.001302889, 
    -0.001423191, -0.001524284, -0.001597997, -0.001672297, -0.001694722, 
    -0.001669523, -0.001739283, -0.00173251, -0.001651618, -0.001621491, 
    -0.001522108, -0.001353857, -0.001305461, -0.001222205, -0.001106472, 
    -0.001052756, -0.0009602867, -0.0008269171, -0.0008056353,
  -0.0006668865, -0.0007018593, -0.001057585, -0.001498972, -0.002022353, 
    -0.002576054, -0.002921389, -0.003070273, -0.003385498, -0.00354019, 
    -0.003523123, -0.003460474, -0.003287568, -0.003004499, -0.002663218, 
    -0.002204006, -0.001628396, -0.001431771, -0.001329598, -0.001313086, 
    -0.0009471183, -0.00079303, -0.0008482253, -0.0007945186, -0.0008133283, 
    -0.0008908692, -0.0007147547, -0.0006697674, -0.0007270286, 
    -0.0006627021, -0.0006865216, -0.0008152856, -0.0009303386, -0.001056364, 
    -0.00119738, -0.00133692, -0.001458081, -0.00155328, -0.001651142, 
    -0.001695304, -0.001689709, -0.001774579, -0.001778271, -0.001703024, 
    -0.001668952, -0.00156396, -0.001388407, -0.001321439, -0.001219744, 
    -0.001085535, -0.001014623, -0.0009036157, -0.0007505189, -0.0007213026,
  -0.0005565076, -0.0005922705, -0.0009415788, -0.001367258, -0.001865931, 
    -0.002398053, -0.002733837, -0.002884258, -0.003184726, -0.003327914, 
    -0.003303477, -0.003235409, -0.00305947, -0.002775747, -0.002449077, 
    -0.00201047, -0.00146134, -0.001262222, -0.001151482, -0.001121021, 
    -0.0007683553, -0.0006136735, -0.0006545841, -0.0006052104, 
    -0.0006244632, -0.0006996432, -0.0005512181, -0.0005248059, 
    -0.0005836949, -0.0005019162, -0.0005303629, -0.0006649547, 
    -0.0007989064, -0.0009395594, -0.001090614, -0.001249623, -0.00139109, 
    -0.001508031, -0.001629735, -0.001695892, -0.001710135, -0.001810294, 
    -0.001824575, -0.001755041, -0.001716978, -0.00160631, -0.001423368, 
    -0.001337607, -0.001217254, -0.001064349, -0.0009760374, -0.0008462703, 
    -0.0006732116, -0.0006359664,
  -0.0003488836, -0.0003904197, -0.0007428012, -0.001160655, -0.001638369, 
    -0.002148912, -0.002473517, -0.00262637, -0.002920838, -0.003069983, 
    -0.00306012, -0.003002225, -0.002823144, -0.002538744, -0.002227211, 
    -0.001809952, -0.001288257, -0.001086557, -0.0009669411, -0.0009220273, 
    -0.0005831437, -0.0004278471, -0.0004499295, -0.000398531, -0.0004108098, 
    -0.0004710905, -0.0003369146, -0.0003152427, -0.0003728603, 
    -0.0003218862, -0.0003685735, -0.0005092034, -0.0006633007, 
    -0.0008211961, -0.000983365, -0.00116538, -0.001329827, -0.001469956, 
    -0.001614745, -0.001702648, -0.001736563, -0.001852208, -0.001874878, 
    -0.001808052, -0.001762706, -0.001642438, -0.001444408, -0.001327133, 
    -0.001175837, -0.0009943304, -0.0008740327, -0.0006934038, -0.0004554283, 
    -0.0003978741,
  -0.0001310525, -0.0001780667, -0.000524713, -0.0009266633, -0.001378877, 
    -0.001867758, -0.002183151, -0.0023378, -0.002617798, -0.00275588, 
    -0.002739752, -0.002679958, -0.002510833, -0.002233059, -0.001941158, 
    -0.001548112, -0.001055684, -0.0008510428, -0.0007179977, -0.0006470471, 
    -0.0003086216, -0.000140098, -0.0001411552, -9.14469e-05, -0.0001049771, 
    -0.000167665, -6.753687e-05, -7.233808e-05, -0.0001522332, -0.0001341501, 
    -0.0002014324, -0.0003496735, -0.0005288948, -0.000703776, -0.0008753213, 
    -0.001083372, -0.001274577, -0.001442875, -0.001613102, -0.001722715, 
    -0.001774318, -0.001905961, -0.001933629, -0.001860446, -0.001793171, 
    -0.001645661, -0.001415364, -0.001252297, -0.001055483, -0.0008283462, 
    -0.000669473, -0.0004492381, -0.0001703221, -9.910145e-05,
  1.012876e-05, -4.904123e-05, -0.0003820058, -0.0007601236, -0.001182833, 
    -0.001651909, -0.001961417, -0.002116117, -0.002370706, -0.002471626, 
    -0.002412861, -0.002341275, -0.002170348, -0.001894274, -0.001620261, 
    -0.001250095, -0.0007853279, -0.0005747126, -0.0004274749, -0.0003352331, 
    -7.668339e-06, 0.0001640085, 0.0001800806, 0.0002280302, 0.0002126857, 
    0.0001459146, 0.0002106393, 0.0001785207, 7.35171e-05, 5.758827e-05, 
    -2.920837e-05, -0.0001843766, -0.0003890673, -0.0005816196, 
    -0.0007629197, -0.0009980561, -0.0012171, -0.001414701, -0.001611393, 
    -0.001743592, -0.001813597, -0.001961883, -0.00199475, -0.001914953, 
    -0.001824865, -0.001649014, -0.001385148, -0.001174441, -0.0009302745, 
    -0.0006556668, -0.0004566624, -0.000195224, 0.0001524171, 0.0002478032,
  9.888375e-05, 1.938206e-05, -0.0003132843, -0.0006800938, -0.001080562, 
    -0.001531377, -0.001832249, -0.001987291, -0.002232128, -0.002328082, 
    -0.002269958, -0.002168968, -0.001975222, -0.001689152, -0.001423666, 
    -0.001065745, -0.0006160517, -0.0003869639, -0.0002151404, -9.387276e-05, 
    0.0002308844, 0.0004151965, 0.0004586993, 0.000519493, 0.0005136349, 
    0.0004507592, 0.0004879286, 0.0004314288, 0.000301957, 0.0002487951, 
    9.845469e-05, -8.776944e-05, -0.0003390995, -0.0005664642, -0.0007650439, 
    -0.001039408, -0.001292464, -0.00152124, -0.001736246, -0.001885958, 
    -0.001970984, -0.002133047, -0.002156593, -0.002048841, -0.001910145, 
    -0.001678279, -0.0013493, -0.001053004, -0.0007221529, -0.0003617853, 
    -8.554732e-05, 0.0002702701, 0.0007023027, 0.0008293592,
  -0.0003142593, -0.0004108969, -0.0007006598, -0.001017816, -0.001374988, 
    -0.001807891, -0.002105495, -0.002250101, -0.002445429, -0.002451217, 
    -0.002280384, -0.00207316, -0.001831759, -0.001545505, -0.001291674, 
    -0.0009460063, -0.0005090627, -0.0002584476, -5.374603e-05, 0.0001107074, 
    0.0004469846, 0.0006304802, 0.0006910418, 0.0007606428, 0.0007586767, 
    0.0006860407, 0.0006819731, 0.0005864772, 0.0004022167, 0.0002797622, 
    0.0001239922, -6.065306e-05, -0.0003346857, -0.0005744095, -0.0007757543, 
    -0.001084293, -0.00137334, -0.001640384, -0.001880249, -0.002048326, 
    -0.002145127, -0.002321438, -0.002338736, -0.002203122, -0.002011434, 
    -0.001715682, -0.001312535, -0.0009246582, -0.000503301, -5.271905e-05, 
    0.0002992584, 0.0007327293, 0.001255317, 0.001419443,
  -0.0009943668, -0.001120651, -0.001409906, -0.001714775, -0.002045679, 
    -0.002456895, -0.002735672, -0.002867399, -0.003057286, -0.003067803, 
    -0.002909613, -0.00270365, -0.002434942, -0.002101986, -0.0018217, 
    -0.001448693, -0.0009811756, -0.0006651943, -0.0003927406, -0.0001632845, 
    0.0002037162, 0.0004560771, 0.000594528, 0.0007219188, 0.0007669801, 
    0.0007304525, 0.0007281139, 0.000631951, 0.0004441627, 0.0002238933, 
    -4.656177e-06, -0.0002250873, -0.0005514381, -0.0008291161, -0.001047078, 
    -0.00141182, -0.001751038, -0.002065138, -0.002319541, -0.002503115, 
    -0.002614491, -0.002805013, -0.002798438, -0.002608038, -0.002329901, 
    -0.001937477, -0.001428112, -0.0009092002, -0.0003559777, 0.0002253315, 
    0.0006894897, 0.001245436, 0.00189414, 0.002111342,
  -0.002950786, -0.003083209, -0.003297942, -0.003526236, -0.003793531, 
    -0.004182623, -0.004445854, -0.004543016, -0.004675185, -0.004572792, 
    -0.004267874, -0.003910927, -0.003531806, -0.003126669, -0.002796434, 
    -0.002372187, -0.001848637, -0.001440493, -0.001078557, -0.000769648, 
    -0.000359292, -4.614265e-05, 0.0001728843, 0.0003690743, 0.0004721075, 
    0.0004725278, 0.0004635043, 0.0003571068, 0.0001346223, -6.9527e-05, 
    -0.0002774342, -0.0004940745, -0.0008764098, -0.001194874, -0.001428469, 
    -0.001857712, -0.002254263, -0.002621299, -0.002883137, -0.003079179, 
    -0.003205331, -0.003406948, -0.00337055, -0.003117853, -0.002742697, 
    -0.002244692, -0.001622524, -0.0009630977, -0.0002715028, 0.0004438413, 
    0.001023231, 0.001698362, 0.002474484, 0.002745586,
  -0.005432389, -0.005564137, -0.005709537, -0.005867993, -0.006077835, 
    -0.006455366, -0.006707133, -0.006769469, -0.006855841, -0.006646795, 
    -0.006195065, -0.005680127, -0.005252803, -0.004807665, -0.004428135, 
    -0.003942536, -0.003346683, -0.002820608, -0.002320196, -0.001850852, 
    -0.001308338, -0.0008745015, -0.0005474777, -0.0002591128, -7.510863e-05, 
    -1.443276e-05, -1.708732e-05, -0.0001212357, -0.0003654044, 
    -0.0006442326, -0.0009067919, -0.00113435, -0.001515288, -0.001817799, 
    -0.002025254, -0.002522532, -0.002997849, -0.003453716, -0.003731834, 
    -0.003940284, -0.00407582, -0.004285246, -0.004221863, -0.003902875, 
    -0.00340852, -0.002779309, -0.002014206, -0.001171074, -0.000315615, 
    0.0005455039, 0.001257571, 0.002067847, 0.002980488, 0.003305258,
  -0.008399032, -0.008528712, -0.008630881, -0.008770955, -0.008960012, 
    -0.009340224, -0.009573524, -0.009610323, -0.009736783, -0.00958334, 
    -0.009191068, -0.008702184, -0.008180286, -0.007622022, -0.00712284, 
    -0.006512814, -0.005784924, -0.00506519, -0.004371717, -0.003715301, 
    -0.003025733, -0.002413898, -0.001875131, -0.001425185, -0.001088393, 
    -0.0008795241, -0.000814808, -0.0008487252, -0.001050298, -0.001387989, 
    -0.001704326, -0.001957099, -0.002397144, -0.002717733, -0.00288814, 
    -0.003500864, -0.004084267, -0.004642331, -0.004876933, -0.005063201, 
    -0.005194301, -0.005374951, -0.005243053, -0.004820086, -0.00415129, 
    -0.003358727, -0.002440229, -0.001373946, -0.0003386805, 0.0006571004, 
    0.001505717, 0.002451143, 0.003495607, 0.003855904,
  -0.01176244, -0.01191217, -0.01206375, -0.01222779, -0.01243878, -0.012894, 
    -0.01317115, -0.01321115, -0.01338287, -0.01321098, -0.01274651, 
    -0.01216067, -0.01153185, -0.01085824, -0.01021458, -0.009457988, 
    -0.008579452, -0.007632492, -0.006711862, -0.005830413, -0.004951842, 
    -0.00413329, -0.003369014, -0.002758723, -0.002264295, -0.001902862, 
    -0.001821158, -0.001826958, -0.001958039, -0.002287326, -0.002623852, 
    -0.002883501, -0.003394017, -0.003716446, -0.003801688, -0.004556614, 
    -0.005269459, -0.005943663, -0.006090571, -0.006219163, -0.006318852, 
    -0.006440495, -0.006219745, -0.005677199, -0.004793344, -0.003812819, 
    -0.002729289, -0.001404922, -0.0001830758, 0.0009263614, 0.001904084, 
    0.002979332, 0.004145813, 0.00452162,
  -0.01458343, -0.01477674, -0.01502575, -0.01528286, -0.01557972, 
    -0.01615361, -0.016503, -0.01657323, -0.0168428, -0.01672683, 
    -0.01627454, -0.01567286, -0.01498554, -0.01421258, -0.01341389, 
    -0.01249972, -0.01146137, -0.01026655, -0.009091006, -0.007943586, 
    -0.006819834, -0.005738374, -0.004695273, -0.003912972, -0.003246101, 
    -0.002704581, -0.002627847, -0.002624138, -0.002724005, -0.003170533, 
    -0.00355123, -0.003802993, -0.004405955, -0.004707173, -0.004641237, 
    -0.005566957, -0.006435182, -0.007244709, -0.007260634, -0.007297414, 
    -0.007343736, -0.007395242, -0.007078101, -0.006408593, -0.005264645, 
    -0.00406812, -0.002809913, -0.001199846, 0.000214303, 0.001421647, 
    0.002514283, 0.003701474, 0.004971394, 0.005348008,
  -0.01653155, -0.01679101, -0.01719534, -0.01759966, -0.01802574, 
    -0.01874116, -0.01917525, -0.0192904, -0.0196949, -0.01970121, 
    -0.01934451, -0.01880707, -0.01811243, -0.0172619, -0.01630927, 
    -0.01523395, -0.01403017, -0.01258027, -0.01113231, -0.009684117, 
    -0.00825064, -0.006842487, -0.005461787, -0.004505388, -0.003666337, 
    -0.002937387, -0.002911674, -0.002947643, -0.003052409, -0.003649411, 
    -0.004127845, -0.004409375, -0.005211526, -0.005505195, -0.005229906, 
    -0.006360029, -0.007410086, -0.008373179, -0.008222572, -0.008152965, 
    -0.008154741, -0.008180246, -0.00780192, -0.007034633, -0.005605881, 
    -0.004173167, -0.002730349, -0.0008216198, 0.0007928149, 0.002101201, 
    0.003289889, 0.004559204, 0.005905071, 0.006280207,
  -0.01756562, -0.01789854, -0.01847284, -0.01904487, -0.01962607, 
    -0.02050097, -0.02103301, -0.02119926, -0.02173845, -0.02186503, 
    -0.02160063, -0.02111988, -0.02041306, -0.01948212, -0.01837891, 
    -0.01713256, -0.01574134, -0.01403441, -0.01231171, -0.0105587, 
    -0.00876653, -0.006983401, -0.00522186, -0.004110817, -0.003134552, 
    -0.002269207, -0.002394821, -0.002586575, -0.002831804, -0.003700451, 
    -0.004344735, -0.0046607, -0.005762434, -0.006064955, -0.005499082, 
    -0.006868859, -0.008135121, -0.009286964, -0.008952395, -0.008805107, 
    -0.008837716, -0.008979029, -0.00866926, -0.007924275, -0.00624953, 
    -0.004585062, -0.002926316, -0.0006920599, 0.00114821, 0.002587353, 
    0.003862836, 0.005219001, 0.006660474, 0.007066691,
  -0.01779038, -0.01819261, -0.01890526, -0.0196622, -0.02046197, 
    -0.02151638, -0.0221641, -0.02239332, -0.02307528, -0.02331231, 
    -0.02312515, -0.02267983, -0.0219494, -0.02092792, -0.01970074, 
    -0.01825022, -0.01657774, -0.01458042, -0.0125439, -0.01044925, 
    -0.008183704, -0.005941875, -0.003744046, -0.002493764, -0.001436781, 
    -0.0005402789, -0.0009414793, -0.001438132, -0.002003982, -0.003259524, 
    -0.004134453, -0.004530663, -0.006008739, -0.006311888, -0.005454332, 
    -0.00708893, -0.008605896, -0.009989624, -0.009509807, -0.009328452, 
    -0.009445372, -0.009733299, -0.009531198, -0.008846833, -0.006975878, 
    -0.005155093, -0.003397048, -0.0009254455, 0.001061125, 0.002569569, 
    0.003870943, 0.005220232, 0.006667488, 0.00713217,
  -0.01734996, -0.01792934, -0.01888408, -0.01986201, -0.02087567, 
    -0.02217185, -0.02296998, -0.02325796, -0.02404376, -0.02430141, 
    -0.02406322, -0.0235443, -0.02273424, -0.02162111, -0.02027079, 
    -0.0185956, -0.01659484, -0.01434586, -0.01200821, -0.009555501, 
    -0.006700373, -0.003958843, -0.001355975, 1.698876e-05, 0.001088462, 
    0.001887745, 0.001137066, 0.0002539162, -0.0007167619, -0.002326995, 
    -0.003385663, -0.004196223, -0.006390012, -0.007179155, -0.006421099, 
    -0.008193101, -0.009778433, -0.01123653, -0.01052541, -0.01036255, 
    -0.01072208, -0.0112697, -0.01122912, -0.01066772, -0.008851524, 
    -0.007160712, -0.005649806, -0.003615229, -0.001954307, -0.0006635745, 
    0.0004431276, 0.00154245, 0.002765837, 0.003271171,
  -0.01772479, -0.01851436, -0.01978852, -0.02112143, -0.02252645, 
    -0.02415112, -0.02535792, -0.02611058, -0.02722327, -0.02762105, 
    -0.02731372, -0.02660239, -0.02555004, -0.02419424, -0.0228111, 
    -0.0208641, -0.0183575, -0.01575187, -0.01308202, -0.01037116, 
    -0.00736184, -0.004680705, -0.002339787, -0.001097851, -0.0003842048, 
    -0.0002986453, -0.001771411, -0.003396015, -0.005403629, -0.008506973, 
    -0.0105921, -0.01146683, -0.01345141, -0.01383264, -0.01244226, 
    -0.01380028, -0.01513902, -0.01650952, -0.01548083, -0.0152829, 
    -0.01589826, -0.0168527, -0.01728112, -0.01724755, -0.01566073, 
    -0.01417414, -0.01282545, -0.01106192, -0.009555442, -0.00832051, 
    -0.007366062, -0.006220855, -0.004805113, -0.004140875,
  -0.01836369, -0.01934242, -0.02102031, -0.02283597, -0.02480108, 
    -0.02684791, -0.0285145, -0.02977249, -0.03135783, -0.03230022, 
    -0.03260494, -0.03249694, -0.0319674, -0.0310329, -0.03033028, 
    -0.02873051, -0.02622497, -0.02390786, -0.02114593, -0.01799949, 
    -0.01454943, -0.01151685, -0.00888016, -0.00716392, -0.006230166, 
    -0.006139861, -0.007430251, -0.009047784, -0.01117537, -0.01442753, 
    -0.01663068, -0.01765999, -0.01991012, -0.02004953, -0.01800585, 
    -0.01900894, -0.02013334, -0.02140129, -0.02024143, -0.0201321, 
    -0.02106524, -0.02239346, -0.02322531, -0.02359837, -0.02213972, 
    -0.02063499, -0.01909604, -0.01691918, -0.01503768, -0.01347283, 
    -0.01230265, -0.01083699, -0.009053068, -0.00813977,
  -0.0194362, -0.02057746, -0.02264613, -0.02493924, -0.02746631, 
    -0.02997778, -0.03209166, -0.03378466, -0.0357841, -0.03714564, 
    -0.03788298, -0.03818371, -0.0381455, -0.03777337, -0.03761691, 
    -0.03650097, -0.03442273, -0.03271825, -0.03008461, -0.02654631, 
    -0.02215902, -0.01813618, -0.01447391, -0.01177364, -0.01018723, 
    -0.009738931, -0.0106558, -0.01228513, -0.01470873, -0.01814753, 
    -0.02043508, -0.02150012, -0.02393596, -0.02386281, -0.02122601, 
    -0.02207469, -0.02312452, -0.0243748, -0.02315438, -0.02314824, 
    -0.02436195, -0.02636216, -0.02774366, -0.02852826, -0.02690297, 
    -0.02500561, -0.02283813, -0.01964107, -0.01696004, -0.01481654, 
    -0.0136066, -0.01198806, -0.009960488, -0.008785993,
  -0.02066245, -0.02191226, -0.02431705, -0.02695487, -0.02982906, 
    -0.03259313, -0.03498669, -0.0370038, -0.03933585, -0.04108734, 
    -0.0422604, -0.04286093, -0.04314785, -0.04312178, -0.04340589, 
    -0.04253387, -0.04050617, -0.0393557, -0.0365972, -0.03223667, 
    -0.02624445, -0.02084359, -0.01603903, -0.01236246, -0.01028306, 
    -0.009803236, -0.0105871, -0.01247956, -0.015494, -0.01944774, 
    -0.0220362, -0.02323804, -0.02591396, -0.02542495, -0.021771, 
    -0.02265509, -0.02382014, -0.02526615, -0.02452672, -0.02497864, 
    -0.0266219, -0.02956969, -0.03168488, -0.03296747, -0.03096207, 
    -0.02833198, -0.02507721, -0.02018525, -0.01627066, -0.01333343, 
    -0.01225031, -0.01057858, -0.008318231, -0.006753175,
  -0.001369803, -0.001268756, -0.001189453, -0.001376109, -0.001878729, 
    -0.002287412, -0.002536214, -0.002626961, -0.002738723, -0.002509303, 
    -0.002125111, -0.001970329, -0.001896097, -0.001785068, -0.0018592, 
    -0.001593119, -0.0009668187, -0.0008816529, -0.0006716789, -0.0003976356, 
    -4.294842e-05, -7.405259e-05, -0.0004350843, -0.000417271, -0.0004647868, 
    -0.0006535689, -0.00061273, -0.0007310167, -0.0008658079, -0.0006789761, 
    -0.0005419381, -0.0007116714, -0.0008609729, -0.001114082, -0.001400293, 
    -0.001442316, -0.001341199, -0.001142753, -0.0009863115, -0.0008831235, 
    -0.0008045717, -0.0008589203, -0.0007906641, -0.0006732624, 
    -0.0006855141, -0.000654846, -0.0005830016, -0.0006632039, -0.000690048, 
    -0.0006692009, -0.0006756135, -0.0007121121, -0.0007596953, -0.0006795931,
  -0.0006358178, -0.0006852887, -0.0009616676, -0.001328646, -0.001831662, 
    -0.002246169, -0.002505544, -0.002611447, -0.002761019, -0.002786765, 
    -0.002686067, -0.002557539, -0.002398698, -0.002211073, -0.001999928, 
    -0.001605932, -0.001015481, -0.0009424792, -0.000943913, -0.00107503, 
    -0.0007345749, -0.0006586827, -0.0008418309, -0.0008424667, 
    -0.0009216272, -0.001083598, -0.0008871402, -0.0008303273, -0.000910843, 
    -0.0009278141, -0.00117731, -0.001557172, -0.001582015, -0.001671676, 
    -0.001829454, -0.001821875, -0.001775708, -0.001687677, -0.001643903, 
    -0.001531278, -0.00135239, -0.001408772, -0.001362285, -0.001213062, 
    -0.001221986, -0.001118007, -0.0009019342, -0.000938013, -0.000929129, 
    -0.0008731171, -0.0008748645, -0.0008848719, -0.0008915918, -0.0008725795,
  -0.0006509876, -0.0006997723, -0.0009580462, -0.001329557, -0.001816532, 
    -0.002220691, -0.00248104, -0.002599142, -0.002747918, -0.002777906, 
    -0.002685625, -0.002562153, -0.002404755, -0.002216357, -0.002022018, 
    -0.001646449, -0.00108883, -0.001016067, -0.001032045, -0.001137726, 
    -0.0008139773, -0.0007404462, -0.0009104527, -0.0009186972, -0.001002543, 
    -0.001166485, -0.001003917, -0.0009808418, -0.001151304, -0.001217469, 
    -0.001315358, -0.001521964, -0.001541416, -0.001624854, -0.001775294, 
    -0.001768919, -0.001728978, -0.001652421, -0.001622979, -0.001527296, 
    -0.001367743, -0.001424791, -0.001382779, -0.001241833, -0.001246125, 
    -0.00114318, -0.0009337357, -0.0009895036, -0.0009872033, -0.0009248537, 
    -0.0009673231, -0.0009907892, -0.0009748561, -0.0009881941,
  -0.0006622649, -0.0007100757, -0.0009705143, -0.001335196, -0.00180573, 
    -0.002195095, -0.002452027, -0.002580137, -0.002730599, -0.002766543, 
    -0.002679164, -0.002560826, -0.002406411, -0.002217894, -0.002035877, 
    -0.001682789, -0.001157679, -0.001084139, -0.001094883, -0.001190587, 
    -0.0008855252, -0.0008154698, -0.0009732011, -0.0009885989, -0.001077035, 
    -0.001242645, -0.001109692, -0.001108562, -0.001228101, -0.001209301, 
    -0.00130156, -0.001483474, -0.001494705, -0.001573925, -0.001721725, 
    -0.001722235, -0.001692903, -0.001629956, -0.001618054, -0.001541639, 
    -0.001403639, -0.001466499, -0.001431225, -0.001299425, -0.001300323, 
    -0.001200264, -0.001001747, -0.001053967, -0.00104453, -0.0009754224, 
    -0.001009503, -0.001014842, -0.0009876717, -0.000989028,
  -0.000670133, -0.0007165081, -0.0009759637, -0.001329821, -0.001779568, 
    -0.002150398, -0.002401272, -0.002535529, -0.002680276, -0.002720328, 
    -0.002650468, -0.002548915, -0.002404772, -0.002217729, -0.002046492, 
    -0.00171409, -0.001219643, -0.00114511, -0.001150589, -0.001236707, 
    -0.0009434292, -0.000866723, -0.001003764, -0.001017941, -0.001098824, 
    -0.00124244, -0.001108787, -0.001103693, -0.00121553, -0.001186675, 
    -0.001253478, -0.001425649, -0.00144405, -0.001526972, -0.001674963, 
    -0.001681769, -0.001661677, -0.001611196, -0.001616221, -0.00155787, 
    -0.001438849, -0.00150816, -0.001482188, -0.001362424, -0.001363317, 
    -0.001267172, -0.0010763, -0.001114897, -0.001095641, -0.001020366, 
    -0.001041725, -0.001035691, -0.0009987804, -0.0009898078,
  -0.0006640318, -0.0007094292, -0.0009703443, -0.001317106, -0.001749563, 
    -0.002102671, -0.00234544, -0.002484874, -0.002632226, -0.002674609, 
    -0.002607082, -0.00250803, -0.002364202, -0.002177501, -0.002017209, 
    -0.00170477, -0.001239643, -0.001163453, -0.001160527, -0.001228895, 
    -0.0009457746, -0.0008678237, -0.0009887897, -0.001004871, -0.001081778, 
    -0.001215818, -0.001099592, -0.001092492, -0.001170944, -0.001135109, 
    -0.001207102, -0.00137487, -0.00139312, -0.001464519, -0.001604599, 
    -0.001615692, -0.001607986, -0.00157543, -0.001602593, -0.001564492, 
    -0.00146548, -0.001545185, -0.001530401, -0.001422469, -0.001423859, 
    -0.001331437, -0.001148143, -0.001177033, -0.001149004, -0.001065637, 
    -0.001075716, -0.001058483, -0.001007921, -0.0009917429,
  -0.0006438963, -0.000687112, -0.0009436091, -0.001276678, -0.001686177, 
    -0.002018223, -0.002250869, -0.002390639, -0.002529298, -0.002581833, 
    -0.002539821, -0.002465045, -0.002327902, -0.002139398, -0.001986788, 
    -0.001690653, -0.00125049, -0.001171115, -0.001161033, -0.001218408, 
    -0.000947873, -0.0008623222, -0.0009592361, -0.0009701624, -0.001036066, 
    -0.001148886, -0.001035034, -0.001028046, -0.00111075, -0.00108897, 
    -0.001141842, -0.001284309, -0.001301354, -0.001380222, -0.001524033, 
    -0.001543114, -0.001546758, -0.001529327, -0.001577823, -0.001561666, 
    -0.001484912, -0.00157879, -0.001578589, -0.001485557, -0.001490923, 
    -0.001403015, -0.001224569, -0.001243746, -0.001205772, -0.001112117, 
    -0.001110742, -0.001080591, -0.001016057, -0.0009934527,
  -0.0006254187, -0.0006666324, -0.0009190753, -0.001239578, -0.00162801, 
    -0.001940729, -0.002164085, -0.002304164, -0.002434847, -0.002483196, 
    -0.00244136, -0.002367077, -0.002237325, -0.002053809, -0.001911334, 
    -0.001632769, -0.001218209, -0.001137045, -0.001117515, -0.001154672, 
    -0.0008831032, -0.0007911069, -0.0008744432, -0.0008871303, -0.000951463, 
    -0.001059925, -0.0009650417, -0.0009689073, -0.001055512, -0.001000199, 
    -0.001047807, -0.001190023, -0.001217143, -0.001302864, -0.001450098, 
    -0.00147651, -0.001490569, -0.001487018, -0.001555091, -0.001559073, 
    -0.001502745, -0.00160963, -0.001622811, -0.001543452, -0.001552467, 
    -0.0014687, -0.001294704, -0.001304968, -0.001257867, -0.001154772, 
    -0.001142886, -0.001100879, -0.001023523, -0.0009940324,
  -0.0005428722, -0.00058506, -0.0008417467, -0.001157251, -0.001528198, 
    -0.00181999, -0.002029633, -0.002169, -0.002303359, -0.002374459, 
    -0.002348137, -0.002274321, -0.002143887, -0.001958424, -0.001821871, 
    -0.001557205, -0.00116451, -0.001078955, -0.001051387, -0.001077202, 
    -0.0008167108, -0.0007236802, -0.0007941612, -0.0008085154, 
    -0.0008713609, -0.0009756976, -0.000882815, -0.0008779468, -0.0009375032, 
    -0.0009017431, -0.0009587718, -0.001100752, -0.001134779, -0.001216485, 
    -0.001361271, -0.001393901, -0.001421184, -0.001436051, -0.001527745, 
    -0.001553539, -0.001518302, -0.001640821, -0.001667397, -0.001599979, 
    -0.00161111, -0.00152948, -0.001356074, -0.001351972, -0.001289636, 
    -0.001171578, -0.001142169, -0.001071333, -0.0009560029, -0.0009172597,
  -0.0004494184, -0.0004904441, -0.0007412562, -0.001042035, -0.00138965, 
    -0.001659797, -0.001857334, -0.001993278, -0.002117506, -0.002182841, 
    -0.002176395, -0.00213473, -0.002024083, -0.001846625, -0.001720822, 
    -0.001473442, -0.001105495, -0.001018448, -0.0009807664, -0.0009841814, 
    -0.0007186703, -0.0006104778, -0.000658016, -0.0006662944, -0.0007208996, 
    -0.0008105993, -0.0007383929, -0.0007502426, -0.0008217638, 
    -0.0008052654, -0.0008542427, -0.0009806529, -0.001017713, -0.001109576, 
    -0.001260382, -0.001302442, -0.001343269, -0.001376306, -0.00149335, 
    -0.001543693, -0.001531852, -0.001674085, -0.001716139, -0.001659825, 
    -0.001669819, -0.001584127, -0.001403663, -0.001380195, -0.001297456, 
    -0.001157774, -0.001110323, -0.001019611, -0.000882791, -0.0008385051,
  -0.000353054, -0.0003947018, -0.0006395692, -0.0009254474, -0.001249452, 
    -0.001497696, -0.001682983, -0.001815463, -0.001929441, -0.001988941, 
    -0.001982093, -0.001940616, -0.001830246, -0.001652982, -0.001533642, 
    -0.001300097, -0.000953279, -0.0008609949, -0.0008141239, -0.0008050484, 
    -0.0005507399, -0.0004429788, -0.0004803023, -0.0004910917, 
    -0.0005480435, -0.0006408099, -0.0005922511, -0.000621018, -0.000696274, 
    -0.0006667058, -0.000719007, -0.0008480568, -0.0008992549, -0.001001395, 
    -0.001158293, -0.001209894, -0.001264427, -0.001315849, -0.001458545, 
    -0.00153373, -0.001545564, -0.001707744, -0.001765462, -0.001720383, 
    -0.001729227, -0.001639424, -0.001451818, -0.001408754, -0.001305369, 
    -0.001143806, -0.001078099, -0.0009672729, -0.0008087079, -0.0007588133,
  -0.0001554013, -0.0002024394, -0.0004514646, -0.000730805, -0.00103518, 
    -0.00126118, -0.001431666, -0.001560355, -0.001673457, -0.00174669, 
    -0.001763902, -0.001739499, -0.001629416, -0.001452354, -0.001339708, 
    -0.001120498, -0.0007955714, -0.0006978616, -0.0006414698, -0.0006194532, 
    -0.0003767518, -0.0002694377, -0.0002923133, -0.0002994873, 
    -0.0003521851, -0.0004379288, -0.0004012757, -0.0004358515, 
    -0.0005146292, -0.0005119891, -0.000578895, -0.00071068, -0.0007773411, 
    -0.0008926426, -0.00105707, -0.001119244, -0.001188487, -0.001259305, 
    -0.001429275, -0.001530212, -0.001566054, -0.001750125, -0.001821618, 
    -0.001784256, -0.001788359, -0.001690121, -0.001487046, -0.001411528, 
    -0.001274696, -0.001080533, -0.0009822194, -0.0008193144, -0.0005941552, 
    -0.0005266694,
  5.202551e-05, -5.975933e-08, -0.0002440114, -0.0005083883, -0.0007884474, 
    -0.0009920225, -0.001149451, -0.001273054, -0.001376156, -0.001445085, 
    -0.001465332, -0.00144807, -0.001354395, -0.001187172, -0.001085888, 
    -0.0008829634, -0.0005798672, -0.0004765484, -0.000406367, -0.0003603225, 
    -0.0001148326, 3.999324e-06, -4.789471e-06, -1.213433e-05, -7.049889e-05, 
    -0.0001686745, -0.0001616439, -0.0002216941, -0.0003245477, 
    -0.0003526612, -0.0004399205, -0.0005758607, -0.0006605837, 
    -0.0007869213, -0.0009568032, -0.001029572, -0.001115272, -0.001208968, 
    -0.001411912, -0.001540928, -0.001599555, -0.001809607, -0.001893656, 
    -0.001855046, -0.001839801, -0.001713722, -0.001474567, -0.001351488, 
    -0.001165495, -0.0009201632, -0.0007833118, -0.0005800149, -0.0003123718, 
    -0.0002341278,
  0.0001891807, 0.0001260569, -0.0001047501, -0.0003463227, -0.000597906, 
    -0.0007799409, -0.0009265387, -0.001042868, -0.001126131, -0.00116853, 
    -0.001160426, -0.00114135, -0.001052737, -0.0008914029, -0.0007998224, 
    -0.0006114191, -0.0003274889, -0.0002156489, -0.0001310329, 
    -6.570102e-05, 0.0001728473, 0.0002931435, 0.0002943381, 0.0002868154, 
    0.0002220119, 0.0001084079, 8.339177e-05, -5.232434e-06, -0.0001406637, 
    -0.0002009451, -0.0003012104, -0.0004373325, -0.0005391164, 
    -0.0006769355, -0.0008524921, -0.0009362835, -0.001039105, -0.001156601, 
    -0.001393848, -0.001552077, -0.001634407, -0.00187149, -0.001968601, 
    -0.001928691, -0.001893318, -0.001738275, -0.001461584, -0.001289026, 
    -0.001051888, -0.0007533247, -0.0005763812, -0.0003310633, 7.553153e-06, 
    0.000106642,
  0.0002782255, 0.0001966404, -3.259814e-05, -0.0002620253, -0.0004909892, 
    -0.0006519437, -0.000784538, -0.0008932376, -0.0009697781, -0.001014611, 
    -0.001019409, -0.0009868287, -0.0008880639, -0.0007258112, -0.0006381251, 
    -0.0004546248, -0.00017598, -4.379717e-05, 6.564717e-05, 0.0001587323, 
    0.0004010612, 0.0005330313, 0.0005527027, 0.0005592728, 0.0004959348, 
    0.0003693981, 0.0003203638, 0.0002060009, 4.082366e-05, -5.076884e-05, 
    -0.0002096249, -0.0003682923, -0.0005055362, -0.0006701121, 
    -0.0008591077, -0.0009574547, -0.001078323, -0.001219871, -0.001494067, 
    -0.001682242, -0.001786488, -0.002055976, -0.002154454, -0.002089889, 
    -0.002007166, -0.001791629, -0.001439255, -0.001177105, -0.0008465734, 
    -0.0004529195, -0.0002008215, 0.0001380397, 0.0005601167, 0.0006848875,
  -0.0001237267, -0.0002187413, -0.0004019013, -0.0005797548, -0.0007640507, 
    -0.0009024202, -0.001025008, -0.001115483, -0.001146122, -0.001112985, 
    -0.00102421, -0.000904303, -0.0007717037, -0.0006193661, -0.0005402862, 
    -0.0003623799, -8.621277e-05, 6.892671e-05, 0.0002114917, 0.0003468697, 
    0.0006078605, 0.0007387492, 0.0007669548, 0.0007841025, 0.0007166002, 
    0.000562285, 0.0004749483, 0.0003180479, 8.714318e-05, -6.953639e-05, 
    -0.0002237195, -0.0003686455, -0.0005161634, -0.0006854259, 
    -0.0008739735, -0.0009820473, -0.001122708, -0.001294402, -0.001612469, 
    -0.001832174, -0.001955285, -0.002258768, -0.002362543, -0.00227334, 
    -0.002138702, -0.001853625, -0.001414712, -0.001056893, -0.0006289692, 
    -0.0001353827, 0.0001896439, 0.0006042062, 0.001117483, 0.001273007,
  -0.0007868812, -0.0009066257, -0.001082973, -0.001243484, -0.001397855, 
    -0.001508462, -0.001605469, -0.001675395, -0.001700209, -0.001678679, 
    -0.001617524, -0.001517839, -0.001378333, -0.001199723, -0.001101209, 
    -0.0008935796, -0.0005753654, -0.0003543613, -0.0001421431, 6.183512e-05, 
    0.0003684204, 0.0005706206, 0.0006672649, 0.0007438556, 0.0007116491, 
    0.0005688603, 0.0004842092, 0.000320708, 7.469134e-05, -0.0001735381, 
    -0.000389331, -0.0005524544, -0.0007350633, -0.0009312714, -0.001132895, 
    -0.001258857, -0.001425515, -0.001634257, -0.002005242, -0.002264083, 
    -0.002411572, -0.002763269, -0.00285945, -0.002714554, -0.002491317, 
    -0.002096484, -0.001526817, -0.001028992, -0.0004566192, 0.0001837526, 
    0.0006145677, 0.001146507, 0.001779202, 0.001975492,
  -0.002714143, -0.002830622, -0.002919963, -0.00299446, -0.00307821, 
    -0.003156137, -0.003227834, -0.003255082, -0.003218418, -0.003094209, 
    -0.002909221, -0.002685897, -0.002462551, -0.002237645, -0.00210238, 
    -0.001844069, -0.001458153, -0.001144748, -0.0008395069, -0.0005486565, 
    -0.000178135, 9.242299e-05, 0.0002631707, 0.0004117932, 0.000424745, 
    0.0002902207, 0.000197915, 1.332536e-05, -0.0002885141, -0.0005134539, 
    -0.0006950803, -0.0008344278, -0.001053082, -0.001277075, -0.001490066, 
    -0.001636666, -0.001833775, -0.002085471, -0.002511871, -0.00281196, 
    -0.002985362, -0.00338865, -0.003473, -0.0032622, -0.002938009, 
    -0.002420957, -0.00170837, -0.001058573, -0.0003325916, 0.0004605901, 
    0.0009987871, 0.0016438, 0.002397869, 0.002632917,
  -0.005173279, -0.005276479, -0.005278339, -0.005268782, -0.005284329, 
    -0.00533614, -0.00538385, -0.005366551, -0.005275084, -0.005052278, 
    -0.004744313, -0.004393633, -0.004150604, -0.003917402, -0.003754474, 
    -0.003439579, -0.002969112, -0.00253772, -0.002087691, -0.00162396, 
    -0.001095446, -0.000693768, -0.0004188561, -0.0001740086, -9.410504e-05, 
    -0.0002001032, -0.0002889543, -0.0004857493, -0.0008359228, -0.001127662, 
    -0.001342808, -0.001458286, -0.001655006, -0.001853029, -0.002039409, 
    -0.002200766, -0.002442666, -0.002768337, -0.003277625, -0.003631451, 
    -0.003829513, -0.00429754, -0.004378792, -0.004092114, -0.003640338, 
    -0.00296499, -0.002063957, -0.001214527, -0.0003040488, 0.0006603632, 
    0.001317732, 0.002083956, 0.002960812, 0.00323013,
  -0.008129088, -0.00821337, -0.008147089, -0.008099307, -0.008078169, 
    -0.008112628, -0.008125878, -0.008070482, -0.007999342, -0.007827038, 
    -0.007589536, -0.007288013, -0.006990054, -0.006693684, -0.006451047, 
    -0.006024143, -0.005406963, -0.004782198, -0.004127509, -0.003452559, 
    -0.002729902, -0.002128017, -0.001645834, -0.001239475, -0.001030343, 
    -0.001034757, -0.001067899, -0.001218573, -0.001560712, -0.001896947, 
    -0.002129518, -0.002213735, -0.002432514, -0.002627504, -0.002775901, 
    -0.002972059, -0.003276697, -0.003693861, -0.004279713, -0.004683542, 
    -0.004903916, -0.005435145, -0.005482663, -0.005070903, -0.004429705, 
    -0.003549012, -0.002424737, -0.001324192, -0.0001995126, 0.0009400283, 
    0.001715647, 0.002601187, 0.00359479, 0.003869441,
  -0.01153912, -0.01160987, -0.01154369, -0.01147613, -0.0114397, 
    -0.01150824, -0.01153179, -0.01145445, -0.01139376, -0.01119807, 
    -0.0109114, -0.0105485, -0.01019402, -0.009846844, -0.009516151, 
    -0.008961977, -0.008177011, -0.007327024, -0.006430869, -0.005499429, 
    -0.004523525, -0.003682629, -0.00297675, -0.002413459, -0.002078267, 
    -0.001989672, -0.002018757, -0.002173206, -0.002496886, -0.002801805, 
    -0.003004079, -0.003016408, -0.003256013, -0.003426696, -0.003493849, 
    -0.003734662, -0.004118655, -0.004648061, -0.005312985, -0.005761361, 
    -0.005991343, -0.006588566, -0.006592201, -0.006028443, -0.005150159, 
    -0.004025014, -0.002644039, -0.001246986, 0.0001114283, 0.001419856, 
    0.002302766, 0.003299947, 0.004399999, 0.004653766,
  -0.01447437, -0.0145334, -0.01448915, -0.01444824, -0.01443952, -0.0145732, 
    -0.01462601, -0.01454757, -0.01454456, -0.01439779, -0.01414723, 
    -0.01380515, -0.01344925, -0.01308033, -0.01266753, -0.01198076, 
    -0.01101371, -0.009920503, -0.008754436, -0.007522237, -0.006220817, 
    -0.005079367, -0.004102172, -0.003379986, -0.00291734, -0.002726436, 
    -0.002775258, -0.002957059, -0.003310738, -0.00367755, -0.003844816, 
    -0.003748568, -0.004022467, -0.004146916, -0.004075689, -0.004372245, 
    -0.004858615, -0.005531119, -0.006288916, -0.006788951, -0.007032272, 
    -0.007730919, -0.00769582, -0.006955134, -0.005782809, -0.004363333, 
    -0.002684723, -0.0009455389, 0.0006738446, 0.002159294, 0.00313334, 
    0.004223512, 0.005413092, 0.005621506,
  -0.01661164, -0.0166655, -0.0166902, -0.01671802, -0.01676855, -0.01698974, 
    -0.01708747, -0.01702716, -0.01712179, -0.01708358, -0.01693942, 
    -0.01668617, -0.01637661, -0.01601408, -0.01553398, -0.01471266, 
    -0.01354686, -0.01220735, -0.01075708, -0.009193746, -0.007486519, 
    -0.005977011, -0.004677704, -0.003805646, -0.003232115, -0.002955599, 
    -0.003070495, -0.003333779, -0.003767762, -0.004212469, -0.004364518, 
    -0.004152414, -0.004551985, -0.004635613, -0.00436982, -0.004737679, 
    -0.005354994, -0.006211052, -0.007094864, -0.007686416, -0.007991324, 
    -0.008896207, -0.008880457, -0.007974745, -0.006469647, -0.004702394, 
    -0.002664293, -0.0005317127, 0.001394648, 0.003098093, 0.004148939, 
    0.00531042, 0.006572965, 0.006719056,
  -0.01786526, -0.01790879, -0.01802664, -0.01813931, -0.01825774, 
    -0.01857311, -0.01872842, -0.01870554, -0.01892195, -0.01901716, 
    -0.01900243, -0.01885526, -0.018601, -0.01824768, -0.01771517, 
    -0.01674826, -0.01534726, -0.0137734, -0.01204292, -0.01014473, 
    -0.007948139, -0.006003918, -0.0043342, -0.003332716, -0.002691968, 
    -0.002396716, -0.002659653, -0.003105408, -0.003739077, -0.004330323, 
    -0.00449558, -0.004147636, -0.004744194, -0.004808249, -0.004282688, 
    -0.004740772, -0.005528088, -0.006628983, -0.007701979, -0.008472523, 
    -0.008948458, -0.01023567, -0.01038782, -0.009427016, -0.007621941, 
    -0.00548963, -0.003023658, -0.0004207786, 0.001886516, 0.003888486, 
    0.005022346, 0.006269501, 0.007630451, 0.00772072,
  -0.01814218, -0.01817246, -0.018404, -0.01860255, -0.01877015, -0.01915835, 
    -0.01935683, -0.01936675, -0.01973871, -0.02001113, -0.02018304, 
    -0.02020859, -0.02004018, -0.01969008, -0.01913043, -0.01799514, 
    -0.01628737, -0.01450992, -0.01250487, -0.01025539, -0.007429889, 
    -0.004949273, -0.00283961, -0.0017138, -0.001061565, -0.0008574337, 
    -0.001359492, -0.002103863, -0.003072152, -0.003858411, -0.004054317, 
    -0.003587845, -0.004419658, -0.004440526, -0.00368821, -0.004246082, 
    -0.005200722, -0.006540264, -0.007820711, -0.008782379, -0.009431003, 
    -0.01109695, -0.01149067, -0.0106036, -0.008622719, -0.006255602, 
    -0.003496736, -0.000519195, 0.002092779, 0.004340416, 0.005545459, 
    0.006895543, 0.008385983, 0.008484509,
  -0.01680728, -0.01691758, -0.01734511, -0.01772142, -0.01803534, 
    -0.0185621, -0.01888825, -0.01902608, -0.01964319, -0.02011707, 
    -0.02042959, -0.02054065, -0.02042701, -0.02009232, -0.01951973, 
    -0.01822703, -0.0162165, -0.01429881, -0.01205046, -0.00944424, 
    -0.005981697, -0.002996339, -0.0005161059, 0.0007699434, 0.001397692, 
    0.001383441, 0.0005753271, -0.0005190186, -0.001853735, -0.002882357, 
    -0.003122316, -0.002957647, -0.004610718, -0.005299064, -0.004794791, 
    -0.005434851, -0.006230588, -0.007279339, -0.008248164, -0.009061082, 
    -0.00966406, -0.01138217, -0.01176468, -0.01086074, -0.008805216, 
    -0.006393409, -0.003652782, -0.0008406521, 0.001686918, 0.003933656, 
    0.005050758, 0.006227788, 0.007552321, 0.007622677,
  -0.01507635, -0.01530034, -0.01588822, -0.01645598, -0.01699751, 
    -0.01780144, -0.01842244, -0.01886356, -0.0198478, -0.02065273, 
    -0.02125929, -0.02150459, -0.02150424, -0.02127981, -0.02092064, 
    -0.01970324, -0.01762791, -0.01561638, -0.01324783, -0.01057269, 
    -0.00716362, -0.004351705, -0.002111482, -0.0009064383, -0.0006180116, 
    -0.001349101, -0.002856641, -0.004770211, -0.007383614, -0.01001499, 
    -0.01156099, -0.0118355, -0.0136444, -0.01408246, -0.01300097, 
    -0.0133361, -0.01372082, -0.01421667, -0.01432758, -0.01444405, 
    -0.01453028, -0.01582619, -0.01606569, -0.01530277, -0.01310878, 
    -0.01067768, -0.008034721, -0.005413503, -0.002990036, -0.0007799426, 
    0.0003216421, 0.001553498, 0.002952414, 0.00294249,
  -0.01353696, -0.0139357, -0.01487791, -0.01579791, -0.01669764, 
    -0.01774718, -0.01869689, -0.0195429, -0.02085435, -0.02203352, 
    -0.0230636, -0.02372963, -0.02411445, -0.0242444, -0.02441453, 
    -0.02357454, -0.02172344, -0.02024994, -0.01829799, -0.01590598, 
    -0.01268792, -0.01015223, -0.008297267, -0.007167249, -0.007060143, 
    -0.008042301, -0.009774798, -0.01189223, -0.01457155, -0.01723834, 
    -0.01878531, -0.01908257, -0.02091993, -0.02107332, -0.01947025, 
    -0.01963102, -0.01981854, -0.02005855, -0.01962443, -0.01932065, 
    -0.01914567, -0.02067381, -0.02120264, -0.02078196, -0.01846715, 
    -0.01585573, -0.01295693, -0.009860804, -0.007134074, -0.004798823, 
    -0.003690558, -0.002536996, -0.001322513, -0.001282124,
  -0.01137528, -0.01183311, -0.01293976, -0.01410502, -0.01531905, 
    -0.01666579, -0.01796801, -0.01923382, -0.02082993, -0.02247943, 
    -0.02415375, -0.02557242, -0.02678723, -0.02781319, -0.02922837, 
    -0.02924092, -0.02785742, -0.02743047, -0.02588308, -0.02325115, 
    -0.01956372, -0.01652975, -0.01413612, -0.01252346, -0.01219522, 
    -0.01319071, -0.01456176, -0.01670427, -0.01975282, -0.02240577, 
    -0.0238708, -0.02407633, -0.02571985, -0.02535762, -0.0229766, 
    -0.02278353, -0.02282085, -0.02308325, -0.02293949, -0.02302267, 
    -0.02335409, -0.02557969, -0.02656111, -0.02633913, -0.02359609, 
    -0.02044868, -0.01689351, -0.01276335, -0.009202678, -0.006238495, 
    -0.005393143, -0.00441085, -0.003290274, -0.003254484,
  -0.011168, -0.01141308, -0.01257805, -0.01386545, -0.01527551, -0.01678868, 
    -0.01845448, -0.02027084, -0.02216487, -0.02435635, -0.02683435, 
    -0.02944029, -0.03232622, -0.0355, -0.03906537, -0.04011731, -0.03866333, 
    -0.03942344, -0.0374087, -0.03262757, -0.02578416, -0.02017727, 
    -0.01582181, -0.01246179, -0.01130296, -0.01234809, -0.01327673, 
    -0.01557297, -0.0192419, -0.02222205, -0.02386646, -0.02414845, 
    -0.02590232, -0.02505979, -0.02162086, -0.02110543, -0.02102003, 
    -0.02136469, -0.0222237, -0.02352368, -0.0252646, -0.03028716, 
    -0.03307343, -0.0336234, -0.03121795, -0.02724958, -0.02171827, 
    -0.01554652, -0.01029023, -0.005949402, -0.005315721, -0.004446652, 
    -0.003342198, -0.003301376 ;

 v_east =
  -0.001153907, -8.673617e-19, -8.673617e-19, 0, -8.673617e-19, 0, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 0, 0, 0, 
    -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.001418448, -8.673617e-19, -8.673617e-19, 0, -8.673617e-19, 0, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 0, 0, 0, 
    -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.001644929, -8.673617e-19, -8.673617e-19, 0, -8.673617e-19, 0, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 0, 0, 0, 
    -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.001839962, -8.673617e-19, -8.673617e-19, 0, -8.673617e-19, 0, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 0, 0, 0, 
    -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.002083743, -8.673617e-19, -8.673617e-19, 0, -8.673617e-19, 0, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 0, 0, 0, 
    -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.002687964, -8.673617e-19, -8.673617e-19, 0, -8.673617e-19, 0, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 0, 0, 0, 
    -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.003229869, -8.673617e-19, -8.673617e-19, 0, -8.673617e-19, 0, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 0, 0, 0, 
    -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.003728156, -8.673617e-19, -8.673617e-19, 0, -8.673617e-19, 0, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 0, 0, 0, 
    -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.004200587, -8.673617e-19, -8.673617e-19, 0, -8.673617e-19, 0, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 0, 0, 0, 
    -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.004589796, -8.673617e-19, -8.673617e-19, 0, -8.673617e-19, 0, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 0, 0, 0, 
    -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.004905125, -8.673617e-19, -8.673617e-19, 0, -8.673617e-19, 0, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 0, 0, 0, 
    -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.005231532, -8.673617e-19, -8.673617e-19, 0, -8.673617e-19, 0, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 0, 0, 0, 
    -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.005588669, -8.673617e-19, -8.673617e-19, 0, -8.673617e-19, 0, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 0, 0, 0, 
    -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.006385055, -8.673617e-19, -8.673617e-19, 0, -8.673617e-19, 0, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 0, 0, 0, 
    -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.007196248, -8.673617e-19, -8.673617e-19, 0, -8.673617e-19, 0, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 0, 0, 0, 
    -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.008533215, -8.673617e-19, -8.673617e-19, 0, -8.673617e-19, 0, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 0, 0, 0, 
    -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.009760018, -8.673617e-19, -8.673617e-19, 0, -8.673617e-19, 0, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 0, 0, 0, 
    -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.00974746, -8.673617e-19, -8.673617e-19, 0, -8.673617e-19, 0, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 0, 0, 0, 
    -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.01016604, -8.673617e-19, -8.673617e-19, 0, -8.673617e-19, 0, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 0, 0, 0, 
    -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.01126966, -8.673617e-19, -8.673617e-19, 0, -8.673617e-19, 0, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 0, 0, 0, 
    -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.01275358, -8.673617e-19, -8.673617e-19, 0, -8.673617e-19, 0, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 0, 0, 0, 
    -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.01543826, -8.673617e-19, -8.673617e-19, 0, -8.673617e-19, 0, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 0, 0, 0, 
    -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.01757964, -8.673617e-19, -8.673617e-19, 0, -8.673617e-19, 0, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 0, 0, 0, 
    -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.0212019, -8.673617e-19, -8.673617e-19, 0, -8.673617e-19, 0, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 0, 0, 0, 
    -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.02426313, -8.673617e-19, -8.673617e-19, 0, -8.673617e-19, 0, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 0, 0, 0, 
    -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.02671312, -8.673617e-19, -8.673617e-19, 0, -8.673617e-19, 0, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 0, 0, 0, 
    -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.02829143, -8.673617e-19, -8.673617e-19, 0, -8.673617e-19, 0, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 0, 0, 0, 
    -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.02829143, -8.673617e-19, -8.673617e-19, 0, -8.673617e-19, 0, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 0, 0, 0, 
    -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.02829143, -8.673617e-19, -8.673617e-19, 0, -8.673617e-19, 0, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 0, 0, 0, 
    -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.02829143, -8.673617e-19, -8.673617e-19, 0, -8.673617e-19, 0, 
    8.673617e-19, 8.673617e-19, 8.673617e-19, -8.673617e-19, 0, 0, 0, 
    -8.673617e-19, 8.673617e-19, 8.673617e-19, 0, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  0.0009126041, 0, -1.734723e-18, 0, -8.673617e-19, 2.602085e-18, 
    1.734723e-18, 0, 0, 1.734723e-18, 1.734723e-18, 1.734723e-18, 0, 
    -8.673617e-19, 1.734723e-18, -8.673617e-19, 1.734723e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  0.0006527598, 0, -1.734723e-18, 0, -8.673617e-19, 2.602085e-18, 
    1.734723e-18, 0, 0, 1.734723e-18, 1.734723e-18, 1.734723e-18, 0, 
    -8.673617e-19, 1.734723e-18, -8.673617e-19, 1.734723e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  0.0004303, 0, -1.734723e-18, 0, -8.673617e-19, 2.602085e-18, 1.734723e-18, 
    0, 0, 1.734723e-18, 1.734723e-18, 1.734723e-18, 0, -8.673617e-19, 
    1.734723e-18, -8.673617e-19, 1.734723e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18,
  0.0002387293, 0, -1.734723e-18, 0, -8.673617e-19, 2.602085e-18, 
    1.734723e-18, 0, 0, 1.734723e-18, 1.734723e-18, 1.734723e-18, 0, 
    -8.673617e-19, 1.734723e-18, -8.673617e-19, 1.734723e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  8.022677e-06, 0, -1.734723e-18, 0, -8.673617e-19, 2.602085e-18, 
    1.734723e-18, 0, 0, 1.734723e-18, 1.734723e-18, 1.734723e-18, 0, 
    -8.673617e-19, 1.734723e-18, -8.673617e-19, 1.734723e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.0005317287, 0, -1.734723e-18, 0, -8.673617e-19, 2.602085e-18, 
    1.734723e-18, 0, 0, 1.734723e-18, 1.734723e-18, 1.734723e-18, 0, 
    -8.673617e-19, 1.734723e-18, -8.673617e-19, 1.734723e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.001015814, 0, -1.734723e-18, 0, -8.673617e-19, 2.602085e-18, 
    1.734723e-18, 0, 0, 1.734723e-18, 1.734723e-18, 1.734723e-18, 0, 
    -8.673617e-19, 1.734723e-18, -8.673617e-19, 1.734723e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.001460935, 0, -1.734723e-18, 0, -8.673617e-19, 2.602085e-18, 
    1.734723e-18, 0, 0, 1.734723e-18, 1.734723e-18, 1.734723e-18, 0, 
    -8.673617e-19, 1.734723e-18, -8.673617e-19, 1.734723e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.001882958, 0, -1.734723e-18, 0, -8.673617e-19, 2.602085e-18, 
    1.734723e-18, 0, 0, 1.734723e-18, 1.734723e-18, 1.734723e-18, 0, 
    -8.673617e-19, 1.734723e-18, -8.673617e-19, 1.734723e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.002275933, 0, -1.734723e-18, 0, -8.673617e-19, 2.602085e-18, 
    1.734723e-18, 0, 0, 1.734723e-18, 1.734723e-18, 1.734723e-18, 0, 
    -8.673617e-19, 1.734723e-18, -8.673617e-19, 1.734723e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.002651452, 0, -1.734723e-18, 0, -8.673617e-19, 2.602085e-18, 
    1.734723e-18, 0, 0, 1.734723e-18, 1.734723e-18, 1.734723e-18, 0, 
    -8.673617e-19, 1.734723e-18, -8.673617e-19, 1.734723e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.003040162, 0, -1.734723e-18, 0, -8.673617e-19, 2.602085e-18, 
    1.734723e-18, 0, 0, 1.734723e-18, 1.734723e-18, 1.734723e-18, 0, 
    -8.673617e-19, 1.734723e-18, -8.673617e-19, 1.734723e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.003463293, 0, -1.734723e-18, 0, -8.673617e-19, 2.602085e-18, 
    1.734723e-18, 0, 0, 1.734723e-18, 1.734723e-18, 1.734723e-18, 0, 
    -8.673617e-19, 1.734723e-18, -8.673617e-19, 1.734723e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.004349034, 0, -1.734723e-18, 0, -8.673617e-19, 2.602085e-18, 
    1.734723e-18, 0, 0, 1.734723e-18, 1.734723e-18, 1.734723e-18, 0, 
    -8.673617e-19, 1.734723e-18, -8.673617e-19, 1.734723e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.005251244, 0, -1.734723e-18, 0, -8.673617e-19, 2.602085e-18, 
    1.734723e-18, 0, 0, 1.734723e-18, 1.734723e-18, 1.734723e-18, 0, 
    -8.673617e-19, 1.734723e-18, -8.673617e-19, 1.734723e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.006366655, 0, -1.734723e-18, 0, -8.673617e-19, 2.602085e-18, 
    1.734723e-18, 0, 0, 1.734723e-18, 1.734723e-18, 1.734723e-18, 0, 
    -8.673617e-19, 1.734723e-18, -8.673617e-19, 1.734723e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.007360656, 0, -1.734723e-18, 0, -8.673617e-19, 2.602085e-18, 
    1.734723e-18, 0, 0, 1.734723e-18, 1.734723e-18, 1.734723e-18, 0, 
    -8.673617e-19, 1.734723e-18, -8.673617e-19, 1.734723e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.007446561, 0, -1.734723e-18, 0, -8.673617e-19, 2.602085e-18, 
    1.734723e-18, 0, 0, 1.734723e-18, 1.734723e-18, 1.734723e-18, 0, 
    -8.673617e-19, 1.734723e-18, -8.673617e-19, 1.734723e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.008146564, 0, -1.734723e-18, 0, -8.673617e-19, 2.602085e-18, 
    1.734723e-18, 0, 0, 1.734723e-18, 1.734723e-18, 1.734723e-18, 0, 
    -8.673617e-19, 1.734723e-18, -8.673617e-19, 1.734723e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.009827083, 0, -1.734723e-18, 0, -8.673617e-19, 2.602085e-18, 
    1.734723e-18, 0, 0, 1.734723e-18, 1.734723e-18, 1.734723e-18, 0, 
    -8.673617e-19, 1.734723e-18, -8.673617e-19, 1.734723e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.01180771, 0, -1.734723e-18, 0, -8.673617e-19, 2.602085e-18, 
    1.734723e-18, 0, 0, 1.734723e-18, 1.734723e-18, 1.734723e-18, 0, 
    -8.673617e-19, 1.734723e-18, -8.673617e-19, 1.734723e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.01494399, 0, -1.734723e-18, 0, -8.673617e-19, 2.602085e-18, 
    1.734723e-18, 0, 0, 1.734723e-18, 1.734723e-18, 1.734723e-18, 0, 
    -8.673617e-19, 1.734723e-18, -8.673617e-19, 1.734723e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.01744559, 0, -1.734723e-18, 0, -8.673617e-19, 2.602085e-18, 
    1.734723e-18, 0, 0, 1.734723e-18, 1.734723e-18, 1.734723e-18, 0, 
    -8.673617e-19, 1.734723e-18, -8.673617e-19, 1.734723e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.02159326, 0, -1.734723e-18, 0, -8.673617e-19, 2.602085e-18, 
    1.734723e-18, 0, 0, 1.734723e-18, 1.734723e-18, 1.734723e-18, 0, 
    -8.673617e-19, 1.734723e-18, -8.673617e-19, 1.734723e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.02509251, 0, -1.734723e-18, 0, -8.673617e-19, 2.602085e-18, 
    1.734723e-18, 0, 0, 1.734723e-18, 1.734723e-18, 1.734723e-18, 0, 
    -8.673617e-19, 1.734723e-18, -8.673617e-19, 1.734723e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.02789306, 0, -1.734723e-18, 0, -8.673617e-19, 2.602085e-18, 
    1.734723e-18, 0, 0, 1.734723e-18, 1.734723e-18, 1.734723e-18, 0, 
    -8.673617e-19, 1.734723e-18, -8.673617e-19, 1.734723e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.0296925, 0, -1.734723e-18, 0, -8.673617e-19, 2.602085e-18, 1.734723e-18, 
    0, 0, 1.734723e-18, 1.734723e-18, 1.734723e-18, 0, -8.673617e-19, 
    1.734723e-18, -8.673617e-19, 1.734723e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.0296925, 0, -1.734723e-18, 0, -8.673617e-19, 2.602085e-18, 1.734723e-18, 
    0, 0, 1.734723e-18, 1.734723e-18, 1.734723e-18, 0, -8.673617e-19, 
    1.734723e-18, -8.673617e-19, 1.734723e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.0296925, 0, -1.734723e-18, 0, -8.673617e-19, 2.602085e-18, 1.734723e-18, 
    0, 0, 1.734723e-18, 1.734723e-18, 1.734723e-18, 0, -8.673617e-19, 
    1.734723e-18, -8.673617e-19, 1.734723e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.0296925, 0, -1.734723e-18, 0, -8.673617e-19, 2.602085e-18, 1.734723e-18, 
    0, 0, 1.734723e-18, 1.734723e-18, 1.734723e-18, 0, -8.673617e-19, 
    1.734723e-18, -8.673617e-19, 1.734723e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18 ;

 v_south =
  -0.002053349, -0.002232674, -0.00257489, -0.003046317, -0.003558519, 
    -0.003940778, -0.004115353, -0.004436044, -0.005051654, -0.005588714, 
    -0.006111963, -0.006013229, -0.005305474, -0.004635567, -0.004091095, 
    -0.003657248, -0.00321911, -0.002828628, -0.002590592, -0.002374522, 
    -0.002150663, -0.001900998, -0.001652628, -0.001366461, -0.001003114, 
    -0.0005792573, -0.0002656453, -2.970293e-05, 0.0002033381, 0.0003372525, 
    0.0004304121, 0.0005712219, 0.0006166759, 0.0005493091, 0.0004578765, 
    0.0002645368, 1.74565e-05, -0.0002158243, -0.000427264, -0.0006965995, 
    -0.001071399, -0.001387975, -0.00143774, -0.00123382, -0.001122162, 
    -0.0009449027, -0.0003406468, -0.0001278573, -2.666071e-05, 
    -0.0002690725, -0.0004120498, -0.0002926496, -0.0001140157, 
    -0.0007223942, -0.002307813, -0.001153907,
  -0.0009936204, -0.0009547506, -0.001354037, -0.001876029, -0.00248574, 
    -0.003247505, -0.004177494, -0.005240373, -0.005990713, -0.006517528, 
    -0.007005468, -0.006790339, -0.006025404, -0.00522816, -0.004495075, 
    -0.003848777, -0.003196434, -0.002639435, -0.002388867, -0.002149342, 
    -0.001876249, -0.001555096, -0.00123121, -0.0009266738, -0.0005812812, 
    -0.0002230267, 6.042036e-05, 0.0003160779, 0.0005713619, 0.0007025342, 
    0.0007647762, 0.0008420494, 0.0008681939, 0.0007749898, 0.0006681144, 
    0.0003426897, -0.000189194, -0.0007151664, -0.001105537, -0.001473593, 
    -0.001827293, -0.00181704, -0.001508578, -0.001273061, -0.001047287, 
    -0.0006775317, -0.0002551764, 7.324323e-05, -0.0002506819, -0.0004314595, 
    -0.0005218355, -0.0003534999, -0.0002493233, -0.00102298, -0.002836895, 
    -0.001418448,
  -0.0009881345, -0.000949075, -0.001353847, -0.001850687, -0.002345843, 
    -0.00310019, -0.00413444, -0.005154299, -0.005826725, -0.006317762, 
    -0.006815941, -0.006610912, -0.005839287, -0.005060729, -0.004355893, 
    -0.003722808, -0.003084179, -0.002528108, -0.002253539, -0.001989346, 
    -0.00169986, -0.001368523, -0.001033748, -0.0007166195, -0.0003561712, 
    1.846349e-05, 0.0003119753, 0.0005719459, 0.0008314765, 0.0009659154, 
    0.001027762, 0.00110716, 0.001128917, 0.001030205, 0.0009082331, 
    0.0005815312, 5.944907e-05, -0.0004572175, -0.0008444691, -0.001211678, 
    -0.001565737, -0.001618111, -0.001419131, -0.00124011, -0.0009465492, 
    -0.0005807236, -0.0001576686, -5.784886e-05, -0.0004688656, 
    -0.0005854516, -0.0006506416, -0.000579821, -0.0004791759, -0.00128022, 
    -0.003289857, -0.001644929,
  -0.0009793601, -0.0009403558, -0.001348121, -0.001850111, -0.002352624, 
    -0.003086744, -0.004068193, -0.005030028, -0.005653301, -0.006106529, 
    -0.006568523, -0.00636322, -0.005628441, -0.004884052, -0.004204252, 
    -0.003587384, -0.002963668, -0.002404687, -0.002108633, -0.001825933, 
    -0.00152062, -0.001177435, -0.0008314252, -0.0005015055, -0.0001319194, 
    0.0002507314, 0.0005509804, 0.0008163358, 0.001081286, 0.001219422, 
    0.001280818, 0.00135838, 0.001366952, 0.001237838, 0.001085027, 
    0.0007546723, 0.0002457662, -0.0002607005, -0.0006487001, -0.001020737, 
    -0.001382902, -0.001467488, -0.001286498, -0.001119442, -0.0008453129, 
    -0.0005109044, -6.599428e-05, -0.0003163332, -0.0006563948, 
    -0.0007178281, -0.00076139, -0.0007956019, -0.0007665944, -0.001644504, 
    -0.003679924, -0.001839962,
  -0.0009674193, -0.0009291182, -0.001337797, -0.001840626, -0.002343948, 
    -0.003052209, -0.003979859, -0.004889355, -0.005468989, -0.005883302, 
    -0.006305726, -0.006099514, -0.005406487, -0.004704559, -0.004054647, 
    -0.003455227, -0.002849462, -0.002294147, -0.001982892, -0.001685681, 
    -0.00136741, -0.001013614, -0.0006569183, -0.0003173414, 5.288095e-05, 
    0.0004312051, 0.0007298551, 0.0009967342, 0.001263401, 0.001400576, 
    0.001455864, 0.001520215, 0.00149778, 0.001344549, 0.001177177, 
    0.0008463623, 0.0003445688, -0.000154963, -0.0005374214, -0.0009005229, 
    -0.001254482, -0.001341115, -0.001171531, -0.001037752, -0.00081743, 
    -0.0004860368, -3.460961e-05, -0.0005404171, -0.0008189849, 
    -0.0008326193, -0.0008574477, -0.0009828159, -0.001016066, -0.001987571, 
    -0.004167487, -0.002083743,
  -0.0009430419, -0.0009050758, -0.001313132, -0.001817825, -0.002326507, 
    -0.003014653, -0.003889554, -0.004740944, -0.005275385, -0.005657175, 
    -0.006048339, -0.005844691, -0.005188161, -0.004520602, -0.003898859, 
    -0.003321414, -0.002737281, -0.002189684, -0.001871655, -0.001567325, 
    -0.001243556, -0.0008868937, -0.0005275343, -0.0001837848, 0.0001884289, 
    0.0005681754, 0.0008668791, 0.001132354, 0.001397631, 0.001531884, 
    0.001581735, 0.001640015, 0.001605269, 0.001438259, 0.0012581, 
    0.0009268813, 0.0004313338, -6.210797e-05, -0.0004397003, -0.0007949545, 
    -0.001172801, -0.001312914, -0.001214027, -0.001110372, -0.0008553144, 
    -0.000464198, -0.0002931413, -0.0007524041, -0.0009744847, -0.0009640575, 
    -0.000972306, -0.001147382, -0.001235455, -0.002289428, -0.005375927, 
    -0.002687964,
  -0.0009055574, -0.0008693087, -0.001275268, -0.001776217, -0.00228089, 
    -0.002942855, -0.003767714, -0.004570663, -0.005066909, -0.005415716, 
    -0.005773258, -0.005573178, -0.004958863, -0.004334266, -0.003745865, 
    -0.003192252, -0.0026324, -0.002095605, -0.001772125, -0.001461425, 
    -0.001132736, -0.0007735099, -0.0004117675, -6.428456e-05, 0.0003097114, 
    0.0006907308, 0.0009855318, 0.00124997, 0.001514547, 0.00164462, 
    0.001684241, 0.001719654, 0.00163674, 0.001410144, 0.001182187, 
    0.000842093, 0.0003588168, -0.0001275168, -0.0005082262, -0.0008756107, 
    -0.001245348, -0.001380187, -0.001279985, -0.001175353, -0.0008892132, 
    -0.000553504, -0.0005244855, -0.0009512053, -0.001122211, -0.001111383, 
    -0.001245443, -0.001429802, -0.00145549, -0.002560028, -0.006459739, 
    -0.003229869,
  -0.0008711594, -0.0008364866, -0.001240522, -0.001738035, -0.00223903, 
    -0.002876968, -0.003655906, -0.004414403, -0.004875599, -0.00519414, 
    -0.005520828, -0.005324022, -0.004748447, -0.004163273, -0.003604253, 
    -0.003072241, -0.002532603, -0.002003207, -0.001678719, -0.001371322, 
    -0.001045415, -0.0006884045, -0.0003284341, 1.573923e-05, 0.0003723693, 
    0.0007276372, 0.001007779, 0.001261216, 0.001514781, 0.001631727, 
    0.001657354, 0.001679069, 0.001578772, 0.001336313, 0.001092572, 
    0.0007492707, 0.0002672912, -0.0002175342, -0.0005915494, -0.0009506446, 
    -0.001311924, -0.001441923, -0.001340514, -0.001260408, -0.001031776, 
    -0.0007934725, -0.0007367991, -0.001133663, -0.001257806, -0.001246629, 
    -0.001496233, -0.001772573, -0.001785469, -0.003225574, -0.007456313, 
    -0.003728156,
  -0.0007742649, -0.000738371, -0.001136715, -0.001633913, -0.002141648, 
    -0.002762342, -0.003487502, -0.00418384, -0.004603869, -0.004899732, 
    -0.005205357, -0.005019511, -0.004482908, -0.003932558, -0.003409397, 
    -0.002913094, -0.002409678, -0.00190359, -0.001588715, -0.001289779, 
    -0.0009726061, -0.0006254481, -0.0002755294, 6.1519e-05, 0.0004102378, 
    0.0007576957, 0.001028844, 0.001271864, 0.001515004, 0.001619519, 
    0.001631896, 0.001640642, 0.001523886, 0.001266408, 0.001007723, 
    0.0006613844, 0.0001806325, -0.0003027649, -0.0006704419, -0.001021689, 
    -0.001391833, -0.0015663, -0.001539288, -0.00150939, -0.001272503, 
    -0.001020686, -0.0009978493, -0.001306433, -0.001386209, -0.001374715, 
    -0.001733777, -0.002097297, -0.002098148, -0.004586473, -0.008401173, 
    -0.004200587,
  -0.0006668865, -0.0006319136, -0.001023917, -0.001511576, -0.002009021, 
    -0.00260202, -0.003280514, -0.003932254, -0.004320451, -0.004590106, 
    -0.004868819, -0.004693246, -0.004203192, -0.003700373, -0.003218457, 
    -0.002757145, -0.002289224, -0.001805975, -0.00150052, -0.001209875, 
    -0.0009012607, -0.0005637569, -0.0002236878, 0.0001063788, 0.0004473453, 
    0.0007871502, 0.00104864, 0.001281386, 0.001514347, 0.001606153, 
    0.001603921, 0.001594578, 0.001448225, 0.001157518, 0.0008679246, 
    0.0005094103, 2.459995e-05, -0.0004642785, -0.0008376199, -0.001209197, 
    -0.001594368, -0.001780339, -0.001768188, -0.001753372, -0.001508394, 
    -0.001243336, -0.001281408, -0.00149153, -0.001527378, -0.00150024, 
    -0.001966581, -0.002415563, -0.002404639, -0.005920589, -0.009179591, 
    -0.004589796,
  -0.0005565076, -0.0005207448, -0.0009060917, -0.001387783, -0.001874815, 
    -0.002439789, -0.003071062, -0.003677673, -0.004031557, -0.004276793, 
    -0.004528275, -0.004363096, -0.003920147, -0.003454929, -0.003005008, 
    -0.002580062, -0.002143837, -0.00167135, -0.001369345, -0.001093822, 
    -0.0008056314, -0.0004874034, -0.0001650335, 0.000152969, 0.0004804299, 
    0.000803599, 0.001049058, 0.001266403, 0.001483945, 0.001556573, 
    0.001535609, 0.001508108, 0.001336754, 0.0010252, 0.0007146564, 
    0.0003448526, -0.0001507251, -0.0006500447, -0.001025159, -0.001405981, 
    -0.001799315, -0.001996925, -0.001999813, -0.002000256, -0.001754873, 
    -0.001534637, -0.001568338, -0.001689011, -0.00173391, -0.00186471, 
    -0.002355044, -0.002737577, -0.002714723, -0.007270253, -0.00981025, 
    -0.004905125,
  -0.0003488836, -0.0003073474, -0.0006741835, -0.001137646, -0.001618106, 
    -0.002156131, -0.002725765, -0.003262256, -0.003575923, -0.003798505, 
    -0.004031201, -0.003883925, -0.003487285, -0.00307179, -0.002674819, 
    -0.002299773, -0.001914435, -0.001480812, -0.001207104, -0.0009575587, 
    -0.0006930668, -0.0003977734, -9.870012e-05, 0.0002022124, 0.000513004, 
    0.0008198945, 0.001049491, 0.001250879, 0.001452447, 0.001505206, 
    0.001464835, 0.001418521, 0.001221263, 0.0008881105, 0.0005558621, 
    0.0001743617, -0.0003323716, -0.0008425087, -0.001219461, -0.00160986, 
    -0.001996247, -0.002188324, -0.002205897, -0.002246014, -0.002044515, 
    -0.001839469, -0.001858079, -0.001893601, -0.001947867, -0.002265691, 
    -0.002933195, -0.003328242, -0.004051844, -0.008579791, -0.01046306, 
    -0.005231532,
  -0.0001310525, -8.403836e-05, -0.0004315037, -0.0008701578, -0.001324093, 
    -0.001821242, -0.002335241, -0.002819451, -0.003099126, -0.003294872, 
    -0.003499708, -0.003368366, -0.003028088, -0.002670855, -0.002329293, 
    -0.002006465, -0.001674379, -0.001281424, -0.001034542, -0.000809114, 
    -0.0005720028, -0.0003035649, -2.928595e-05, 0.0002537427, 0.0005565091, 
    0.0008617725, 0.001086252, 0.001277615, 0.001468818, 0.001508632, 
    0.001459833, 0.001417026, 0.001230615, 0.0009234408, 0.0006078078, 
    0.0002201639, -0.0003131585, -0.0008445567, -0.001232637, -0.001649095, 
    -0.002074768, -0.002320402, -0.002400965, -0.002501795, -0.002347602, 
    -0.00215845, -0.002110954, -0.002123796, -0.002171733, -0.002685208, 
    -0.003538006, -0.003946485, -0.005894303, -0.00926575, -0.01117734, 
    -0.005588669,
  1.012876e-05, 6.929875e-05, -0.0002415124, -0.0006328876, -0.001039073, 
    -0.001481422, -0.001930024, -0.002350201, -0.002587166, -0.002749783, 
    -0.002921405, -0.002801816, -0.002511356, -0.00220163, -0.001909129, 
    -0.001639831, -0.001359388, -0.0009987276, -0.000782864, -0.0005935331, 
    -0.0003855214, -0.0001414689, 0.0001064209, 0.0003799616, 0.0006760419, 
    0.0009739479, 0.001197804, 0.00139379, 0.001589634, 0.001629069, 
    0.001581815, 0.001539868, 0.001335861, 0.001015146, 0.0006869474, 
    0.000287305, -0.0002643574, -0.0008143138, -0.001224928, -0.001686637, 
    -0.002156456, -0.002457807, -0.002590038, -0.002718981, -0.002585367, 
    -0.002378282, -0.002374021, -0.002483472, -0.002675774, -0.003371199, 
    -0.004250653, -0.004589429, -0.007810055, -0.009978855, -0.01277011, 
    -0.006385055,
  9.888375e-05, 0.0001783854, -8.538185e-05, -0.0004219437, -0.0007713183, 
    -0.001146515, -0.001518279, -0.001865464, -0.002055334, -0.002179507, 
    -0.002311467, -0.002198481, -0.001955637, -0.001696126, -0.001456655, 
    -0.001242401, -0.0010185, -0.0007019078, -0.0005263969, -0.0003738496, 
    -0.0001954912, 2.371192e-05, 0.0002462374, 0.0005090336, 0.0007978494, 
    0.001078682, 0.001306171, 0.00151671, 0.001726689, 0.001776039, 
    0.001744363, 0.001729762, 0.001554947, 0.001284366, 0.001001563, 
    0.0006090874, 3.367242e-05, -0.0005342678, -0.0009679082, -0.001469033, 
    -0.0019691, -0.002308957, -0.002517153, -0.002767052, -0.002723286, 
    -0.002595278, -0.002719897, -0.002849981, -0.003294049, -0.004359873, 
    -0.005366941, -0.006681153, -0.009018054, -0.01122858, -0.0143925, 
    -0.007196248,
  -0.0003142593, -0.0002176218, -0.0004131503, -0.000643539, -0.000869787, 
    -0.001135677, -0.001430878, -0.001721907, -0.001864343, -0.001922858, 
    -0.001984687, -0.001856445, -0.001653486, -0.001447255, -0.001258998, 
    -0.001089602, -0.000920053, -0.0006573431, -0.0005403919, -0.0004251774, 
    -0.0002557342, -3.382847e-05, 0.0001875756, 0.0004706689, 0.0007832362, 
    0.001102308, 0.001384124, 0.001663278, 0.001941958, 0.002055342, 
    0.002091683, 0.002142471, 0.001997395, 0.00175417, 0.001500594, 
    0.001118045, 0.0005380262, -3.566894e-05, -0.0005145348, -0.001091792, 
    -0.001668132, -0.002111241, -0.002442888, -0.002811783, -0.002877225, 
    -0.002886372, -0.003135129, -0.003545963, -0.00415567, -0.005464253, 
    -0.006490802, -0.008858933, -0.009951418, -0.01299489, -0.01706643, 
    -0.008533215,
  -0.0009943668, -0.0008680827, -0.0009878421, -0.001132806, -0.001274375, 
    -0.001443027, -0.00162615, -0.0018058, -0.001874155, -0.001867836, 
    -0.00186426, -0.001714303, -0.001526019, -0.001335007, -0.001172625, 
    -0.001039623, -0.0009310965, -0.0007672078, -0.0007614372, -0.0007015275, 
    -0.000523111, -0.0002745406, -3.617184e-05, 0.0002702412, 0.0005721721, 
    0.0008755261, 0.001209356, 0.00159006, 0.001970237, 0.00217691, 
    0.002310349, 0.002453003, 0.002360879, 0.00217597, 0.001995289, 
    0.001650239, 0.001085516, 0.0005262209, 6.019531e-06, -0.0006409651, 
    -0.001284812, -0.001833746, -0.002317223, -0.002841192, -0.00306009, 
    -0.003195914, -0.003794209, -0.004330654, -0.005362791, -0.007036764, 
    -0.008712401, -0.01064164, -0.01185996, -0.01542975, -0.01952004, 
    -0.009760018,
  -0.002950786, -0.002818362, -0.002853931, -0.002858099, -0.002832587, 
    -0.002847656, -0.002927176, -0.003035146, -0.003040297, -0.002924391, 
    -0.002803462, -0.002596319, -0.002418596, -0.002264529, -0.002142236, 
    -0.002040793, -0.00195953, -0.001778753, -0.001780367, -0.001738314, 
    -0.001566634, -0.001304328, -0.001050252, -0.0006711037, -0.0002595938, 
    0.000153086, 0.0006149783, 0.00114816, 0.001680912, 0.002034767, 
    0.002324915, 0.002622538, 0.002635715, 0.002543996, 0.002418877, 
    0.002118276, 0.001593073, 0.001065608, 0.0004983961, -0.0002315137, 
    -0.0009633388, -0.00165501, -0.002329998, -0.003030783, -0.00346088, 
    -0.003874376, -0.004600991, -0.005641152, -0.006894052, -0.008919518, 
    -0.01097187, -0.01264956, -0.01420295, -0.01761262, -0.01949492, 
    -0.00974746,
  -0.005432389, -0.005300641, -0.00526894, -0.005154851, -0.004984715, 
    -0.00485641, -0.004838049, -0.004881436, -0.004833595, -0.004608055, 
    -0.004368598, -0.004102294, -0.003936378, -0.00382583, -0.003756349, 
    -0.003701191, -0.003692364, -0.003601686, -0.00374505, -0.003787879, 
    -0.003613141, -0.00331009, -0.003025181, -0.002576129, -0.002123797, 
    -0.001685222, -0.001092858, -0.000336739, 0.0004192497, 0.0009855443, 
    0.001499379, 0.002002165, 0.002149514, 0.002167941, 0.002217332, 
    0.002023207, 0.001571, 0.001117016, 0.0005466651, -0.000209047, 
    -0.0009662443, -0.00173632, -0.002537876, -0.003359891, -0.004016005, 
    -0.004744666, -0.005913174, -0.007109403, -0.008626545, -0.01104471, 
    -0.01338513, -0.0155003, -0.01705705, -0.01767022, -0.02033209, 
    -0.01016604,
  -0.008399032, -0.008269353, -0.008191363, -0.008003925, -0.007765041, 
    -0.007555981, -0.00741027, -0.007348787, -0.007248223, -0.006925149, 
    -0.006582255, -0.006263497, -0.006103777, -0.006022583, -0.00600778, 
    -0.006018837, -0.006097991, -0.006096958, -0.006406454, -0.006570059, 
    -0.006424189, -0.00610286, -0.00580793, -0.005293095, -0.004802877, 
    -0.00434822, -0.003618663, -0.002610018, -0.001601015, -0.0007908734, 
    -1.499145e-05, 0.000724919, 0.001037243, 0.001176334, 0.001380479, 
    0.001325973, 0.0009897805, 0.0006433782, 9.459139e-05, -0.0006669037, 
    -0.001436563, -0.002288288, -0.003229878, -0.004170954, -0.004984145, 
    -0.005855672, -0.00742832, -0.008788267, -0.01094545, -0.01420312, 
    -0.01713342, -0.0191236, -0.01726171, -0.01902674, -0.02253933, 
    -0.01126966,
  -0.01176244, -0.01161271, -0.01152318, -0.01134062, -0.01110589, 
    -0.0108233, -0.01061728, -0.01047203, -0.01033764, -0.009965701, 
    -0.009578555, -0.009259418, -0.009127175, -0.009055188, -0.009108079, 
    -0.009254743, -0.009453665, -0.009465865, -0.009876939, -0.01017606, 
    -0.01015325, -0.009911359, -0.00968973, -0.009107583, -0.008443597, 
    -0.007913499, -0.007031781, -0.00574765, -0.004462605, -0.003381104, 
    -0.002302503, -0.001284298, -0.0007588297, -0.0004779754, -0.0001038305, 
    8.786312e-06, -0.0001958851, -0.0004195879, -0.0009139039, -0.001648763, 
    -0.002402588, -0.0033056, -0.004346755, -0.00535681, -0.006330686, 
    -0.007473555, -0.009251929, -0.01118511, -0.01406131, -0.01835002, 
    -0.02129914, -0.02041313, -0.0185816, -0.02121415, -0.02550717, 
    -0.01275358,
  -0.01458343, -0.01439012, -0.0143041, -0.01413769, -0.01392778, 
    -0.01361381, -0.01336382, -0.01316623, -0.01305114, -0.01266516, 
    -0.01226486, -0.01199156, -0.01195471, -0.01197813, -0.01219993, 
    -0.01258628, -0.01302901, -0.01320572, -0.01392911, -0.0145345, 
    -0.0147336, -0.01464175, -0.01457182, -0.01400205, -0.01330436, 
    -0.01264992, -0.01157872, -0.01001668, -0.008453965, -0.007091896, 
    -0.005658033, -0.004269951, -0.003381635, -0.00286746, -0.002306618, 
    -0.002012613, -0.002098844, -0.00220921, -0.002616095, -0.00329729, 
    -0.004018614, -0.004956169, -0.006076508, -0.00713581, -0.008223999, 
    -0.00966038, -0.01158993, -0.01433107, -0.0181261, -0.0230152, 
    -0.0234799, -0.02201523, -0.02099263, -0.02568503, -0.03087651, 
    -0.01543826,
  -0.01653155, -0.0162721, -0.01618899, -0.01604776, -0.01588372, 
    -0.01555413, -0.01525727, -0.01498682, -0.01489389, -0.01451014, 
    -0.0141191, -0.01392208, -0.01399867, -0.01411321, -0.0145321, 
    -0.01523186, -0.01597421, -0.01632821, -0.01741098, -0.01840981, 
    -0.01895291, -0.0191343, -0.01933222, -0.01885426, -0.01815331, 
    -0.01750522, -0.01636775, -0.01457382, -0.01277893, -0.01120798, 
    -0.00945488, -0.007756171, -0.006632057, -0.005944004, -0.005180239, 
    -0.004746586, -0.004834935, -0.004941361, -0.005255961, -0.005862625, 
    -0.006499368, -0.007441981, -0.008612568, -0.009717661, -0.01087449, 
    -0.01265245, -0.01514628, -0.01845619, -0.0227043, -0.02595203, 
    -0.02557703, -0.02526267, -0.02590621, -0.03133323, -0.03515927, 
    -0.01757964,
  -0.01756562, -0.0172327, -0.01714664, -0.01701301, -0.01687372, 
    -0.01650615, -0.01614727, -0.01579008, -0.01570112, -0.01528317, 
    -0.01486666, -0.01472728, -0.01489755, -0.01507435, -0.01568482, 
    -0.01672369, -0.0177812, -0.01830729, -0.0197737, -0.02121146, 
    -0.02218066, -0.02273118, -0.02328865, -0.02296841, -0.02229135, 
    -0.02166413, -0.02052343, -0.01856711, -0.01660989, -0.01491762, 
    -0.01287574, -0.01088008, -0.009586629, -0.008785347, -0.007922545, 
    -0.007484693, -0.007735183, -0.008001192, -0.008370739, -0.009099045, 
    -0.009875535, -0.01085813, -0.01208922, -0.01327974, -0.01448334, 
    -0.01661208, -0.01971501, -0.02295083, -0.02581351, -0.02860464, 
    -0.02969206, -0.03034728, -0.03180045, -0.03704233, -0.04240381, 
    -0.0212019,
  -0.01779038, -0.01738815, -0.01725632, -0.01706342, -0.01688528, 
    -0.01649473, -0.01611283, -0.0157257, -0.01560032, -0.01504978, 
    -0.01450738, -0.01435033, -0.01455149, -0.01473515, -0.01549471, 
    -0.01684, -0.01818286, -0.01886801, -0.02073154, -0.02261288, 
    -0.02403327, -0.02500037, -0.02596579, -0.0258464, -0.025243, 
    -0.02467851, -0.02359756, -0.0215508, -0.01950338, -0.01776804, 
    -0.0154543, -0.01316899, -0.01177934, -0.01085331, -0.00988624, 
    -0.009548984, -0.01009919, -0.01065822, -0.01124371, -0.01226187, 
    -0.01333706, -0.01456426, -0.01591799, -0.01724554, -0.01852608, 
    -0.02087371, -0.02412828, -0.02591742, -0.02865508, -0.03342839, 
    -0.03522338, -0.03620924, -0.03847112, -0.04459344, -0.04852627, 
    -0.02426313,
  -0.01734996, -0.01677058, -0.01650878, -0.01617595, -0.01586863, 
    -0.01522736, -0.01457735, -0.01385594, -0.0135846, -0.01308097, 
    -0.01258689, -0.01246651, -0.01263043, -0.01274826, -0.01354618, 
    -0.01504849, -0.01651815, -0.01721475, -0.01917868, -0.02121823, 
    -0.02289878, -0.02416024, -0.02540819, -0.02550809, -0.02504779, 
    -0.02460507, -0.02375349, -0.02196812, -0.02018177, -0.01872121, 
    -0.01642609, -0.0141426, -0.01283219, -0.01187147, -0.01087696, 
    -0.0107309, -0.01159905, -0.01246187, -0.01332967, -0.01466583, 
    -0.01603157, -0.01741825, -0.0188353, -0.02026976, -0.02159525, 
    -0.02385167, -0.02651836, -0.02933141, -0.03332462, -0.03943283, 
    -0.04099134, -0.04388175, -0.04629406, -0.05060396, -0.05342625, 
    -0.02671312,
  -0.01772479, -0.01693521, -0.01644392, -0.01571845, -0.01501347, 
    -0.01401404, -0.01301939, -0.01200087, -0.01147179, -0.01083471, 
    -0.01020957, -0.0101191, -0.01048016, -0.01082572, -0.01187834, 
    -0.01363828, -0.01539286, -0.01639439, -0.01860094, -0.0208197, 
    -0.02255381, -0.02380153, -0.02504969, -0.02520961, -0.02487114, 
    -0.02453333, -0.02369048, -0.02183376, -0.01997741, -0.01843041, 
    -0.01612582, -0.01381599, -0.01251574, -0.0116056, -0.01071961, 
    -0.01069607, -0.01178977, -0.01289933, -0.01407529, -0.01579538, 
    -0.01759524, -0.01947297, -0.0213718, -0.02321159, -0.02484338, 
    -0.0276447, -0.03117156, -0.03401501, -0.03956896, -0.04512876, 
    -0.05049801, -0.05246136, -0.05255504, -0.05545008, -0.05658286, 
    -0.02829143,
  -0.01836369, -0.01738496, -0.01681421, -0.01590475, -0.01499597, 
    -0.01389872, -0.01285621, -0.01181595, -0.01124129, -0.01052647, 
    -0.009810916, -0.009798326, -0.01033636, -0.01088201, -0.01219444, 
    -0.0142681, -0.01635421, -0.01760926, -0.02006609, -0.02249746, 
    -0.02429291, -0.02548237, -0.02667868, -0.02666862, -0.02623423, 
    -0.02580024, -0.0249877, -0.02320372, -0.02141924, -0.02005534, 
    -0.01783661, -0.01563708, -0.01470559, -0.01412266, -0.01353038, 
    -0.01364191, -0.01490152, -0.01617117, -0.01755309, -0.01981726, 
    -0.02213232, -0.0243354, -0.02632719, -0.02825623, -0.03002127, 
    -0.03310093, -0.03709323, -0.04049384, -0.04783232, -0.05757898, 
    -0.05994023, -0.05939956, -0.05642529, -0.05630662, -0.05658286, 
    -0.02829143,
  -0.0194362, -0.01829494, -0.01773357, -0.01677342, -0.01580735, 
    -0.01466058, -0.01357812, -0.0125013, -0.011985, -0.01122462, 
    -0.01046307, -0.01052341, -0.01125261, -0.01199368, -0.01360865, 
    -0.01608869, -0.01858381, -0.02015459, -0.02314526, -0.02610737, 
    -0.02829031, -0.02973119, -0.03117836, -0.03105103, -0.03044649, 
    -0.0298529, -0.02886337, -0.02686324, -0.02486317, -0.02342522, 
    -0.02117014, -0.01893754, -0.01808918, -0.01768821, -0.01726603, 
    -0.01788948, -0.01969323, -0.02150504, -0.02321768, -0.02572007, 
    -0.0282586, -0.03053179, -0.03269213, -0.03499031, -0.03739835, 
    -0.04162931, -0.04741015, -0.05325287, -0.06075946, -0.06805205, 
    -0.06567291, -0.06105821, -0.05642529, -0.05630662, -0.05658286, 
    -0.02829143,
  -0.02066245, -0.01941263, -0.01893786, -0.01804687, -0.01715242, 
    -0.01606033, -0.01505893, -0.01406259, -0.01368481, -0.0128512, 
    -0.01201664, -0.01217852, -0.0131969, -0.01422254, -0.01629631, 
    -0.01941303, -0.02253854, -0.02458083, -0.02853861, -0.03247919, 
    -0.03552177, -0.03768793, -0.03985658, -0.03955393, -0.03855268, 
    -0.03751893, -0.03575277, -0.03275124, -0.02974973, -0.02714372, 
    -0.0234003, -0.0196567, -0.01766573, -0.01621798, -0.01477043, 
    -0.01569494, -0.01848387, -0.02127272, -0.02450894, -0.02842406, 
    -0.03233904, -0.03668452, -0.04146057, -0.04623676, -0.0503104, 
    -0.05479553, -0.05927774, -0.06202606, -0.06552998, -0.06902567, 
    -0.06567291, -0.06105821, -0.05642529, -0.05630662, -0.05658286, 
    -0.02829143,
  -0.001369803, -0.001470851, -0.001667305, -0.001955943, -0.002290061, 
    -0.002524431, -0.002627004, -0.002802501, -0.003188644, -0.003555028, 
    -0.003908563, -0.003901996, -0.003557956, -0.003255426, -0.002998062, 
    -0.002758401, -0.002537632, -0.002380978, -0.002313672, -0.002211668, 
    -0.002085392, -0.001956344, -0.001832868, -0.001747799, -0.001680773, 
    -0.001621158, -0.001594196, -0.001528397, -0.001462683, -0.001435909, 
    -0.001403663, -0.001369967, -0.001245804, -0.001144869, -0.001069219, 
    -0.001021747, -0.001020785, -0.001003454, -0.00110317, -0.001368602, 
    -0.001725698, -0.001960843, -0.001871611, -0.001523043, -0.001389241, 
    -0.001184627, -0.0003844813, 0.0002598934, 0.001123349, 0.001861701, 
    0.002534999, 0.00304923, 0.002909161, 0.002518567, 0.001825208, 
    0.0009126041,
  -0.0006358178, -0.0005863469, -0.0007954627, -0.001055259, -0.001393613, 
    -0.001860413, -0.002425019, -0.003055943, -0.003548527, -0.00398837, 
    -0.00440433, -0.004400879, -0.00409643, -0.003768921, -0.003440062, 
    -0.003130263, -0.00281267, -0.002477895, -0.002307243, -0.002151428, 
    -0.002013475, -0.001876716, -0.001736768, -0.001662139, -0.001543778, 
    -0.001412557, -0.001353497, -0.00128625, -0.00121936, -0.001192118, 
    -0.0011579, -0.001109484, -0.001006047, -0.0009377975, -0.0008855203, 
    -0.0009983539, -0.001369843, -0.001736796, -0.001955161, -0.002227525, 
    -0.002477343, -0.002339258, -0.001898175, -0.001545541, -0.001257094, 
    -0.0007838986, -0.0001747655, 0.0008404907, 0.001088416, 0.002107221, 
    0.002819658, 0.003256213, 0.002907059, 0.00229734, 0.00130552, 
    0.0006527598,
  -0.0006509876, -0.0006022028, -0.0008165505, -0.001056557, -0.001294138, 
    -0.001733373, -0.002360168, -0.002974428, -0.003408016, -0.003808955, 
    -0.004216604, -0.004217113, -0.003909636, -0.003593609, -0.003283886, 
    -0.002980833, -0.002670638, -0.00234061, -0.002150157, -0.001973622, 
    -0.001822575, -0.001677942, -0.001529318, -0.001442904, -0.001309467, 
    -0.001161714, -0.001093936, -0.001024935, -0.0009563458, -0.0009298934, 
    -0.0009011924, -0.0008561626, -0.0007594554, -0.000705887, -0.0006768483, 
    -0.0007913178, -0.001140935, -0.001486397, -0.001684798, -0.001930325, 
    -0.002155209, -0.002079803, -0.001754775, -0.001431635, -0.001019546, 
    -0.0005433733, 0.0002405907, 0.0009743027, 0.001273688, 0.002413123, 
    0.003084044, 0.003253978, 0.002787802, 0.002108013, 0.0008606, 0.0004303,
  -0.0006622649, -0.0006144542, -0.0008313825, -0.001074553, -0.001317552, 
    -0.001736784, -0.002313664, -0.002873583, -0.003259619, -0.003623278, 
    -0.0039949, -0.003987875, -0.003705781, -0.003412461, -0.003118141, 
    -0.00282395, -0.002521117, -0.002189878, -0.00198158, -0.001790575, 
    -0.0016262, -0.001470881, -0.001312294, -0.00121397, -0.001072571, 
    -0.0009179889, -0.000845618, -0.0007741778, -0.0007031171, -0.0006775006, 
    -0.0006548314, -0.0006171229, -0.0005348113, -0.0005189425, 
    -0.0005281561, -0.0006458632, -0.0009707725, -0.001294605, -0.001475801, 
    -0.001696411, -0.001895143, -0.001818054, -0.001478318, -0.001148821, 
    -0.0007656739, -0.0002931971, 0.0006735816, 0.0009148791, 0.00143293, 
    0.002676087, 0.003311366, 0.003230323, 0.002592912, 0.001776818, 
    0.0004774586, 0.0002387293,
  -0.000670133, -0.000623758, -0.0008410701, -0.001083191, -0.001325163, 
    -0.001719526, -0.002246535, -0.002757845, -0.003102073, -0.003428577, 
    -0.003762448, -0.003747618, -0.003494477, -0.00323094, -0.002956594, 
    -0.002672488, -0.002380379, -0.002055023, -0.001834746, -0.001632308, 
    -0.001457273, -0.001292628, -0.001124645, -0.001017292, -0.0008749875, 
    -0.0007242759, -0.0006553006, -0.0005857777, -0.0005164317, 
    -0.0004965932, -0.0004859897, -0.0004676755, -0.0004175811, 
    -0.0004324816, -0.0004625981, -0.0005788199, -0.0008841287, -0.001188437, 
    -0.001342338, -0.001522156, -0.001681726, -0.001583172, -0.001238683, 
    -0.0009098395, -0.0005297249, 3.961848e-05, 0.0009928079, 0.000863364, 
    0.001570995, 0.002904117, 0.003508533, 0.003209799, 0.002423752, 
    0.001457752, 1.604535e-05, 8.022677e-06,
  -0.0006640318, -0.0006186344, -0.0008347688, -0.001076775, -0.001322203, 
    -0.001697522, -0.00217633, -0.002635383, -0.002938078, -0.003234288, 
    -0.003538539, -0.003519428, -0.003290818, -0.003049972, -0.002793405, 
    -0.002522604, -0.002243364, -0.001925984, -0.001701583, -0.00149468, 
    -0.001315314, -0.001147668, -0.0009769176, -0.0008661687, -0.0007231251, 
    -0.0005722665, -0.0005058385, -0.0004413309, -0.0003769876, 
    -0.0003649846, -0.0003658204, -0.000359484, -0.0003222262, -0.0003565548, 
    -0.0004050272, -0.0005199448, -0.0008080413, -0.001095204, -0.001225135, 
    -0.00136913, -0.001520009, -0.00143462, -0.00109869, -0.0007388291, 
    -0.0003059641, 0.0003318982, 0.0009392396, 0.0009164239, 0.001735358, 
    0.003108406, 0.003651449, 0.003191758, 0.002274991, 0.001177013, 
    -0.001063457, -0.0005317287,
  -0.0006438963, -0.0006006805, -0.000814137, -0.001050515, -0.001290087, 
    -0.001641645, -0.00207724, -0.002494423, -0.002762871, -0.003030143, 
    -0.003304907, -0.00328305, -0.003082351, -0.002870246, -0.002635509, 
    -0.002379529, -0.002115681, -0.001809649, -0.001582435, -0.001371538, 
    -0.001188297, -0.001017964, -0.0008447376, -0.0007309502, -0.0005872452, 
    -0.0004362547, -0.000375616, -0.0003154961, -0.0002551997, -0.0002517818, 
    -0.0002682353, -0.0002903033, -0.0003017313, -0.0004020739, -0.000505364, 
    -0.000626148, -0.0008905654, -0.001159288, -0.00126871, -0.001387944, 
    -0.001495676, -0.001366199, -0.0009871449, -0.0005858109, -0.000105744, 
    0.0004747299, 0.0008913045, 0.001022825, 0.00191153, 0.003295108, 
    0.003609697, 0.003035848, 0.002115142, 0.0009253444, -0.002031629, 
    -0.001015814,
  -0.0006254187, -0.000584205, -0.000795204, -0.001026416, -0.001260616, 
    -0.001590369, -0.001986308, -0.002365071, -0.002602091, -0.002842808, 
    -0.003090513, -0.003066135, -0.00289105, -0.002705318, -0.002489597, 
    -0.002246963, -0.001995327, -0.001697069, -0.001470455, -0.00126383, 
    -0.001083314, -0.000914272, -0.0007420224, -0.0006315213, -0.0005039392, 
    -0.0003767879, -0.0003330927, -0.0002884126, -0.0002435682, 
    -0.0002593976, -0.0002974757, -0.0003407784, -0.0003699293, 
    -0.0004925178, -0.0006178659, -0.0007388186, -0.0009913502, -0.001247892, 
    -0.001328152, -0.001406116, -0.001473346, -0.001303411, -0.0008847807, 
    -0.0004679629, -3.108172e-05, 0.0004334769, 0.0008473126, 0.00112048, 
    0.002073233, 0.003466502, 0.003571361, 0.002806367, 0.001823726, 
    0.0003669162, -0.00292187, -0.001460935,
  -0.0005428722, -0.0005006843, -0.0007056151, -0.0009350374, -0.001174559, 
    -0.00149053, -0.00184154, -0.002168387, -0.002371418, -0.002595076, 
    -0.002826676, -0.00280699, -0.002656946, -0.002492856, -0.00230058, 
    -0.002082422, -0.001855872, -0.001578827, -0.001362431, -0.001164672, 
    -0.0009918627, -0.0008303584, -0.000665863, -0.0005623291, -0.0004433219, 
    -0.0003247088, -0.000292831, -0.0002627696, -0.0002325553, -0.0002666083, 
    -0.0003251609, -0.0003885691, -0.0004345006, -0.0005781521, 
    -0.0007243855, -0.0008454978, -0.001086776, -0.001331784, -0.001384432, 
    -0.001423321, -0.001469615, -0.001309113, -0.0009197519, -0.0005059934, 
    -6.388787e-05, 0.0003944166, 0.0008664925, 0.001212949, 0.002226362, 
    0.003628823, 0.00353505, 0.002588969, 0.001547587, -0.0007348852, 
    -0.003765916, -0.001882958,
  -0.0004494184, -0.0004083927, -0.0006066324, -0.0008250108, -0.001052767, 
    -0.001345577, -0.001660308, -0.00195261, -0.002130531, -0.002334746, 
    -0.002546333, -0.002531207, -0.002411958, -0.002279666, -0.002115362, 
    -0.001921188, -0.00171922, -0.001462962, -0.001256579, -0.001067507, 
    -0.0009022495, -0.0007481311, -0.0005912342, -0.0004945273, 
    -0.0003839226, -0.0002736762, -0.0002535653, -0.0002380071, 
    -0.0002222192, -0.0002746169, -0.0003547033, -0.0004429047, 
    -0.0005183401, -0.00070294, -0.0008893555, -0.001020161, -0.001257577, 
    -0.001500081, -0.001537247, -0.00156461, -0.001594162, -0.001405787, 
    -0.0009858368, -0.00054326, -9.60351e-05, 0.0003561408, 0.0009134181, 
    0.001322988, 0.002374667, 0.003787896, 0.003499463, 0.002375894, 
    0.001276914, -0.001815003, -0.004551867, -0.002275933,
  -0.000353054, -0.0003114062, -0.0005026633, -0.0007136743, -0.0009295259, 
    -0.001198897, -0.001476917, -0.001734264, -0.001884866, -0.002071318, 
    -0.002262653, -0.002252141, -0.002164053, -0.00205486, -0.00191033, 
    -0.001741156, -0.001560204, -0.001313219, -0.001110597, -0.0009353741, 
    -0.0007872758, -0.0006480207, -0.0005047102, -0.000418251, -0.0003183075, 
    -0.0002205657, -0.0002181777, -0.0002228234, -0.0002272576, 
    -0.0003069323, -0.0004164631, -0.0005334576, -0.0006359931, 
    -0.0008516116, -0.001068916, -0.001208377, -0.001449363, -0.001695029, 
    -0.001711848, -0.001715016, -0.001720193, -0.001503612, -0.001052708, 
    -0.00058097, -0.0001210127, 0.0003835233, 0.0009609018, 0.001446865, 
    0.002517444, 0.003713343, 0.003304671, 0.00216031, 0.001003068, 
    -0.002907708, -0.005302904, -0.002651452,
  -0.0001554013, -0.0001083631, -0.0002814345, -0.0004736518, -0.0006824963, 
    -0.0009323499, -0.00116345, -0.001366211, -0.0014882, -0.001662145, 
    -0.001844229, -0.001845769, -0.001787154, -0.001710482, -0.001603019, 
    -0.00146985, -0.001325937, -0.001111788, -0.0009349378, -0.0007830836, 
    -0.0006541747, -0.000531528, -0.0004051809, -0.0003329885, -0.0002482244, 
    -0.0001654579, -0.0001815139, -0.0002070921, -0.0002324777, 
    -0.0003404131, -0.0004804499, -0.0006272757, -0.0007578884, -0.001005644, 
    -0.001254951, -0.00140338, -0.001648063, -0.001897006, -0.001892743, 
    -0.001870846, -0.001840623, -0.001588338, -0.001117112, -0.0006482811, 
    -0.0001136096, 0.0004149337, 0.0010153, 0.001575202, 0.002665355, 
    0.003612873, 0.002920385, 0.001642654, -6.525819e-05, -0.003999529, 
    -0.006080324, -0.003040162,
  5.202551e-05, 0.0001041108, -4.993028e-05, -0.0002166163, -0.0003982502, 
    -0.0006156968, -0.0008073315, -0.0009734943, -0.001073111, -0.001231192, 
    -0.001396588, -0.001408439, -0.001387391, -0.001350108, -0.001281433, 
    -0.001185943, -0.001080789, -0.0009010013, -0.0007489508, -0.0006189908, 
    -0.0005120439, -0.0004092258, -0.0003010292, -0.0002437661, 
    -0.0001638519, -7.779587e-05, -9.946213e-05, -0.0001399011, 
    -0.0001805262, -0.0003108478, -0.0004719404, -0.000627339, -0.0007508434, 
    -0.0009878086, -0.0012375, -0.001393163, -0.00166417, -0.001933936, 
    -0.001922868, -0.001900918, -0.001882633, -0.001642625, -0.001181543, 
    -0.0007226259, -0.0001058629, 0.0004478018, 0.001107022, 0.001704773, 
    0.002820116, 0.003507759, 0.002518378, 0.001100739, -0.001525236, 
    -0.004834577, -0.006926587, -0.003463293,
  0.0001891807, 0.0002523046, 0.0001336798, 1.352876e-05, -0.0001211187, 
    -0.0002945779, -0.0004393437, -0.0005600958, -0.0006323452, 
    -0.0007701878, -0.0009151315, -0.0009338554, -0.0009449744, 
    -0.0009386512, -0.0009038303, -0.0008470276, -0.0007795909, 
    -0.0006248979, -0.000499265, -0.0003988662, -0.0003114804, -0.0002204205, 
    -0.0001259986, -6.940928e-05, 1.094897e-05, 9.629846e-05, 7.410551e-05, 
    3.42911e-05, -5.687998e-06, -0.0001480438, -0.0003240963, -0.0004951078, 
    -0.0006447743, -0.0009142314, -0.001194935, -0.001363907, -0.001654518, 
    -0.001944027, -0.001936279, -0.0019297, -0.001926337, -0.001699102, 
    -0.001239186, -0.0007700328, -8.913255e-05, 0.0005132961, 0.001202442, 
    0.001804382, 0.002707472, 0.003134249, 0.002003851, 0.0005371741, 
    -0.003043292, -0.00570267, -0.008698069, -0.004349034,
  0.0002782255, 0.0003598106, 0.0002864538, 0.0002200317, 0.0001410702, 
    2.163237e-05, -6.713378e-05, -0.0001351339, -0.0001775135, -0.0002915361, 
    -0.0004116987, -0.0004333507, -0.0004743129, -0.0005001865, 
    -0.0005017992, -0.0004847905, -0.0004585789, -0.0003369398, 
    -0.0002448276, -0.0001745525, -0.0001071001, -2.802207e-05, 5.396692e-05, 
    0.0001087725, 0.0001890763, 0.000266248, 0.0002498213, 0.0002211568, 
    0.0001918575, 4.750862e-05, -0.0001298826, -0.0002896087, -0.0004199546, 
    -0.0006611147, -0.0009199351, -0.001089768, -0.00141266, -0.001728486, 
    -0.001733187, -0.001748448, -0.001762623, -0.001547986, -0.001118034, 
    -0.000712286, -6.041183e-05, 0.000581998, 0.001255004, 0.001905884, 
    0.002487061, 0.002447083, 0.001029703, -0.001239472, -0.004277576, 
    -0.007160407, -0.01050249, -0.005251244,
  -0.0001237267, -2.871204e-05, -3.657124e-05, 6.623475e-07, 4.214035e-05, 
    1.66769e-05, -1.731322e-05, -5.05129e-05, -6.589659e-05, -0.0001304441, 
    -0.000196716, -0.0002014703, -0.0002677826, -0.000333138, -0.0003730627, 
    -0.000388067, -0.0004041579, -0.0003266924, -0.0002872311, -0.0002466516, 
    -0.0001737696, -7.245308e-05, 2.754815e-05, 0.0001196148, 0.0002404165, 
    0.0003718454, 0.0004168911, 0.0004577434, 0.0004980584, 0.0004047227, 
    0.000274651, 0.0001595214, 3.805571e-05, -0.0002044422, -0.0004618814, 
    -0.0006346463, -0.0009775107, -0.001314398, -0.001358997, -0.001435833, 
    -0.001511728, -0.001362148, -0.001000356, -0.0006693766, -6.490888e-05, 
    0.0005824754, 0.001264391, 0.001662032, 0.001991262, 0.001616508, 
    4.632342e-05, -0.003087682, -0.005387079, -0.009182463, -0.01273331, 
    -0.006366655,
  -0.0007868812, -0.0006671366, -0.000602355, -0.000482206, -0.0003585742, 
    -0.0003030218, -0.0002469947, -0.0001902887, -0.0001529492, 
    -0.0001692426, -0.0001869667, -0.00017008, -0.0002385852, -0.0003062745, 
    -0.000359852, -0.0003997525, -0.0004659549, -0.0004775156, -0.0005435845, 
    -0.0005513128, -0.000454932, -0.000306464, -0.0001694257, -3.514235e-05, 
    9.404857e-05, 0.0002306601, 0.0003403502, 0.0004872925, 0.0006335743, 
    0.0006220855, 0.0005689189, 0.0005267434, 0.000433983, 0.0002184499, 
    6.319065e-07, -0.0001589649, -0.0005132584, -0.0008621579, -0.0009548798, 
    -0.001104776, -0.001255324, -0.001192931, -0.0009323871, -0.0006965343, 
    -0.0001369274, 0.0005537063, 0.0009773619, 0.001302616, 0.001089698, 
    0.0002072371, -0.00202851, -0.004993218, -0.007558343, -0.01153942, 
    -0.01472131, -0.007360656,
  -0.002714143, -0.002597664, -0.002452021, -0.002192347, -0.001903237, 
    -0.001711161, -0.001571477, -0.001462275, -0.001385905, -0.001311139, 
    -0.001230171, -0.001160014, -0.001233001, -0.00133188, -0.001420247, 
    -0.001486312, -0.001574094, -0.001557467, -0.001623422, -0.00164231, 
    -0.001537914, -0.001352206, -0.001175722, -0.0009405029, -0.0006721035, 
    -0.0003976931, -0.000140712, 0.0001695988, 0.0004793733, 0.000605667, 
    0.0006877517, 0.0007787413, 0.0007558869, 0.0005963717, 0.0004009498, 
    0.0002568596, -9.026098e-05, -0.0004390203, -0.000591167, -0.0008348616, 
    -0.001087988, -0.001157077, -0.001052641, -0.0009614375, -0.0005165954, 
    4.705341e-05, 0.000484974, 0.0002803023, -0.0002688241, -0.001615791, 
    -0.004275209, -0.007225301, -0.01002891, -0.01352483, -0.01489312, 
    -0.007446561,
  -0.005173279, -0.005070079, -0.004858568, -0.004476597, -0.004039468, 
    -0.003717734, -0.003494687, -0.003333973, -0.003227662, -0.003061595, 
    -0.002880685, -0.002757769, -0.002841537, -0.002983063, -0.003124437, 
    -0.003237474, -0.003398942, -0.003468317, -0.003678023, -0.003782829, 
    -0.003662008, -0.003409507, -0.003176572, -0.002834935, -0.002482749, 
    -0.002137214, -0.001711963, -0.001151166, -0.0005907044, -0.0002527087, 
    3.401206e-05, 0.0003128677, 0.000383126, 0.000290849, 0.0002217928, 
    0.0001382219, -0.0001848655, -0.0005092376, -0.0006974244, -0.001001121, 
    -0.001312259, -0.001455636, -0.001439587, -0.001434042, -0.001124596, 
    -0.0007519118, -0.0006972533, -0.001026749, -0.001944555, -0.003782823, 
    -0.006899771, -0.01034912, -0.01269716, -0.01351754, -0.01629313, 
    -0.008146564,
  -0.008129088, -0.008044805, -0.007786204, -0.007319318, -0.006802484, 
    -0.006408796, -0.006066101, -0.00580753, -0.005670496, -0.005424038, 
    -0.005157473, -0.004991009, -0.00508515, -0.005259158, -0.005460294, 
    -0.005647041, -0.005903971, -0.006062251, -0.006448059, -0.006684539, 
    -0.006585569, -0.006291175, -0.006024853, -0.005574516, -0.005130589, 
    -0.004712053, -0.004096779, -0.003238286, -0.00237981, -0.001789901, 
    -0.001257046, -0.0007545101, -0.0005634231, -0.000585155, -0.000553873, 
    -0.0005556907, -0.0008246856, -0.001102755, -0.001317057, -0.001681042, 
    -0.002062148, -0.00231955, -0.002453279, -0.002580184, -0.002320552, 
    -0.001914513, -0.002241387, -0.002708508, -0.004413663, -0.007232021, 
    -0.01091246, -0.01358707, -0.01268081, -0.01558204, -0.01965417, 
    -0.009827083,
  -0.01153912, -0.01146837, -0.01119507, -0.01070869, -0.01017078, 
    -0.009697657, -0.009278418, -0.008919118, -0.008766617, -0.008477351, 
    -0.00817266, -0.008011702, -0.008141224, -0.008332036, -0.008615073, 
    -0.008958469, -0.009355726, -0.009534927, -0.01004751, -0.01044549, 
    -0.01047642, -0.01024778, -0.01004068, -0.009469095, -0.008773987, 
    -0.00820758, -0.00736957, -0.006167251, -0.0049646, -0.004083998, 
    -0.003259709, -0.002486769, -0.00212958, -0.002067575, -0.001929464, 
    -0.001833649, -0.002049105, -0.002281384, -0.002504704, -0.002915703, 
    -0.00335841, -0.003722033, -0.003988934, -0.004221099, -0.004063562, 
    -0.003833883, -0.004274254, -0.005379568, -0.007875649, -0.01168009, 
    -0.01462323, -0.01461335, -0.01453375, -0.01897346, -0.02361541, 
    -0.01180771,
  -0.01447437, -0.01441534, -0.01414997, -0.01365136, -0.01310802, 
    -0.01258713, -0.0120907, -0.01164608, -0.01152473, -0.01120331, 
    -0.01086801, -0.0107445, -0.01095565, -0.01122563, -0.01167639, 
    -0.01227569, -0.01293123, -0.0132861, -0.01416845, -0.01493508, 
    -0.01523292, -0.01517947, -0.01514831, -0.01453535, -0.01371785, 
    -0.0129354, -0.01180361, -0.01020908, -0.008614316, -0.007408947, 
    -0.00622463, -0.005079236, -0.004425032, -0.004208575, -0.00395593, 
    -0.003760446, -0.003957969, -0.004175975, -0.004394983, -0.004849595, 
    -0.005361229, -0.005838405, -0.006243454, -0.006589283, -0.006513682, 
    -0.006503998, -0.007016363, -0.008966806, -0.01230085, -0.01588056, 
    -0.0164455, -0.01662433, -0.01815246, -0.02430748, -0.02988798, 
    -0.01494399,
  -0.01661164, -0.01655779, -0.01631814, -0.01582953, -0.0153128, 
    -0.01475602, -0.01417316, -0.01361978, -0.01352812, -0.01316782, 
    -0.01280047, -0.01272917, -0.0130077, -0.01332151, -0.01393824, 
    -0.0148384, -0.01577894, -0.01631661, -0.0176274, -0.01886158, 
    -0.01958017, -0.01987481, -0.02018465, -0.01962234, -0.0187302, 
    -0.01788585, -0.01656529, -0.01458879, -0.01261189, -0.01112191, 
    -0.009575107, -0.008073504, -0.007230861, -0.006912418, -0.006532535, 
    -0.006285474, -0.006604194, -0.006938248, -0.007179629, -0.007702169, 
    -0.008267458, -0.008857405, -0.009399438, -0.009887693, -0.009872314, 
    -0.01013691, -0.01119347, -0.01351675, -0.01640612, -0.01841681, 
    -0.01893319, -0.02126792, -0.02392302, -0.03055274, -0.03489117, 
    -0.01744559,
  -0.01786526, -0.01782172, -0.01762415, -0.01714151, -0.01664727, 
    -0.01603962, -0.01535109, -0.01466813, -0.01458052, -0.01413944, 
    -0.01369963, -0.01365739, -0.01395566, -0.01425775, -0.01500621, 
    -0.01620037, -0.01740968, -0.01812638, -0.01989805, -0.02165087, 
    -0.02290086, -0.02369206, -0.02448731, -0.02406503, -0.02316633, 
    -0.02231932, -0.02087317, -0.0185741, -0.01627463, -0.01456276, 
    -0.01264804, -0.01077131, -0.009791846, -0.009395917, -0.008947887, 
    -0.008752846, -0.009331845, -0.009923525, -0.01033759, -0.01115678, 
    -0.0120376, -0.01281542, -0.0135382, -0.01423535, -0.0142617, 
    -0.01474706, -0.01625186, -0.01736004, -0.01926993, -0.02161445, 
    -0.02462445, -0.02767606, -0.03041776, -0.03692668, -0.04318651, 
    -0.02159326,
  -0.01814218, -0.0181119, -0.01794165, -0.017414, -0.01689964, -0.01621129, 
    -0.01536284, -0.01448925, -0.0143509, -0.01379673, -0.01325154, 
    -0.01320677, -0.01346283, -0.01369198, -0.01452143, -0.01596718, 
    -0.01740192, -0.01828239, -0.02049336, -0.02274155, -0.02455769, 
    -0.02593257, -0.02730038, -0.02710347, -0.02631073, -0.02556561, 
    -0.02409188, -0.02159523, -0.01909817, -0.0172644, -0.01502101, 
    -0.01280209, -0.01175558, -0.01126348, -0.0107349, -0.01065338, 
    -0.01156634, -0.01248687, -0.013187, -0.0144394, -0.01572962, 
    -0.01671453, -0.01750199, -0.01834395, -0.0183102, -0.01852359, 
    -0.01936872, -0.02047086, -0.02313202, -0.02832445, -0.03202217, 
    -0.03473979, -0.03790673, -0.04544931, -0.05018502, -0.02509251,
  -0.01680728, -0.01669698, -0.01642278, -0.01571215, -0.01505522, 
    -0.01424956, -0.01318671, -0.01205567, -0.01171988, -0.01102857, 
    -0.0103599, -0.01026329, -0.01040653, -0.01047216, -0.01127219, 
    -0.01284924, -0.01436986, -0.0153103, -0.01762872, -0.02007416, 
    -0.02220613, -0.02392641, -0.02562629, -0.02566609, -0.02500113, 
    -0.0243422, -0.02290359, -0.02047585, -0.01804843, -0.01626325, 
    -0.01389781, -0.01150326, -0.0103698, -0.009752079, -0.009200842, 
    -0.00931378, -0.01055777, -0.01179413, -0.01289698, -0.01471508, 
    -0.0166085, -0.01827464, -0.01966815, -0.02103049, -0.0212981, 
    -0.02189832, -0.02311102, -0.02565787, -0.02995433, -0.03699359, 
    -0.03964449, -0.04376496, -0.04679377, -0.05223314, -0.05578612, 
    -0.02789306,
  -0.01507635, -0.01485235, -0.0144259, -0.01344822, -0.01250221, 
    -0.01149134, -0.01021356, -0.008887227, -0.008353014, -0.007463353, 
    -0.006589608, -0.006362895, -0.006527869, -0.006646339, -0.007553841, 
    -0.00927236, -0.01095903, -0.0120474, -0.0145855, -0.0171994, -0.0193945, 
    -0.0211156, -0.02282642, -0.02284894, -0.02222882, -0.021584, 
    -0.02030823, -0.01802395, -0.01573994, -0.01420307, -0.01204186, 
    -0.009863566, -0.009165678, -0.009157538, -0.009192468, -0.00976638, 
    -0.01154626, -0.01335583, -0.01507968, -0.01769184, -0.02043471, 
    -0.02283098, -0.02481099, -0.02669172, -0.02724246, -0.0285014, 
    -0.0308101, -0.03301387, -0.03977935, -0.04530321, -0.05112894, 
    -0.05374107, -0.05390639, -0.05770276, -0.05938499, -0.0296925,
  -0.01353696, -0.01313822, -0.01264737, -0.01152011, -0.01041419, 
    -0.00925343, -0.007872249, -0.006464271, -0.005898115, -0.005160019, 
    -0.004424037, -0.004364876, -0.004685556, -0.004996878, -0.006069874, 
    -0.007905872, -0.009735674, -0.0110469, -0.01394778, -0.01686613, 
    -0.01937197, -0.02145613, -0.02353522, -0.0237838, -0.02348379, 
    -0.02320732, -0.02229965, -0.02029604, -0.01829117, -0.01715635, 
    -0.01534843, -0.01358175, -0.01373759, -0.01424006, -0.01471465, 
    -0.01584077, -0.01824107, -0.02066005, -0.02285515, -0.0259791, 
    -0.0291866, -0.03208698, -0.03448929, -0.0367818, -0.03737604, 
    -0.03880777, -0.041749, -0.04436039, -0.05182424, -0.0606414, 
    -0.06234463, -0.06180862, -0.0582882, -0.05865494, -0.05938499, -0.0296925,
  -0.01137528, -0.01091745, -0.0104146, -0.009225722, -0.008052643, 
    -0.006873852, -0.005551537, -0.004213117, -0.003861725, -0.003460936, 
    -0.003059977, -0.003439258, -0.004417752, -0.005412239, -0.007155619, 
    -0.009627871, -0.01212103, -0.01430577, -0.01787898, -0.02140432, 
    -0.02437397, -0.02684116, -0.02931746, -0.02986106, -0.02987777, 
    -0.02993299, -0.0293696, -0.02773819, -0.02610482, -0.02557884, 
    -0.02430847, -0.02310887, -0.02410766, -0.02534769, -0.02652519, 
    -0.02820586, -0.03110954, -0.03404226, -0.03636805, -0.03957402, 
    -0.04285251, -0.04615667, -0.04927384, -0.05225703, -0.05323664, 
    -0.05524506, -0.05936907, -0.06331872, -0.06903841, -0.07350741, 
    -0.06915011, -0.06372725, -0.0582882, -0.05865494, -0.05938499, -0.0296925,
  -0.011168, -0.01092292, -0.01082621, -0.009928421, -0.009024217, 
    -0.007804603, -0.00628587, -0.004768915, -0.004695355, -0.004333754, 
    -0.003971286, -0.004568148, -0.005759081, -0.006954384, -0.009192388, 
    -0.01247079, -0.01575695, -0.01900352, -0.02409841, -0.0291787, 
    -0.03380602, -0.03800162, -0.04219681, -0.04345107, -0.04386142, 
    -0.04422602, -0.04382206, -0.04237097, -0.04091989, -0.04092176, 
    -0.03978365, -0.03864539, -0.04029267, -0.04194067, -0.04358883, 
    -0.04623856, -0.0505375, -0.05483638, -0.0582884, -0.0626262, 
    -0.06696386, -0.07067639, -0.07376382, -0.07685139, -0.07751536, 
    -0.0778706, -0.07822324, -0.07608602, -0.07539912, -0.07470489, 
    -0.06915011, -0.06372725, -0.0582882, -0.05865494, -0.05938499, -0.0296925 ;

 v_north =
  -0.0004091309, -0.0003311469, -0.000393715, -0.00063217, -0.0007742811, 
    -0.0006616398, -0.0004406187, -0.0002988141, -0.0003778972, 
    -0.0005306175, -0.0006818859, -0.000697663, -0.0005508081, -0.0003629736, 
    1.425777e-05, 0.0001702391, 0.000283393, 0.0002407248, 0.0002349741, 
    0.0003028092, 0.0003557904, 0.0003143993, 0.0003297645, 0.0005593741, 
    0.002649494, 0.00571339, 0.008017274, 0.009916961, 0, 8.673617e-19, 
    -8.673617e-19, -1.734723e-18, 0, 1.734723e-18, 8.673617e-19, 0, 
    8.673617e-19, 0, -8.673617e-19, 0, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18,
  -0.0007257851, -0.0007227993, -0.0008222297, -0.0008791936, -0.0007857079, 
    -0.0006840323, -0.0006092073, -0.0006064775, -0.0007636705, 
    -0.0008601076, -0.0009552408, -0.0008290236, -0.0005579228, 
    -0.0002861402, 0.0001350895, 0.0002835469, 0.0004207557, 0.0004056111, 
    0.0003898476, 0.0003743869, 0.0003409325, 0.0003290634, 0.000306788, 
    0.0009690252, 0.003334302, 0.006394592, 0.008657211, 0.009945949, 0, 
    8.673617e-19, -8.673617e-19, -1.734723e-18, 0, 1.734723e-18, 
    8.673617e-19, 0, 8.673617e-19, 0, -8.673617e-19, 0, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.0009088299, -0.0009510079, -0.0009327102, -0.0008410601, -0.000741843, 
    -0.0007016098, -0.0007191743, -0.0007285398, -0.0008204354, 
    -0.0008394118, -0.0008492682, -0.0007168335, -0.000452764, -0.0001880832, 
    0.0002139107, 0.0003539751, 0.0004838053, 0.0004605078, 0.0004154943, 
    0.0003706794, 0.0003319033, 0.0003443249, 0.0002871499, 0.001319215, 
    0.003919866, 0.007094427, 0.00920508, 0.009970799, 0, 8.673617e-19, 
    -8.673617e-19, -1.734723e-18, 0, 1.734723e-18, 8.673617e-19, 0, 
    8.673617e-19, 0, -8.673617e-19, 0, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18,
  -0.0009050265, -0.0009341846, -0.0009054743, -0.0008096927, -0.0007190976, 
    -0.0006825708, -0.000689569, -0.0006890558, -0.0007588991, -0.000762099, 
    -0.0007569205, -0.0006204207, -0.0003623934, -0.0001005123, 0.0002925122, 
    0.0004323267, 0.0005558321, 0.0005209151, 0.0004463214, 0.000381254, 
    0.000347093, 0.0003584441, 0.0002702702, 0.001734966, 0.004692433, 
    0.007732151, 0.009676876, 0.01214854, 0, 8.673617e-19, -8.673617e-19, 
    -1.734723e-18, 0, 1.734723e-18, 8.673617e-19, 0, 8.673617e-19, 0, 
    -8.673617e-19, 0, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.000901702, -0.0009195466, -0.0008839237, -0.0007929376, -0.0007040417, 
    -0.0006660669, -0.0006639057, -0.000654829, -0.0007044478, -0.0006931214, 
    -0.0006754282, -0.0005330369, -0.0002703866, -2.30608e-06, 0.0003794041, 
    0.000521405, 0.0006483732, 0.0006177165, 0.000510245, 0.0004115153, 
    0.0003602608, 0.0003841696, 0.0005617571, 0.002420022, 0.005412862, 
    0.008285695, 0.01003414, 0.01425077, 0, 8.673617e-19, -8.673617e-19, 
    -1.734723e-18, 0, 1.734723e-18, 8.673617e-19, 0, 8.673617e-19, 0, 
    -8.673617e-19, 0, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.0008971078, -0.0009051768, -0.0008675726, -0.0007782234, -0.0006908196, 
    -0.0006339756, -0.0006200801, -0.000601606, -0.0006450036, -0.0006265028, 
    -0.0006021023, -0.0004544949, -0.0001877919, 8.394398e-05, 0.0004557178, 
    0.000599639, 0.0007296484, 0.0007027329, 0.0005663862, 0.0004380927, 
    0.0003718259, 0.0004067651, 0.0008733275, 0.003021934, 0.006046073, 
    0.008772504, 0.01007951, 0.01610438, 0, 8.673617e-19, -8.673617e-19, 
    -1.734723e-18, 0, 1.734723e-18, 8.673617e-19, 0, 8.673617e-19, 0, 
    -8.673617e-19, 0, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.0008929326, -0.0008923188, -0.0008529417, -0.0007486739, -0.000617757, 
    -0.0005679587, -0.0005606881, -0.0005491827, -0.0005918106, 
    -0.0005668899, -0.0005364869, -0.0003842116, -0.0001138817, 0.0001611256, 
    0.0005310484, 0.0006897062, 0.0008098641, 0.0007788109, 0.0006166248, 
    0.0004693703, 0.0004355171, 0.0004269866, 0.001152196, 0.003560784, 
    0.00661313, 0.009242048, 0.0101202, 0.01776941, 0, 8.673617e-19, 
    -8.673617e-19, -1.734723e-18, 0, 1.734723e-18, 8.673617e-19, 0, 
    8.673617e-19, 0, -8.673617e-19, 0, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18,
  -0.0008880975, -0.0008785119, -0.0008038479, -0.0006683349, -0.0005487826, 
    -0.0005073732, -0.0005061824, -0.000501072, -0.0005429934, -0.0005121807, 
    -0.0004748866, -0.0002846366, 1.877006e-05, 0.0003297773, 0.0007179913, 
    0.0008745974, 0.0009953537, 0.0009578125, 0.0007507309, 0.0005742437, 
    0.0004951952, 0.0005017522, 0.001408173, 0.004055493, 0.007177123, 
    0.009718472, 0.01015761, 0.01846175, 0, 8.673617e-19, -8.673617e-19, 
    -1.734723e-18, 0, 1.734723e-18, 8.673617e-19, 0, 8.673617e-19, 0, 
    -8.673617e-19, 0, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.0008056353, -0.0007843534, -0.0007159277, -0.0005922663, -0.000483474, 
    -0.0004500074, -0.0004521743, -0.0004053639, -0.0004145803, 
    -0.0003569463, -0.0002874974, -9.625684e-05, 0.0002060273, 0.0005153801, 
    0.0008950041, 0.001049668, 0.00117099, 0.00113938, 0.0008922476, 
    0.0006735463, 0.0005517038, 0.0008269649, 0.001849626, 0.004755252, 
    0.007809481, 0.01016993, 0.01019309, 0.01878751, 0, 8.673617e-19, 
    -8.673617e-19, -1.734723e-18, 0, 1.734723e-18, 8.673617e-19, 0, 
    8.673617e-19, 0, -8.673617e-19, 0, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18,
  -0.0007213026, -0.0006920862, -0.0006297735, -0.0005177254, -0.0003416345, 
    -0.0002665861, -0.0002520814, -0.0002176183, -0.000239478, -0.000177148, 
    -0.0001038697, 8.83418e-05, 0.0003895262, 0.000697258, 0.001068464, 
    0.001221225, 0.001343102, 0.001317304, 0.001030924, 0.0007708561, 
    0.0006070787, 0.001145657, 0.002477252, 0.005517075, 0.008429251, 
    0.01061245, 0.01140403, 0.019107, 0, 8.673617e-19, -8.673617e-19, 
    -1.734723e-18, 0, 1.734723e-18, 8.673617e-19, 0, 8.673617e-19, 0, 
    -8.673617e-19, 0, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.0006359664, -0.0005987211, -0.0005149462, -0.0003025115, -0.0001155072, 
    -5.322507e-05, -4.960873e-05, -2.763974e-05, -6.229343e-05, 4.788457e-06, 
    8.194162e-05, 0.0002751354, 0.0005752068, 0.0008812983, 0.001273525, 
    0.001438331, 0.001548763, 0.00150942, 0.001178433, 0.0009372316, 
    0.0009943112, 0.001468134, 0.003112324, 0.006287914, 0.009056329, 
    0.01106016, 0.01386148, 0.01943014, 0, 8.673617e-19, -8.673617e-19, 
    -1.734723e-18, 0, 1.734723e-18, 8.673617e-19, 0, 8.673617e-19, 0, 
    -8.673617e-19, 0, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.0003978741, -0.00034032, -0.0002312633, -4.465598e-05, 0.0001187685, 
    0.0001678238, 0.0001601592, 0.0001691833, 0.0001385505, 0.000231561, 
    0.0003391812, 0.0005624328, 0.0008872387, 0.001220401, 0.001614142, 
    0.0017789, 0.001894162, 0.001892514, 0.001585192, 0.00135962, 
    0.001396072, 0.001905498, 0.003770216, 0.007086388, 0.009706432, 
    0.01115279, 0.01640527, 0.02553676, 0, 8.673617e-19, -8.673617e-19, 
    -1.734723e-18, 0, 1.734723e-18, 8.673617e-19, 0, 8.673617e-19, 0, 
    -8.673617e-19, 0, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -9.910145e-05, -2.788076e-05, 6.558855e-05, 0.0002251678, 0.0004375819, 
    0.000526287, 0.000531889, 0.0005692688, 0.0005273267, 0.0006171745, 
    0.0007201271, 0.0009367327, 0.001254363, 0.001579484, 0.001970557, 
    0.002135265, 0.002255582, 0.002293378, 0.002010818, 0.0018016, 
    0.001816463, 0.002815442, 0.004710187, 0.008078902, 0.01047934, 
    0.01121293, 0.01898959, 0.03422154, 0, 8.673617e-19, -8.673617e-19, 
    -1.734723e-18, 0, 1.734723e-18, 8.673617e-19, 0, 8.673617e-19, 0, 
    -8.673617e-19, 0, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  0.0002478032, 0.0003431894, 0.000484763, 0.0007270293, 0.0009452706, 
    0.001015347, 0.0009983783, 0.001009393, 0.0009317743, 0.001018332, 
    0.001116428, 0.001326118, 0.001636282, 0.001963891, 0.002381845, 
    0.002569326, 0.002691833, 0.002755137, 0.002504497, 0.002407094, 
    0.00275074, 0.003762025, 0.005881221, 0.009200088, 0.01128315, 
    0.01127547, 0.01976383, 0.04324285, 0, 8.673617e-19, -8.673617e-19, 
    -1.734723e-18, 0, 1.734723e-18, 8.673617e-19, 0, 8.673617e-19, 0, 
    -8.673617e-19, 0, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  0.0008293592, 0.0009564157, 0.001078869, 0.001281123, 0.001462614, 
    0.001532767, 0.00150899, 0.001519142, 0.001420155, 0.00151394, 
    0.001621112, 0.001846358, 0.002179344, 0.002524141, 0.002961842, 
    0.00319442, 0.003370961, 0.003558046, 0.003485795, 0.003545801, 
    0.003894303, 0.004983849, 0.007074472, 0.01034305, 0.01197456, 
    0.01440581, 0.02055247, 0.04295902, 0, 8.673617e-19, -8.673617e-19, 
    -1.734723e-18, 0, 1.734723e-18, 8.673617e-19, 0, 8.673617e-19, 0, 
    -8.673617e-19, 0, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  0.001419443, 0.001583569, 0.001720193, 0.001942741, 0.002149284, 
    0.002216302, 0.002161761, 0.002135807, 0.001983383, 0.002070286, 
    0.002168467, 0.002390922, 0.002728946, 0.003076922, 0.003536056, 
    0.003819517, 0.004049717, 0.004351384, 0.004454012, 0.004714403, 
    0.0053056, 0.006510374, 0.008527997, 0.01157706, 0.01234232, 0.01793243, 
    0.03573227, 0.04203144, 0, 8.673617e-19, -8.673617e-19, -1.734723e-18, 0, 
    1.734723e-18, 8.673617e-19, 0, 8.673617e-19, 0, -8.673617e-19, 0, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  0.002111342, 0.002328543, 0.002454122, 0.002639377, 0.002812759, 
    0.002866994, 0.002779146, 0.002711602, 0.002491637, 0.002568451, 
    0.002653435, 0.002876026, 0.003232527, 0.0036004, 0.004107421, 
    0.004479611, 0.004807959, 0.005314863, 0.005755627, 0.006334029, 
    0.006989451, 0.008073906, 0.009917274, 0.01271249, 0.0151462, 0.0194024, 
    0.05106993, 0.04312289, 0, 8.673617e-19, -8.673617e-19, -1.734723e-18, 0, 
    1.734723e-18, 8.673617e-19, 0, 8.673617e-19, 0, -8.673617e-19, 0, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  0.002745586, 0.003016689, 0.003134007, 0.003286961, 0.003427266, 
    0.003466299, 0.003336771, 0.003223558, 0.002931751, 0.003001866, 
    0.003071139, 0.003265308, 0.003608417, 0.003951569, 0.004463761, 
    0.004901127, 0.005332278, 0.00607341, 0.00689303, 0.007821172, 
    0.008642909, 0.009633209, 0.01119329, 0.01351942, 0.0220193, 0.02867593, 
    0.05007729, 0.04564645, 0, 8.673617e-19, -8.673617e-19, -1.734723e-18, 0, 
    1.734723e-18, 8.673617e-19, 0, 8.673617e-19, 0, -8.673617e-19, 0, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  0.003305258, 0.003630027, 0.003739598, 0.003854279, 0.003940701, 0.0039331, 
    0.003718381, 0.003501875, 0.0030472, 0.003060102, 0.003069086, 
    0.003244275, 0.003590056, 0.003935841, 0.0044942, 0.005003709, 
    0.005508439, 0.0064811, 0.007769249, 0.009143161, 0.01011105, 0.01091047, 
    0.01219064, 0.02037869, 0.02445277, 0.04830395, 0.05065713, 0.04821419, 
    0, 8.673617e-19, -8.673617e-19, -1.734723e-18, 0, 1.734723e-18, 
    8.673617e-19, 0, 8.673617e-19, 0, -8.673617e-19, 0, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18,
  0.003855904, 0.004216201, 0.004284468, 0.004330819, 0.004374748, 
    0.004311309, 0.003983061, 0.003635335, 0.002957101, 0.00286885, 
    0.00276154, 0.002820047, 0.003054279, 0.003268183, 0.003740309, 
    0.004224406, 0.004753586, 0.005999716, 0.007921569, 0.009874075, 
    0.01115616, 0.01180296, 0.0150487, 0.02823835, 0.03470651, 0.0471534, 
    0.05368268, 0.05386879, 0, 8.673617e-19, -8.673617e-19, -1.734723e-18, 0, 
    1.734723e-18, 8.673617e-19, 0, 8.673617e-19, 0, -8.673617e-19, 0, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  0.00452162, 0.004897428, 0.004925404, 0.00490219, 0.004836023, 0.004658295, 
    0.004167055, 0.00366533, 0.002708221, 0.002482433, 0.002228964, 
    0.002125552, 0.002175865, 0.002180266, 0.002462834, 0.002820088, 
    0.003269758, 0.004743299, 0.007380534, 0.009982254, 0.01157418, 
    0.01348293, 0.02741744, 0.03121191, 0.04315787, 0.04833487, 0.057462, 
    0.05855403, 0, 8.673617e-19, -8.673617e-19, -1.734723e-18, 0, 
    1.734723e-18, 8.673617e-19, 0, 8.673617e-19, 0, -8.673617e-19, 0, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  0.005348008, 0.005724621, 0.005709933, 0.005628425, 0.005496819, 
    0.005220433, 0.004511091, 0.003785311, 0.002460073, 0.002053944, 
    0.001632109, 0.00131896, 0.001097249, 0.0008061976, 0.0007666165, 
    0.0008707944, 0.001098928, 0.002723739, 0.006140195, 0.009464887, 
    0.01301984, 0.02097558, 0.0297257, 0.03857556, 0.0424727, 0.0510475, 
    0.06386958, 0.06398309, 0, 8.673617e-19, -8.673617e-19, -1.734723e-18, 0, 
    1.734723e-18, 8.673617e-19, 0, 8.673617e-19, 0, -8.673617e-19, 0, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  0.006280207, 0.006655343, 0.00658495, 0.006433909, 0.006261137, 
    0.005957565, 0.005066158, 0.004169795, 0.002476358, 0.0018881, 
    0.001282447, 0.0006898342, 5.691504e-05, -0.0006694979, -0.001245602, 
    -0.001580585, -0.001771024, -9.859996e-05, 0.004165699, 0.008289541, 
    0.01388392, 0.02173754, 0.03263018, 0.03827453, 0.04651425, 0.05679614, 
    0.06898049, 0.06997381, 0, 8.673617e-19, -8.673617e-19, -1.734723e-18, 0, 
    1.734723e-18, 8.673617e-19, 0, 8.673617e-19, 0, -8.673617e-19, 0, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  0.007066691, 0.007472908, 0.007403419, 0.007240133, 0.007093791, 
    0.006863752, 0.005855608, 0.004859428, 0.002882016, 0.002173299, 
    0.001457601, 0.0004455574, -0.0008992646, -0.002365117, -0.00371921, 
    -0.004584947, -0.005275685, -0.003676344, 0.001546915, 0.0066474, 
    0.01355442, 0.02324532, 0.03274816, 0.04199411, 0.05086095, 0.06319769, 
    0.07652815, 0.07477986, 0, 8.673617e-19, -8.673617e-19, -1.734723e-18, 0, 
    1.734723e-18, 8.673617e-19, 0, 8.673617e-19, 0, -8.673617e-19, 0, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  0.00713217, 0.007596852, 0.007400143, 0.006944837, 0.006541848, 
    0.006294188, 0.00529277, 0.004281072, 0.002291195, 0.001473849, 
    0.0004517113, -0.001387262, -0.003706442, -0.006031462, -0.007972136, 
    -0.008880235, -0.009510872, -0.007717863, -0.001429395, 0.004629245, 
    0.01230055, 0.02193025, 0.03611703, 0.04651922, 0.05749697, 0.07042881, 
    0.0828719, 0.07865075, 0, 8.673617e-19, -8.673617e-19, -1.734723e-18, 0, 
    1.734723e-18, 8.673617e-19, 0, 8.673617e-19, 0, -8.673617e-19, 0, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  0.003271171, 0.003776504, 0.003059014, 0.001690226, 0.0004414479, 
    -0.0001938088, -0.00133166, -0.002649051, -0.004924986, -0.006074819, 
    -0.00730653, -0.008864309, -0.01054189, -0.0120192, -0.01348756, 
    -0.01382427, -0.01414538, -0.01201322, -0.005000557, 0.0021192, 0.011948, 
    0.02545537, 0.04116382, 0.05302013, 0.0638717, 0.07836709, 0.08794902, 
    0.08094758, 0, 8.673617e-19, -8.673617e-19, -1.734723e-18, 0, 
    1.734723e-18, 8.673617e-19, 0, 8.673617e-19, 0, -8.673617e-19, 0, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.004140875, -0.003476637, -0.003671465, -0.004221047, -0.004703294, 
    -0.0049373, -0.005800429, -0.006728951, -0.008534708, -0.008986856, 
    -0.009420457, -0.01014758, -0.01116277, -0.01214266, -0.01343594, 
    -0.01416748, -0.01488807, -0.01287708, -0.004270758, 0.004408672, 
    0.01541602, 0.03039634, 0.04769529, 0.05923968, 0.07183851, 0.08472323, 
    0.09125938, 0.08094758, 0, 8.673617e-19, -8.673617e-19, -1.734723e-18, 0, 
    1.734723e-18, 8.673617e-19, 0, 8.673617e-19, 0, -8.673617e-19, 0, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.00813977, -0.007226471, -0.00688359, -0.006695424, -0.006412324, 
    -0.006137896, -0.006691633, -0.007203954, -0.008595685, -0.008320129, 
    -0.007995898, -0.008118376, -0.008728512, -0.00931079, -0.01029462, 
    -0.01111392, -0.01202718, -0.01006404, -0.0009259653, 0.008358764, 
    0.02039756, 0.03594945, 0.05477694, 0.06680391, 0.07826923, 0.08851428, 
    0.09125938, 0.08094758, 0, 8.673617e-19, -8.673617e-19, -1.734723e-18, 0, 
    1.734723e-18, 8.673617e-19, 0, 8.673617e-19, 0, -8.673617e-19, 0, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.008785993, -0.007611498, -0.006588971, -0.005648823, -0.004627598, 
    -0.003789008, -0.004030398, -0.00419053, -0.005351146, -0.00439524, 
    -0.003383914, -0.003049196, -0.003442249, -0.003806908, -0.004550591, 
    -0.00552438, -0.006624551, -0.004661437, 0.004629531, 0.01409162, 
    0.02700994, 0.04408745, 0.06243865, 0.07277806, 0.08066304, 0.08851428, 
    0.09125938, 0.08094758, 0, 8.673617e-19, -8.673617e-19, -1.734723e-18, 0, 
    1.734723e-18, 8.673617e-19, 0, 8.673617e-19, 0, -8.673617e-19, 0, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.006753175, -0.005188119, -0.003478352, -0.002154018, -0.0008297403, 
    0.0003573296, 0.000278877, 0.0001999956, -0.001014721, 0.0003921182, 
    0.001798771, 0.002283757, 0.001847242, 0.001410582, 0.0006414159, 
    -0.0005613465, -0.001763411, 0.0002877256, 0.009644025, 0.0189994, 
    0.03190435, 0.04835555, 0.06479701, 0.07277806, 0.08066304, 0.08851428, 
    0.09125938, 0.08094758, 0, 8.673617e-19, -8.673617e-19, -1.734723e-18, 0, 
    1.734723e-18, 8.673617e-19, 0, 8.673617e-19, 0, -8.673617e-19, 0, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18, 
    -4.336809e-18, -4.336809e-18, -4.336809e-18, -4.336809e-18,
  -0.0006795931, -0.0005994909, -0.0006119221, -0.0007300467, -0.0007090982, 
    -0.0005706056, -0.0004618278, -0.0004744254, -0.0006224862, 
    -0.0008268785, -0.001048036, -0.001094171, -0.0008988921, -0.000636252, 
    -0.0004426108, -0.0002738711, -0.0001258799, -0.0001057276, 
    -0.0001147879, -7.718067e-05, -0.0002608603, -0.0007472949, -0.000977118, 
    -0.002369741, -0.0004425011, 0.002635272, 0.004948918, 0.00673482, 
    1.734723e-18, 0, -8.673617e-19, -2.602085e-18, 8.673617e-19, 
    1.734723e-18, -8.673617e-19, 8.673617e-19, 1.734723e-18, -1.734723e-18, 
    0, 0, -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.0008725795, -0.0008535671, -0.0008557298, -0.0008137668, -0.0006878552, 
    -0.0006492329, -0.0007556408, -0.0009724879, -0.001197319, -0.001373479, 
    -0.001564905, -0.001393335, -0.0009869785, -0.0005897566, -0.0003644988, 
    -0.0002244167, -8.867636e-05, -9.484195e-05, -0.0001721956, 
    -0.0003129923, -0.0006123078, -0.0008591063, -0.001555251, -0.002072017, 
    0.0001164267, 0.0032651, 0.005521978, 0.006945455, 1.734723e-18, 0, 
    -8.673617e-19, -2.602085e-18, 8.673617e-19, 1.734723e-18, -8.673617e-19, 
    8.673617e-19, 1.734723e-18, -1.734723e-18, 0, 0, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.0009881941, -0.001001532, -0.0009162325, -0.0007908851, -0.0006639457, 
    -0.0007137586, -0.0009519622, -0.001173829, -0.001287866, -0.001355686, 
    -0.001408983, -0.001237046, -0.0008626941, -0.0004967123, -0.0002954056, 
    -0.0001962915, -0.0001010979, -0.0001871205, -0.0003752763, 
    -0.0006215594, -0.00088672, -0.000938909, -0.002049383, -0.001817509, 
    0.0005943545, 0.003948116, 0.006012591, 0.007126018, 1.734723e-18, 0, 
    -8.673617e-19, -2.602085e-18, 8.673617e-19, 1.734723e-18, -8.673617e-19, 
    8.673617e-19, 1.734723e-18, -1.734723e-18, 0, 0, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.000989028, -0.0009903844, -0.000897584, -0.0007735812, -0.0006656828, 
    -0.0007108015, -0.0009213778, -0.00111695, -0.001203702, -0.001244894, 
    -0.001272734, -0.001102736, -0.0007558874, -0.0004126982, -0.000222504, 
    -0.0001621202, -0.0001093029, -0.000258003, -0.0005292216, -0.0008153042, 
    -0.0009603637, -0.001031815, -0.002474107, -0.001503247, 0.001283916, 
    0.00457962, 0.00643508, 0.007612907, 1.734723e-18, 0, -8.673617e-19, 
    -2.602085e-18, 8.673617e-19, 1.734723e-18, -8.673617e-19, 8.673617e-19, 
    1.734723e-18, -1.734723e-18, 0, 0, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18,
  -0.0009898078, -0.0009808353, -0.0008864395, -0.0007761457, -0.0006741362, 
    -0.0007082381, -0.0008948658, -0.001067644, -0.001128553, -0.00114326, 
    -0.001145374, -0.000971548, -0.0006398862, -0.0003125003, -0.0001359595, 
    -0.0001206282, -0.000112249, -0.0002911725, -0.0005755661, -0.00087377, 
    -0.001024205, -0.001439214, -0.002286631, -0.0009606783, 0.00193412, 
    0.005127764, 0.006778979, 0.00806847, 1.734723e-18, 0, -8.673617e-19, 
    -2.602085e-18, 8.673617e-19, 1.734723e-18, -8.673617e-19, 8.673617e-19, 
    1.734723e-18, -1.734723e-18, 0, 0, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18,
  -0.0009917429, -0.0009755647, -0.0008829333, -0.0007783978, -0.0006815601, 
    -0.0006874703, -0.0008473003, -0.0009938219, -0.001039579, -0.001036748, 
    -0.001022233, -0.0008493627, -0.0005349416, -0.000224501, -5.995102e-05, 
    -8.418739e-05, -0.0001148365, -0.0003203039, -0.0006162684, 
    -0.0009251182, -0.001080276, -0.001797045, -0.0020212, -0.0004839593, 
    0.002505607, 0.005609824, 0.006963205, 0.008470154, 1.734723e-18, 0, 
    -8.673617e-19, -2.602085e-18, 8.673617e-19, 1.734723e-18, -8.673617e-19, 
    8.673617e-19, 1.734723e-18, -1.734723e-18, 0, 0, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.0009934527, -0.0009708487, -0.0008797959, -0.0007639743, -0.000625778, 
    -0.0006296329, -0.0007817214, -0.000921441, -0.0009599621, -0.0009414364, 
    -0.0009120403, -0.0007400252, -0.0004410314, -0.0001457541, 1.799016e-05, 
    -2.280242e-05, -0.0001062218, -0.0003463725, -0.0006526914, 
    -0.0009839351, -0.001381232, -0.00211728, -0.001783628, -5.718577e-05, 
    0.00301739, 0.006067644, 0.007128431, 0.008830973, 1.734723e-18, 0, 
    -8.673617e-19, -2.602085e-18, 8.673617e-19, 1.734723e-18, -8.673617e-19, 
    8.673617e-19, 1.734723e-18, -1.734723e-18, 0, 0, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.0009940324, -0.0009645417, -0.0008415912, -0.0006973271, -0.000572623, 
    -0.0005765539, -0.0007215377, -0.0008550144, -0.0008868944, 
    -0.0008539653, -0.000809375, -0.0005985496, -0.0002727523, 5.988585e-05, 
    0.0002556954, 0.000180214, 6.502972e-05, -0.0002172226, -0.0006747632, 
    -0.001168573, -0.00166318, -0.002301997, -0.001565557, 0.0003346273, 
    0.003538661, 0.006523228, 0.007280358, 0.009123926, 1.734723e-18, 0, 
    -8.673617e-19, -2.602085e-18, 8.673617e-19, 1.734723e-18, -8.673617e-19, 
    8.673617e-19, 1.734723e-18, -1.734723e-18, 0, 0, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.0009172597, -0.0008785164, -0.0007643729, -0.0006342226, -0.0005222932, 
    -0.0005262957, -0.0006620692, -0.0007395721, -0.0007288881, 
    -0.0006574189, -0.0005678441, -0.0003542102, -3.531677e-05, 0.0002899388, 
    0.0004807739, 0.0003724467, 0.0002271845, -7.800889e-05, -0.0006937878, 
    -0.001343404, -0.001930154, -0.001982918, -0.001191322, 0.0009422498, 
    0.004148792, 0.006954936, 0.007424402, 0.009386417, 1.734723e-18, 0, 
    -8.673617e-19, -2.602085e-18, 8.673617e-19, 1.734723e-18, -8.673617e-19, 
    8.673617e-19, 1.734723e-18, -1.734723e-18, 0, 0, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.0008385051, -0.0007942191, -0.0006887055, -0.0005723853, -0.0003930936, 
    -0.0003461791, -0.0004510048, -0.0005279865, -0.0005208006, 
    -0.0004343741, -0.0003311614, -0.0001147751, 0.0001973533, 0.0005153748, 
    0.0007013356, 0.0005608217, 0.0003860853, 5.841099e-05, -0.0007124305, 
    -0.001514726, -0.002191772, -0.001670237, -0.0006603466, 0.00161548, 
    0.004746777, 0.007378102, 0.007564308, 0.009643859, 1.734723e-18, 0, 
    -8.673617e-19, -2.602085e-18, 8.673617e-19, 1.734723e-18, -8.673617e-19, 
    8.673617e-19, 1.734723e-18, -1.734723e-18, 0, 0, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.0007588133, -0.0007089187, -0.000584371, -0.0003679066, -0.0001775794, 
    -0.0001353548, -0.0002374301, -0.0003138846, -0.0003102385, 
    -0.0002086769, -9.166429e-05, 0.000127507, 0.0004327898, 0.0007434909, 
    0.000975215, 0.0008342922, 0.00061256, 0.000219939, -0.0007164071, 
    -0.001542511, -0.001764835, -0.001353842, -0.0001230725, 0.002296678, 
    0.005351813, 0.007806226, 0.007704456, 0.009904233, 1.734723e-18, 0, 
    -8.673617e-19, -2.602085e-18, 8.673617e-19, 1.734723e-18, -8.673617e-19, 
    8.673617e-19, 1.734723e-18, -1.734723e-18, 0, 0, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.0005266694, -0.0004591836, -0.0003107962, -0.0001206346, 4.570077e-05, 
    8.306602e-05, -1.616015e-05, -9.206897e-05, -7.491966e-05, 6.546668e-05, 
    0.0002287054, 0.0004953298, 0.0008495468, 0.001224841, 0.001479015, 
    0.001337858, 0.001123108, 0.0007449845, -0.0001955347, -0.00103565, 
    -0.001321377, -0.0009289201, 0.0004335087, 0.003002297, 0.005978971, 
    0.00807068, 0.007849528, 0.0123026, 1.734723e-18, 0, -8.673617e-19, 
    -2.602085e-18, 8.673617e-19, 1.734723e-18, -8.673617e-19, 8.673617e-19, 
    1.734723e-18, -1.734723e-18, 0, 0, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18,
  -0.0002341278, -0.0001558838, -2.452178e-05, 0.0001381145, 0.0003521425, 
    0.0004360205, 0.0003639863, 0.0003291263, 0.0003489779, 0.0005085916, 
    0.0006887162, 0.0009720182, 0.001344325, 0.001735551, 0.002006183, 
    0.001864781, 0.001657336, 0.001294384, 0.0003494983, -0.0005052797, 
    -0.0008573552, -5.922332e-05, 0.001281676, 0.003921188, 0.006710694, 
    0.0083295, 0.00801558, 0.01566144, 1.734723e-18, 0, -8.673617e-19, 
    -2.602085e-18, 8.673617e-19, 1.734723e-18, -8.673617e-19, 8.673617e-19, 
    1.734723e-18, -1.734723e-18, 0, 0, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18,
  0.000106642, 0.0002057308, 0.0003834041, 0.0006269142, 0.0008449315, 
    0.0009168527, 0.0008373535, 0.000790604, 0.0007899625, 0.0009695781, 
    0.001167268, 0.001467919, 0.001859044, 0.00228653, 0.002629334, 
    0.002529538, 0.002323876, 0.001941124, 0.0009847849, 0.0002143341, 
    0.0001407794, 0.0008454921, 0.002367973, 0.004979029, 0.007471681, 
    0.008598613, 0.008558657, 0.01915043, 1.734723e-18, 0, -8.673617e-19, 
    -2.602085e-18, 8.673617e-19, 1.734723e-18, -8.673617e-19, 8.673617e-19, 
    1.734723e-18, -1.734723e-18, 0, 0, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18,
  0.0006848875, 0.0008096584, 0.0009657082, 0.001167415, 0.001347092, 
    0.00142482, 0.001352658, 0.001317451, 0.001310771, 0.001532115, 
    0.001776283, 0.002146397, 0.002634068, 0.00315405, 0.003561276, 
    0.003543477, 0.003434308, 0.003158607, 0.002273226, 0.001548324, 
    0.001356419, 0.002053513, 0.003474879, 0.006057394, 0.008186967, 
    0.008088293, 0.009111831, 0.01991375, 1.734723e-18, 0, -8.673617e-19, 
    -2.602085e-18, 8.673617e-19, 1.734723e-18, -8.673617e-19, 8.673617e-19, 
    1.734723e-18, -1.734723e-18, 0, 0, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18,
  0.001273007, 0.00142853, 0.001596538, 0.001815053, 0.002013815, 
    0.002089432, 0.00200032, 0.001942361, 0.001900888, 0.002159142, 
    0.002436648, 0.002859693, 0.003421216, 0.004010005, 0.004494056, 
    0.004573411, 0.004554075, 0.00436227, 0.00354449, 0.002921986, 
    0.002887668, 0.003602234, 0.004909915, 0.00721491, 0.008744719, 
    0.007472627, 0.01553952, 0.02047411, 1.734723e-18, 0, -8.673617e-19, 
    -2.602085e-18, 8.673617e-19, 1.734723e-18, -8.673617e-19, 8.673617e-19, 
    1.734723e-18, -1.734723e-18, 0, 0, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18,
  0.001975492, 0.002171783, 0.002323166, 0.002498104, 0.002658642, 
    0.002721397, 0.002610799, 0.002521671, 0.002428389, 0.002730143, 
    0.003049657, 0.003551399, 0.004234547, 0.004951185, 0.005560554, 
    0.005788101, 0.005934299, 0.005948682, 0.005325865, 0.004875388, 
    0.004744651, 0.005237909, 0.00628533, 0.008297805, 0.009399079, 
    0.008313105, 0.0221335, 0.02056597, 1.734723e-18, 0, -8.673617e-19, 
    -2.602085e-18, 8.673617e-19, 1.734723e-18, -8.673617e-19, 8.673617e-19, 
    1.734723e-18, -1.734723e-18, 0, 0, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18,
  0.002632917, 0.002867966, 0.003006825, 0.003142815, 0.003260811, 
    0.003301183, 0.003157586, 0.003031256, 0.002880652, 0.003233681, 
    0.003594217, 0.004149142, 0.004927218, 0.005733117, 0.006444512, 
    0.006810486, 0.007124359, 0.007366466, 0.006975812, 0.006740442, 
    0.006658338, 0.006923267, 0.00756779, 0.009185295, 0.01021495, 
    0.01267265, 0.02284319, 0.02030747, 1.734723e-18, 0, -8.673617e-19, 
    -2.602085e-18, 8.673617e-19, 1.734723e-18, -8.673617e-19, 8.673617e-19, 
    1.734723e-18, -1.734723e-18, 0, 0, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18,
  0.00323013, 0.003499447, 0.003626313, 0.003719443, 0.00377537, 0.003755703, 
    0.003528252, 0.003298317, 0.002988362, 0.003357033, 0.003730508, 
    0.004368529, 0.005279363, 0.006212207, 0.007068581, 0.007581098, 
    0.008052486, 0.008550343, 0.008471024, 0.008514539, 0.008423148, 
    0.00837146, 0.00862838, 0.01128053, 0.01172792, 0.02141583, 0.02324502, 
    0.01989157, 1.734723e-18, 0, -8.673617e-19, -2.602085e-18, 8.673617e-19, 
    1.734723e-18, -8.673617e-19, 8.673617e-19, 1.734723e-18, -1.734723e-18, 
    0, 0, -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  0.003869441, 0.004144092, 0.004219383, 0.004224211, 0.004224204, 
    0.004129413, 0.003782792, 0.003413907, 0.00287407, 0.003217985, 
    0.003552343, 0.004194607, 0.005161728, 0.006136806, 0.007060443, 
    0.007658185, 0.008256233, 0.00905344, 0.009392872, 0.009808123, 
    0.00982664, 0.009509254, 0.01003649, 0.01389716, 0.01681647, 0.02226011, 
    0.02319981, 0.01762827, 1.734723e-18, 0, -8.673617e-19, -2.602085e-18, 
    8.673617e-19, 1.734723e-18, -8.673617e-19, 8.673617e-19, 1.734723e-18, 
    -1.734723e-18, 0, 0, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  0.004653766, 0.004907534, 0.004936021, 0.00485524, 0.004722351, 0.00448267, 
    0.003956811, 0.003412236, 0.002569122, 0.002853427, 0.00311902, 
    0.003738182, 0.004730125, 0.005716475, 0.006642159, 0.007270582, 
    0.007932782, 0.009008541, 0.009806851, 0.01063509, 0.01077925, 
    0.01066855, 0.01385253, 0.01638389, 0.02148798, 0.02255626, 0.02233925, 
    0.01575297, 1.734723e-18, 0, -8.673617e-19, -2.602085e-18, 8.673617e-19, 
    1.734723e-18, -8.673617e-19, 8.673617e-19, 1.734723e-18, -1.734723e-18, 
    0, 0, -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  0.005621506, 0.005829921, 0.005803811, 0.005638928, 0.005413222, 
    0.005030668, 0.004250145, 0.003447477, 0.002194237, 0.002382537, 
    0.002552596, 0.003127958, 0.004125484, 0.005116706, 0.005975761, 
    0.006592273, 0.007250612, 0.008572031, 0.009853749, 0.01115472, 
    0.01194324, 0.01332229, 0.01629301, 0.02047351, 0.02272214, 0.02246451, 
    0.01949064, 0.0145613, 1.734723e-18, 0, -8.673617e-19, -2.602085e-18, 
    8.673617e-19, 1.734723e-18, -8.673617e-19, 8.673617e-19, 1.734723e-18, 
    -1.734723e-18, 0, 0, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  0.006719056, 0.006865148, 0.006765387, 0.006493522, 0.006180756, 
    0.005694803, 0.00465297, 0.003591233, 0.001870401, 0.001962368, 
    0.002041375, 0.002587839, 0.003610883, 0.00463656, 0.005343311, 
    0.00591396, 0.006507329, 0.008050224, 0.009841967, 0.01167479, 
    0.01329166, 0.01521402, 0.01880028, 0.02235251, 0.02221718, 0.02047048, 
    0.01721848, 0.01394003, 1.734723e-18, 0, -8.673617e-19, -2.602085e-18, 
    8.673617e-19, 1.734723e-18, -8.673617e-19, 8.673617e-19, 1.734723e-18, 
    -1.734723e-18, 0, 0, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  0.00772072, 0.007810989, 0.007667462, 0.007316791, 0.0069595, 0.006434074, 
    0.005156377, 0.003867241, 0.001773235, 0.001836702, 0.001896258, 
    0.002524196, 0.003665208, 0.004804751, 0.005343047, 0.005861107, 
    0.006330964, 0.007987898, 0.01024039, 0.01257515, 0.0147683, 0.0173212, 
    0.02093039, 0.02210056, 0.02117464, 0.01789636, 0.01633918, 0.01344162, 
    1.734723e-18, 0, -8.673617e-19, -2.602085e-18, 8.673617e-19, 
    1.734723e-18, -8.673617e-19, 8.673617e-19, 1.734723e-18, -1.734723e-18, 
    0, 0, -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  0.008484509, 0.008583034, 0.008519467, 0.008267226, 0.008038712, 
    0.007581993, 0.006283501, 0.005020938, 0.003014305, 0.003222889, 
    0.003317008, 0.003656419, 0.004456717, 0.00527835, 0.005430668, 
    0.00592987, 0.006528511, 0.008415408, 0.01107027, 0.01375794, 0.01634729, 
    0.01913633, 0.02076513, 0.02116261, 0.0185829, 0.01656985, 0.01573385, 
    0.01304019, 1.734723e-18, 0, -8.673617e-19, -2.602085e-18, 8.673617e-19, 
    1.734723e-18, -8.673617e-19, 8.673617e-19, 1.734723e-18, -1.734723e-18, 
    0, 0, -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  0.007622677, 0.007693034, 0.007061035, 0.005835292, 0.004625385, 
    0.003781008, 0.002379141, 0.0008718729, -0.001128204, -0.0008937059, 
    -0.0006859132, 1.627397e-05, 0.001233947, 0.002411532, 0.002749208, 
    0.003619482, 0.004643115, 0.007065495, 0.01060672, 0.01394163, 
    0.01626835, 0.0177165, 0.01943339, 0.01872153, 0.01671449, 0.0162292, 
    0.01524939, 0.01279999, 1.734723e-18, 0, -8.673617e-19, -2.602085e-18, 
    8.673617e-19, 1.734723e-18, -8.673617e-19, 8.673617e-19, 1.734723e-18, 
    -1.734723e-18, 0, 0, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  0.00294249, 0.002932566, 0.002357947, 0.001414064, 0.0005767203, 
    -8.297568e-05, -0.001504382, -0.003018738, -0.005098674, -0.004981962, 
    -0.00491103, -0.004140923, -0.002610973, -0.001078442, -0.000704018, 
    0.000190189, 0.001189688, 0.003547718, 0.007124958, 0.01056014, 
    0.01344834, 0.01553809, 0.01715428, 0.01665793, 0.0156523, 0.01595644, 
    0.01493291, 0.01279999, 1.734723e-18, 0, -8.673617e-19, -2.602085e-18, 
    8.673617e-19, 1.734723e-18, -8.673617e-19, 8.673617e-19, 1.734723e-18, 
    -1.734723e-18, 0, 0, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.001282124, -0.001241735, -0.0012323, -0.001646867, -0.002036576, 
    -0.002584551, -0.004130213, -0.005726068, -0.007918946, -0.007856165, 
    -0.007813448, -0.006917656, -0.005143076, -0.003369354, -0.002891575, 
    -0.001898011, -0.0008564772, 0.001482475, 0.004774685, 0.007984505, 
    0.01086143, 0.01324543, 0.01488077, 0.01468325, 0.0147949, 0.01579331, 
    0.01493291, 0.01279999, 1.734723e-18, 0, -8.673617e-19, -2.602085e-18, 
    8.673617e-19, 1.734723e-18, -8.673617e-19, 8.673617e-19, 1.734723e-18, 
    -1.734723e-18, 0, 0, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.003254484, -0.003218693, -0.002871384, -0.003063655, -0.003276432, 
    -0.003808061, -0.005543737, -0.007302122, -0.009722355, -0.009688216, 
    -0.009662742, -0.008752269, -0.006953197, -0.005166065, -0.00454647, 
    -0.003443348, -0.002314714, 3.239703e-05, 0.002826679, 0.005562606, 
    0.008178698, 0.01052443, 0.01257289, 0.01312791, 0.01447562, 0.01579331, 
    0.01493291, 0.01279999, 1.734723e-18, 0, -8.673617e-19, -2.602085e-18, 
    8.673617e-19, 1.734723e-18, -8.673617e-19, 8.673617e-19, 1.734723e-18, 
    -1.734723e-18, 0, 0, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18,
  -0.003301376, -0.003260554, -0.002768698, -0.003094466, -0.003420285, 
    -0.003993794, -0.005979522, -0.00796563, -0.01070964, -0.01070035, 
    -0.01069122, -0.009827685, -0.008109592, -0.006391629, -0.005612175, 
    -0.004417185, -0.003221574, -0.0008817723, 0.001461862, 0.003804673, 
    0.006357829, 0.009118357, 0.01187023, 0.01312791, 0.01447562, 0.01579331, 
    0.01493291, 0.01279999, 1.734723e-18, 0, -8.673617e-19, -2.602085e-18, 
    8.673617e-19, 1.734723e-18, -8.673617e-19, 8.673617e-19, 1.734723e-18, 
    -1.734723e-18, 0, 0, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, 
    -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18, -6.071532e-18 ;

 temp_west =
  1.137725, 1.138502, 1.136654, 1.134171, 1.132539, 1.132293, 1.133186, 
    1.134001, 1.132972, 1.129846, 1.125488, 1.120774, 1.117511, 1.115659, 
    1.114885, 1.114359, 1.114028, 1.113606, 1.11334, 1.11447, 1.116616, 
    1.118535, 1.120631, 1.121848, 1.122246, 1.124431, 1.128423, 1.13209, 
    1.139097, 1.155439, 1.173234, 1.191265, 1.203188, 1.215801, 1.225897, 
    1.230901, 1.231603, 1.229766, 1.22669, 1.224867, 1.226371, 1.227922, 
    1.226231, 1.223652, 1.222011, 1.220882, 1.221794, 1.225152, 1.22797, 
    1.228305, 1.228361, 1.231949, 1.239335, 1.246062, 1.245957,
  1.165706, 1.165869, 1.162951, 1.160826, 1.159603, 1.159553, 1.160453, 
    1.161237, 1.160347, 1.156453, 1.149617, 1.141817, 1.135718, 1.132736, 
    1.131714, 1.131402, 1.131398, 1.131247, 1.131173, 1.132387, 1.135486, 
    1.139327, 1.142602, 1.14519, 1.147001, 1.150447, 1.156169, 1.161097, 
    1.168691, 1.192465, 1.220587, 1.236734, 1.252448, 1.271241, 1.285827, 
    1.292801, 1.293334, 1.28976, 1.284302, 1.28098, 1.28309, 1.285208, 
    1.282291, 1.278021, 1.275158, 1.273021, 1.274281, 1.2795, 1.283914, 
    1.28435, 1.284357, 1.289735, 1.300864, 1.310501, 1.310103,
  1.209825, 1.209718, 1.205902, 1.201692, 1.199112, 1.198701, 1.200008, 
    1.201094, 1.199339, 1.192526, 1.180784, 1.167589, 1.161353, 1.158691, 
    1.157714, 1.157151, 1.157052, 1.156755, 1.15662, 1.158592, 1.162381, 
    1.166008, 1.169129, 1.172724, 1.175626, 1.181208, 1.190407, 1.198399, 
    1.210477, 1.234884, 1.276182, 1.300798, 1.316836, 1.333686, 1.346634, 
    1.353082, 1.353789, 1.349381, 1.344143, 1.340921, 1.342727, 1.34453, 
    1.341717, 1.337696, 1.334966, 1.332903, 1.33394, 1.338567, 1.342425, 
    1.342663, 1.342453, 1.347103, 1.36265, 1.378188, 1.377501,
  1.26423, 1.263827, 1.256817, 1.249049, 1.244045, 1.242975, 1.245036, 
    1.246723, 1.243428, 1.231266, 1.219582, 1.207299, 1.197806, 1.193167, 
    1.19136, 1.190238, 1.189782, 1.189076, 1.188707, 1.191774, 1.197881, 
    1.203783, 1.208825, 1.212865, 1.215783, 1.221125, 1.229811, 1.237682, 
    1.256805, 1.295278, 1.335309, 1.362036, 1.388048, 1.415319, 1.436419, 
    1.446209, 1.446395, 1.440163, 1.431095, 1.425319, 1.427641, 1.430112, 
    1.425069, 1.418078, 1.413326, 1.409777, 1.411161, 1.4184, 1.424359, 
    1.424519, 1.424067, 1.431624, 1.447731, 1.461604, 1.460587,
  1.327183, 1.326464, 1.31968, 1.312243, 1.307458, 1.306272, 1.307942, 
    1.309229, 1.305875, 1.294285, 1.274712, 1.252877, 1.23609, 1.228443, 
    1.226767, 1.22578, 1.225507, 1.224976, 1.224733, 1.2277, 1.233692, 
    1.2436, 1.251911, 1.25841, 1.262919, 1.271271, 1.285086, 1.296971, 
    1.31453, 1.349878, 1.413756, 1.450677, 1.474346, 1.499224, 1.51831, 
    1.526931, 1.526666, 1.520461, 1.511686, 1.506011, 1.50794, 1.509921, 
    1.504868, 1.498052, 1.493243, 1.489482, 1.490282, 1.496533, 1.501637, 
    1.501339, 1.500476, 1.507023, 1.521479, 1.535462, 1.534149,
  1.405654, 1.404546, 1.392665, 1.379531, 1.370858, 1.368611, 1.371466, 
    1.373695, 1.36787, 1.349624, 1.331143, 1.310536, 1.294595, 1.286596, 
    1.283243, 1.28102, 1.279815, 1.278272, 1.277334, 1.281842, 1.291185, 
    1.300172, 1.307736, 1.313657, 1.317768, 1.325456, 1.338167, 1.349035, 
    1.375654, 1.433913, 1.49464, 1.528518, 1.55013, 1.587443, 1.618097, 
    1.631998, 1.63172, 1.621846, 1.60776, 1.59854, 1.60116, 1.604042, 
    1.595935, 1.585058, 1.577484, 1.571683, 1.572978, 1.582859, 1.590877, 
    1.590512, 1.589363, 1.599964, 1.622993, 1.642768, 1.640938,
  1.499188, 1.49762, 1.48604, 1.473315, 1.464844, 1.462306, 1.464469, 
    1.465995, 1.459966, 1.440579, 1.408276, 1.372446, 1.346942, 1.339243, 
    1.33592, 1.333698, 1.332524, 1.330993, 1.329984, 1.334078, 1.342625, 
    1.35137, 1.363851, 1.373394, 1.379741, 1.391994, 1.412722, 1.430447, 
    1.456884, 1.510794, 1.575422, 1.630195, 1.664987, 1.701417, 1.729236, 
    1.741476, 1.740534, 1.730575, 1.716726, 1.707442, 1.709338, 1.711383, 
    1.703099, 1.692317, 1.684545, 1.67836, 1.6788, 1.687244, 1.693963, 
    1.692891, 1.691096, 1.700254, 1.721007, 1.738783, 1.736491,
  1.58502, 1.58303, 1.571727, 1.559377, 1.551091, 1.548286, 1.549814, 
    1.550695, 1.544478, 1.525755, 1.49499, 1.460907, 1.434519, 1.420935, 
    1.41482, 1.410476, 1.407588, 1.404257, 1.401981, 1.408287, 1.422311, 
    1.435819, 1.446981, 1.455455, 1.461003, 1.472061, 1.491004, 1.50713, 
    1.531424, 1.599777, 1.690443, 1.740868, 1.772671, 1.80601, 1.831228, 
    1.841943, 1.840392, 1.830354, 1.816723, 1.80738, 1.808612, 1.809889, 
    1.801443, 1.790746, 1.782794, 1.776256, 1.77591, 1.783037, 1.788563, 
    1.786842, 1.784455, 1.792289, 1.810954, 1.828109, 1.825388,
  1.719404, 1.716673, 1.698593, 1.678692, 1.665154, 1.660719, 1.663494, 
    1.665296, 1.655634, 1.625708, 1.577091, 1.544662, 1.519369, 1.506095, 
    1.499818, 1.49523, 1.492063, 1.488463, 1.485827, 1.4912, 1.503739, 
    1.515774, 1.525687, 1.53315, 1.537942, 1.547868, 1.569997, 1.59603, 
    1.635125, 1.715568, 1.799347, 1.845655, 1.874629, 1.918793, 1.956957, 
    1.973582, 1.971984, 1.957718, 1.937938, 1.924411, 1.926282, 1.928464, 
    1.91638, 1.900847, 1.889559, 1.880529, 1.880658, 1.89187, 1.900633, 
    1.898738, 1.895932, 1.908437, 1.937093, 1.961666, 1.958394,
  1.859259, 1.855749, 1.838025, 1.818637, 1.805269, 1.800304, 1.801989, 
    1.802683, 1.792677, 1.763808, 1.716685, 1.664611, 1.624204, 1.602982, 
    1.592939, 1.585473, 1.579946, 1.573877, 1.569512, 1.577932, 1.598076, 
    1.617599, 1.633537, 1.645392, 1.652806, 1.668426, 1.695979, 1.719423, 
    1.755063, 1.829032, 1.915863, 1.985098, 2.028548, 2.073987, 2.10833, 
    2.122746, 2.120312, 2.106001, 2.086602, 2.073029, 2.073863, 2.074894, 
    2.062599, 2.047135, 2.035516, 2.0259, 2.024862, 2.034087, 2.041019, 
    2.038147, 2.034472, 2.045046, 2.070631, 2.092541, 2.088728,
  2.003505, 1.999185, 1.979117, 1.960248, 1.947051, 1.941552, 1.942132, 
    1.941706, 1.931353, 1.903553, 1.858914, 1.80967, 1.771131, 1.750372, 
    1.739949, 1.731938, 1.725748, 1.719084, 1.714016, 1.720718, 1.738248, 
    1.755235, 1.76901, 1.779106, 1.785193, 1.798838, 1.823462, 1.844284, 
    1.876429, 1.974722, 2.088298, 2.151148, 2.190195, 2.231027, 2.261504, 
    2.273685, 2.270406, 2.25605, 2.237034, 2.223415, 2.2232, 2.223067, 
    2.210559, 2.195164, 2.18321, 2.173, 2.170782, 2.177996, 2.183075, 
    2.179215, 2.174662, 2.18328, 2.205759, 2.224973, 2.220614,
  2.230664, 2.224898, 2.200686, 2.17434, 2.155729, 2.148175, 2.149394, 
    2.149296, 2.13534, 2.096834, 2.034321, 1.965167, 1.923359, 1.903078, 
    1.892262, 1.883688, 1.876809, 1.869529, 1.863732, 1.868655, 1.883477, 
    1.897835, 1.909623, 1.924333, 1.933172, 1.952949, 1.988814, 2.019352, 
    2.066318, 2.164618, 2.266952, 2.323184, 2.35767, 2.40836, 2.449283, 
    2.466026, 2.462348, 2.444016, 2.419407, 2.401837, 2.401696, 2.40183, 
    2.385781, 2.365818, 2.350523, 2.337647, 2.335286, 2.345274, 2.3524, 
    2.347902, 2.342565, 2.354606, 2.384929, 2.411027, 2.406135,
  2.468373, 2.461094, 2.437364, 2.411836, 2.393378, 2.384919, 2.384404, 
    2.38258, 2.368296, 2.331948, 2.273983, 2.210025, 2.159558, 2.131534, 
    2.1166, 2.104649, 2.094757, 2.084439, 2.076354, 2.083296, 2.104495, 
    2.125328, 2.142092, 2.154137, 2.161005, 2.177691, 2.208786, 2.235056, 
    2.276223, 2.363334, 2.489286, 2.563045, 2.60835, 2.655581, 2.690393, 
    2.70362, 2.698639, 2.680242, 2.656213, 2.638512, 2.636628, 2.634803, 
    2.618251, 2.598137, 2.582042, 2.567945, 2.563562, 2.57025, 2.574342, 
    2.568267, 2.561585, 2.570658, 2.596298, 2.61842, 2.612982,
  2.775254, 2.765999, 2.736813, 2.705523, 2.68265, 2.67219, 2.671667, 
    2.669617, 2.652398, 2.608073, 2.536834, 2.464765, 2.418084, 2.391267, 
    2.376028, 2.363451, 2.352665, 2.34162, 2.332664, 2.336896, 2.353846, 
    2.370616, 2.383942, 2.393216, 2.398032, 2.417743, 2.457514, 2.49125, 
    2.54407, 2.65563, 2.771487, 2.834893, 2.873055, 2.912774, 2.941228, 
    2.950798, 2.944462, 2.925997, 2.902571, 2.884734, 2.881036, 2.877172, 
    2.860098, 2.839827, 2.8229, 2.807532, 2.801046, 2.8043, 2.805236, 
    2.797522, 2.78944, 2.795425, 2.820537, 2.848446, 2.842401,
  3.123553, 3.112048, 3.083724, 3.053981, 3.03161, 3.020234, 3.017715, 
    3.013731, 2.996715, 2.956358, 2.892657, 2.822315, 2.766174, 2.733838, 
    2.715416, 2.700095, 2.686683, 2.673075, 2.662158, 2.667319, 2.688432, 
    2.709607, 2.726646, 2.738609, 2.744943, 2.762047, 2.794959, 2.822474, 
    2.866724, 2.961263, 3.085148, 3.163843, 3.211107, 3.260133, 3.295207, 
    3.307054, 3.299393, 3.276669, 3.247666, 3.225413, 3.220383, 3.21508, 
    3.193474, 3.167759, 3.14617, 3.126503, 3.117922, 3.121167, 3.12155, 
    3.111715, 3.101613, 3.108693, 3.133798, 3.155715, 3.148876,
  3.559371, 3.545696, 3.511822, 3.476258, 3.44935, 3.43589, 3.433335, 
    3.429035, 3.409059, 3.360882, 3.28425, 3.199647, 3.132374, 3.102112, 
    3.084107, 3.068723, 3.05482, 3.040971, 3.029616, 3.031581, 3.047275, 
    3.067347, 3.088518, 3.103465, 3.111504, 3.13249, 3.172566, 3.206036, 
    3.259716, 3.37398, 3.491772, 3.555281, 3.592036, 3.630072, 3.655783, 
    3.662233, 3.652563, 3.629632, 3.601311, 3.5786, 3.570722, 3.562088, 
    3.539161, 3.512545, 3.489016, 3.466711, 3.454475, 3.452223, 3.447549, 
    3.434917, 3.422435, 3.42484, 3.44752, 3.473412, 3.465548,
  4.023047, 4.007346, 3.975441, 3.942612, 3.917077, 3.902914, 3.898022, 
    3.891366, 3.871838, 3.8291, 3.762476, 3.689149, 3.630002, 3.595009, 
    3.573808, 3.555584, 3.538504, 3.521872, 3.508564, 3.510311, 3.528586, 
    3.547527, 3.563364, 3.574159, 3.579348, 3.594784, 3.625677, 3.650816, 
    3.692876, 3.805308, 3.949027, 4.025674, 4.069403, 4.114581, 4.144781, 
    4.152066, 4.140351, 4.11241, 4.077727, 4.04961, 4.039457, 4.027731, 
    3.998125, 3.963896, 3.93301, 3.903224, 3.886081, 3.880543, 3.871883, 
    3.854603, 3.837617, 3.837986, 3.856843, 3.87338, 3.862947,
  4.731818, 4.71242, 4.669348, 4.624045, 4.588967, 4.569139, 4.56151, 
    4.551352, 4.523611, 4.464725, 4.374134, 4.2756, 4.196838, 4.150838, 
    4.123027, 4.099107, 4.075921, 4.053942, 4.036788, 4.037532, 4.059029, 
    4.081366, 4.100572, 4.113488, 4.119551, 4.13707, 4.173368, 4.20276, 
    4.251678, 4.359194, 4.468636, 4.524206, 4.573597, 4.629857, 4.667295, 
    4.67685, 4.663682, 4.630015, 4.58777, 4.553617, 4.542283, 4.528063, 
    4.49014, 4.446217, 4.40581, 4.366151, 4.343036, 4.333775, 4.319823, 
    4.296099, 4.272552, 4.269271, 4.287901, 4.303104, 4.287123,
  5.654085, 5.625742, 5.557993, 5.486111, 5.430552, 5.399023, 5.386184, 
    5.370083, 5.326245, 5.234464, 5.095635, 4.946298, 4.840849, 4.795218, 
    4.763936, 4.73568, 4.70603, 4.678937, 4.657268, 4.646976, 4.654587, 
    4.66433, 4.687347, 4.70367, 4.710941, 4.73156, 4.776309, 4.812269, 
    4.871254, 5.003207, 5.136427, 5.200052, 5.231337, 5.265146, 5.283628, 
    5.28334, 5.26837, 5.235516, 5.19609, 5.163295, 5.150354, 5.130974, 
    5.088666, 5.041205, 4.992501, 4.94036, 4.904698, 4.878341, 4.846599, 
    4.810831, 4.775123, 4.755386, 4.75584, 4.754798, 4.730273,
  6.825705, 6.781668, 6.675507, 6.57273, 6.508284, 6.462278, 6.430555, 
    6.396846, 6.340583, 6.246028, 6.114827, 5.974074, 5.856639, 5.780448, 
    5.724843, 5.673025, 5.617599, 5.566912, 5.524918, 5.495625, 5.491825, 
    5.492064, 5.495114, 5.493886, 5.488145, 5.489003, 5.510376, 5.526628, 
    5.559396, 5.728868, 5.900308, 5.977363, 6.01307, 6.053519, 6.07349, 
    6.074037, 6.060887, 6.023654, 5.979807, 5.946347, 5.939883, 5.922037, 
    5.870718, 5.812041, 5.746742, 5.672052, 5.62159, 5.580136, 5.527823, 
    5.472351, 5.414687, 5.375057, 5.361985, 5.344921, 5.297616,
  8.676331, 8.595848, 8.471599, 8.346244, 8.237016, 8.157437, 8.100881, 
    8.045774, 7.953738, 7.801104, 7.59687, 7.376722, 7.190806, 7.066184, 
    6.970728, 6.879096, 6.781882, 6.69134, 6.613207, 6.551422, 6.527483, 
    6.510912, 6.499774, 6.485325, 6.467698, 6.456429, 6.474345, 6.487192, 
    6.520079, 6.626163, 6.780048, 6.864777, 6.899669, 6.941815, 6.956142, 
    6.952608, 6.939071, 6.895202, 6.847341, 6.815419, 6.81612, 6.800321, 
    6.74193, 6.674014, 6.592522, 6.494172, 6.427887, 6.368834, 6.293298, 
    6.216701, 6.134738, 6.072187, 6.043503, 6.008234, 5.933947,
  10.92399, 10.7879, 10.60321, 10.42442, 10.26358, 10.14314, 10.05455, 
    9.971041, 9.839475, 9.630086, 9.35834, 9.06506, 8.812864, 8.636262, 
    8.493466, 8.352574, 8.20446, 8.063465, 7.937002, 7.830443, 7.775229, 
    7.732022, 7.69755, 7.661808, 7.625006, 7.593922, 7.601059, 7.602906, 
    7.628404, 7.742479, 7.851549, 7.877754, 7.887586, 7.907933, 7.895561, 
    7.878428, 7.864923, 7.817691, 7.772526, 7.749176, 7.760442, 7.747539, 
    7.682865, 7.608694, 7.511736, 7.388757, 7.303734, 7.221697, 7.118603, 
    7.019697, 6.912338, 6.821233, 6.766976, 6.704464, 6.601238,
  13.22495, 13.02462, 12.7862, 12.5633, 12.35516, 12.19126, 12.06304, 
    11.94365, 11.77647, 11.533, 11.2324, 10.90891, 10.62238, 10.40854, 
    10.22297, 10.03504, 9.838056, 9.647323, 9.469985, 9.309077, 9.204234, 
    9.116638, 9.044448, 8.975874, 8.910616, 8.846611, 8.822427, 8.792747, 
    8.787745, 8.866357, 8.931381, 8.915253, 8.872767, 8.854485, 8.819829, 
    8.797163, 8.795793, 8.753751, 8.717427, 8.712023, 8.750308, 8.747168, 
    8.666633, 8.580659, 8.460798, 8.30255, 8.189425, 8.082174, 7.951546, 
    7.826762, 7.691759, 7.575552, 7.502339, 7.415859, 7.280087,
  15.41727, 15.16509, 14.88535, 14.62688, 14.3758, 14.17178, 14.00721, 
    13.85827, 13.66011, 13.38457, 13.0561, 12.70041, 12.37774, 12.12908, 
    11.90594, 11.67847, 11.43672, 11.20397, 10.98687, 10.78072, 10.6323, 
    10.50602, 10.40455, 10.31126, 10.22533, 10.13736, 10.088, 10.02786, 
    10.0056, 10.06392, 10.08864, 10.03983, 9.969115, 9.923856, 9.867879, 
    9.864956, 9.909823, 9.911548, 9.914508, 9.952141, 10.04151, 10.04889, 
    9.939241, 9.833719, 9.681492, 9.473606, 9.304961, 9.141584, 8.966027, 
    8.79847, 8.621914, 8.465683, 8.354024, 8.229898, 8.053718,
  17.43805, 17.17404, 16.88912, 16.62444, 16.36119, 16.1426, 15.96362, 
    15.80602, 15.59073, 15.2889, 14.93828, 14.55181, 14.18885, 13.90351, 
    13.63924, 13.3659, 13.06507, 12.78186, 12.52409, 12.26156, 12.07919, 
    11.93666, 11.84283, 11.76286, 11.69478, 11.61959, 11.57308, 11.49393, 
    11.47701, 11.5408, 11.5527, 11.49708, 11.4219, 11.38569, 11.29868, 
    11.28216, 11.33744, 11.36676, 11.377, 11.38744, 11.42166, 11.3566, 
    11.18467, 10.99527, 10.77449, 10.51982, 10.29464, 10.0879, 9.896707, 
    9.706484, 9.513761, 9.320834, 9.136243, 8.956052, 8.775131,
  18.46674, 18.20966, 17.9756, 17.7699, 17.55877, 17.37451, 17.21738, 
    17.07159, 16.90451, 16.70299, 16.46736, 16.2, 15.91904, 15.67768, 
    15.42891, 15.16199, 14.87182, 14.59086, 14.3247, 14.04446, 13.84783, 
    13.69808, 13.62572, 13.55577, 13.48407, 13.38997, 13.28324, 13.11452, 
    12.98815, 12.90162, 12.7814, 12.63643, 12.4749, 12.3843, 12.25562, 
    12.18342, 12.16835, 12.13684, 12.06942, 11.9662, 11.86347, 11.69498, 
    11.46032, 11.21737, 10.95553, 10.67453, 10.4106, 10.17247, 9.95995, 
    9.75638, 9.564767, 9.385315, 9.204858, 9.038293, 8.885454,
  18.56439, 18.30234, 18.07619, 17.88571, 17.68764, 17.51923, 17.38043, 
    17.24464, 17.10852, 16.97208, 16.80638, 16.62722, 16.43478, 16.28563, 
    16.1251, 15.95303, 15.75149, 15.56609, 15.39659, 15.20831, 15.03321, 
    14.87021, 14.76188, 14.6301, 14.47402, 14.28348, 14.04729, 13.76406, 
    13.49733, 13.21655, 12.91719, 12.67588, 12.5061, 12.41047, 12.27516, 
    12.19945, 12.18329, 12.14971, 12.08219, 11.98077, 11.87936, 11.71088, 
    11.4753, 11.22666, 10.96312, 10.6847, 10.4199, 10.18171, 9.970098, 
    9.765129, 9.572428, 9.392069, 9.210578, 9.043533, 8.890863,
  18.56682, 18.30254, 18.07548, 17.88565, 17.68724, 17.51835, 17.37898, 
    17.24247, 17.10638, 16.97069, 16.80623, 16.62786, 16.43567, 16.28775, 
    16.13278, 15.97075, 15.77048, 15.59897, 15.45623, 15.27586, 15.10988, 
    14.95826, 14.84643, 14.70333, 14.52896, 14.32355, 14.07619, 13.78688, 
    13.51443, 13.22469, 12.91791, 12.67559, 12.50644, 12.41029, 12.27594, 
    12.20065, 12.18455, 12.15113, 12.08369, 11.98224, 11.88074, 11.71216, 
    11.47647, 11.22828, 10.96492, 10.68638, 10.42157, 10.18371, 9.972793, 
    9.76839, 9.575872, 9.395262, 9.213336, 9.046055, 8.893392,
  18.56869, 18.30292, 18.07522, 17.88556, 17.68716, 17.51835, 17.37912, 
    17.24281, 17.10679, 16.97107, 16.80702, 16.62892, 16.43679, 16.28907, 
    16.13421, 15.9722, 15.77185, 15.60035, 15.45769, 15.27712, 15.11097, 
    14.95922, 14.84743, 14.7038, 14.5283, 14.32252, 14.07509, 13.78605, 
    13.51414, 13.22568, 12.92076, 12.67883, 12.50944, 12.41262, 12.27645, 
    12.20053, 12.18491, 12.15161, 12.08442, 11.9833, 11.88187, 11.71328, 
    11.47752, 11.22914, 10.96571, 10.68723, 10.42243, 10.18459, 9.973706, 
    9.769499, 9.577046, 9.396339, 9.214319, 9.047004, 8.894401,
  18.57084, 18.30304, 18.07437, 17.88482, 17.68601, 17.51711, 17.37812, 
    17.24216, 17.10631, 16.97057, 16.80673, 16.62878, 16.43674, 16.28919, 
    16.13453, 15.97274, 15.77251, 15.60113, 15.4586, 15.27811, 15.11219, 
    14.96083, 14.8494, 14.70617, 14.53114, 14.32548, 14.0782, 13.78929, 
    13.51782, 13.22949, 12.92422, 12.6816, 12.5115, 12.4139, 12.27684, 
    12.20052, 12.18494, 12.15153, 12.08445, 11.98371, 11.88231, 11.71358, 
    11.47752, 11.22887, 10.96525, 10.68665, 10.42182, 10.18405, 9.97333, 
    9.768906, 9.576345, 9.395651, 9.213738, 9.046537, 8.894047,
  1.137597, 1.138368, 1.136519, 1.134045, 1.132428, 1.132173, 1.133031, 
    1.133825, 1.13267, 1.129336, 1.124939, 1.120284, 1.117102, 1.115341, 
    1.114629, 1.114161, 1.11388, 1.113489, 1.113231, 1.114385, 1.116523, 
    1.118395, 1.120454, 1.121654, 1.122057, 1.124231, 1.12822, 1.131908, 
    1.138938, 1.155203, 1.172869, 1.190703, 1.202482, 1.214961, 1.225012, 
    1.229991, 1.230659, 1.228839, 1.225798, 1.224017, 1.225556, 1.227125, 
    1.225449, 1.222935, 1.221345, 1.220256, 1.221151, 1.224493, 1.227316, 
    1.227668, 1.227769, 1.231411, 1.238846, 1.245597, 1.2455,
  1.165555, 1.165723, 1.1628, 1.160666, 1.159443, 1.159371, 1.160226, 
    1.16098, 1.159921, 1.155743, 1.148792, 1.140971, 1.1349, 1.132031, 
    1.13113, 1.130959, 1.131071, 1.13099, 1.130941, 1.132219, 1.13531, 
    1.139072, 1.142298, 1.144866, 1.146687, 1.150106, 1.155804, 1.16074, 
    1.168349, 1.192041, 1.219939, 1.235867, 1.251409, 1.270045, 1.284608, 
    1.291537, 1.292002, 1.28847, 1.283075, 1.279815, 1.281982, 1.284105, 
    1.281176, 1.276991, 1.274182, 1.272072, 1.273261, 1.278428, 1.282854, 
    1.283346, 1.28344, 1.288903, 1.30016, 1.309891, 1.309547,
  1.209679, 1.209597, 1.205782, 1.201553, 1.198959, 1.198508, 1.199744, 
    1.200773, 1.198788, 1.191603, 1.179706, 1.166496, 1.160293, 1.157772, 
    1.156949, 1.156569, 1.156615, 1.156407, 1.156302, 1.158352, 1.162133, 
    1.165665, 1.168716, 1.172268, 1.175159, 1.180686, 1.189857, 1.197883, 
    1.20999, 1.234286, 1.275309, 1.299677, 1.315515, 1.332192, 1.345104, 
    1.35148, 1.352082, 1.347724, 1.342552, 1.339389, 1.341276, 1.343077, 
    1.340209, 1.336262, 1.333565, 1.331499, 1.332423, 1.336998, 1.340906, 
    1.341266, 1.341195, 1.345972, 1.361745, 1.377438, 1.376846,
  1.264199, 1.263831, 1.256801, 1.248982, 1.243938, 1.242802, 1.244763, 
    1.24636, 1.24277, 1.230137, 1.218223, 1.205891, 1.196461, 1.191997, 
    1.190387, 1.189499, 1.189219, 1.188622, 1.188293, 1.191453, 1.197549, 
    1.203333, 1.208282, 1.212263, 1.215158, 1.220424, 1.229091, 1.237035, 
    1.256195, 1.294542, 1.334254, 1.360697, 1.38648, 1.413544, 1.434588, 
    1.444279, 1.444323, 1.438123, 1.429101, 1.42336, 1.425742, 1.428192, 
    1.423092, 1.416184, 1.411474, 1.407932, 1.409201, 1.416408, 1.422455, 
    1.422781, 1.422509, 1.430235, 1.446621, 1.460696, 1.459817,
  1.327358, 1.326673, 1.319858, 1.312347, 1.307485, 1.306191, 1.307716, 
    1.308864, 1.305142, 1.292985, 1.273104, 1.251193, 1.234481, 1.227028, 
    1.225583, 1.224879, 1.224808, 1.224406, 1.224216, 1.227296, 1.233277, 
    1.24306, 1.251267, 1.257695, 1.26217, 1.270429, 1.284228, 1.296201, 
    1.313815, 1.349024, 1.412534, 1.449146, 1.472557, 1.497193, 1.516215, 
    1.524717, 1.524277, 1.518086, 1.509331, 1.503658, 1.505623, 1.50757, 
    1.502454, 1.49572, 1.490963, 1.487231, 1.487931, 1.494176, 1.499403, 
    1.499304, 1.498658, 1.505411, 1.520191, 1.534411, 1.533274,
  1.406091, 1.405018, 1.393074, 1.379819, 1.37102, 1.368624, 1.371294, 
    1.373338, 1.367079, 1.348173, 1.329312, 1.308606, 1.292769, 1.284984, 
    1.281898, 1.280007, 1.279024, 1.277626, 1.276757, 1.281397, 1.290738, 
    1.299588, 1.30703, 1.312864, 1.316925, 1.324499, 1.33719, 1.348157, 
    1.374843, 1.432945, 1.493267, 1.526819, 1.548147, 1.58512, 1.615633, 
    1.629349, 1.628844, 1.618976, 1.604909, 1.595675, 1.598294, 1.601113, 
    1.592958, 1.582194, 1.574706, 1.568971, 1.570179, 1.580051, 1.588208, 
    1.58809, 1.587201, 1.598029, 1.621386, 1.641421, 1.639819,
  1.49994, 1.498409, 1.48675, 1.473869, 1.465218, 1.462478, 1.464405, 
    1.465685, 1.459164, 1.43906, 1.406292, 1.370314, 1.344921, 1.337454, 
    1.334431, 1.332588, 1.331654, 1.330285, 1.329361, 1.333603, 1.34215, 
    1.350746, 1.363089, 1.372529, 1.378811, 1.390927, 1.411629, 1.429464, 
    1.455979, 1.509722, 1.573882, 1.628219, 1.662633, 1.698672, 1.726335, 
    1.738356, 1.737133, 1.727147, 1.713274, 1.703927, 1.705789, 1.70775, 
    1.699404, 1.688726, 1.681051, 1.67496, 1.67535, 1.683836, 1.690751, 
    1.689992, 1.688514, 1.697948, 1.719084, 1.737172, 1.735154,
  1.586061, 1.58411, 1.572714, 1.560174, 1.55166, 1.548604, 1.549848, 
    1.550427, 1.543667, 1.524175, 1.492892, 1.458649, 1.432399, 1.419033, 
    1.413229, 1.40929, 1.40664, 1.40348, 1.401306, 1.407768, 1.421794, 
    1.435152, 1.446164, 1.454521, 1.459985, 1.470887, 1.489802, 1.506051, 
    1.530434, 1.598539, 1.688592, 1.738568, 1.769966, 1.802878, 1.827926, 
    1.838391, 1.836509, 1.826414, 1.81272, 1.803268, 1.804435, 1.80561, 
    1.797088, 1.786489, 1.778642, 1.772225, 1.771864, 1.779078, 1.784853, 
    1.783506, 1.781488, 1.789643, 1.808741, 1.826248, 1.823844,
  1.720763, 1.718073, 1.699879, 1.679747, 1.665924, 1.661185, 1.663624, 
    1.665064, 1.654807, 1.62407, 1.574886, 1.542284, 1.517161, 1.504097, 
    1.498138, 1.493978, 1.491039, 1.487614, 1.485098, 1.490633, 1.503179, 
    1.515067, 1.524819, 1.532151, 1.536841, 1.546594, 1.568674, 1.594799, 
    1.633928, 1.71405, 1.797201, 1.843049, 1.871592, 1.915253, 1.95318, 
    1.969486, 1.96749, 1.953135, 1.933273, 1.919607, 1.921372, 1.923422, 
    1.911272, 1.895859, 1.884705, 1.875834, 1.87598, 1.887301, 1.896347, 
    1.894886, 1.892501, 1.905351, 1.934439, 1.959377, 1.95647,
  1.860936, 1.857469, 1.839615, 1.81996, 1.80625, 1.800924, 1.802215, 
    1.802483, 1.791831, 1.762111, 1.714365, 1.662099, 1.621888, 1.600866, 
    1.591147, 1.584132, 1.578827, 1.572944, 1.568722, 1.577296, 1.597415, 
    1.616766, 1.632511, 1.644203, 1.651483, 1.66689, 1.694366, 1.717906, 
    1.753592, 1.82724, 1.9134, 1.982094, 2.02504, 2.069913, 2.103995, 
    2.118044, 2.11514, 2.100682, 2.081138, 2.067365, 2.068053, 2.068934, 
    2.056569, 2.04122, 2.029752, 2.020331, 2.019362, 2.028757, 2.036033, 
    2.033664, 2.03047, 2.041441, 2.067507, 2.089832, 2.086432,
  2.005498, 2.001224, 1.981014, 1.961842, 1.948246, 1.942327, 1.942457, 
    1.941538, 1.930487, 1.901796, 1.856477, 1.807011, 1.768667, 1.748045, 
    1.737907, 1.730331, 1.724312, 1.717821, 1.71292, 1.719782, 1.737306, 
    1.754149, 1.767733, 1.777655, 1.783586, 1.797008, 1.821554, 1.84248, 
    1.874681, 1.972548, 2.085356, 2.147674, 2.186196, 2.226415, 2.256604, 
    2.268369, 2.264548, 2.249985, 2.230762, 2.216883, 2.21648, 2.216177, 
    2.203594, 2.188311, 2.176524, 2.166547, 2.164451, 2.171896, 2.177382, 
    2.174095, 2.17008, 2.17915, 2.202158, 2.22184, 2.217941,
  2.232812, 2.227111, 2.20278, 2.176147, 2.157132, 2.149135, 2.149867, 
    2.149239, 2.13455, 2.095108, 2.031822, 1.962363, 1.92074, 1.900532, 
    1.88996, 1.881805, 1.875045, 1.867924, 1.86232, 1.867408, 1.882244, 
    1.896489, 1.908084, 1.922584, 1.931228, 1.95075, 1.986491, 2.017087, 
    2.064051, 2.161915, 2.263512, 2.319224, 2.353161, 2.40314, 2.443687, 
    2.45991, 2.455571, 2.436955, 2.412088, 2.394205, 2.393814, 2.393741, 
    2.377645, 2.357834, 2.342755, 2.33017, 2.327989, 2.338249, 2.345834, 
    2.341995, 2.337275, 2.349817, 2.38069, 2.407293, 2.402938,
  2.470685, 2.463491, 2.439658, 2.413851, 2.394994, 2.386079, 2.385047, 
    2.382657, 2.367616, 2.330318, 2.271535, 2.207192, 2.156793, 2.128691, 
    2.113884, 2.102265, 2.092398, 2.082206, 2.074337, 2.081417, 2.10261, 
    2.123352, 2.139921, 2.151768, 2.158428, 2.174891, 2.205877, 2.232195, 
    2.273372, 2.360077, 2.485239, 2.558431, 2.603101, 2.649511, 2.6839, 
    2.696504, 2.690703, 2.671876, 2.647449, 2.629312, 2.627106, 2.625048, 
    2.608459, 2.588505, 2.572664, 2.558929, 2.554845, 2.561926, 2.566595, 
    2.56131, 2.555359, 2.56504, 2.591306, 2.614019, 2.609205,
  2.777702, 2.768599, 2.739361, 2.707825, 2.684595, 2.673689, 2.672635, 
    2.669994, 2.651975, 2.606636, 2.534472, 2.461902, 2.415168, 2.388092, 
    2.372824, 2.360449, 2.349557, 2.338579, 2.329849, 2.334206, 2.351188, 
    2.367947, 2.381114, 2.390201, 2.394798, 2.414294, 2.453926, 2.487663, 
    2.540457, 2.651554, 2.766682, 2.829544, 2.867025, 2.905821, 2.933801, 
    2.94264, 2.93532, 2.916273, 2.892304, 2.873901, 2.869809, 2.865686, 
    2.848583, 2.82848, 2.811848, 2.796915, 2.790852, 2.794626, 2.79626, 
    2.789471, 2.782239, 2.788943, 2.814731, 2.843273, 2.837958,
  3.126121, 3.114862, 3.086569, 3.056649, 3.034028, 3.022257, 3.019199, 
    3.014598, 2.996742, 2.955314, 2.890603, 2.819581, 2.763133, 2.730248, 
    2.711544, 2.696202, 2.682492, 2.668855, 2.658162, 2.663394, 2.684532, 
    2.705767, 2.722679, 2.734467, 2.740576, 2.757565, 2.790396, 2.817911, 
    2.862178, 2.956329, 3.079495, 3.157583, 3.204017, 3.251844, 3.28626, 
    3.297092, 3.288067, 3.26444, 3.234653, 3.211627, 3.206038, 3.20041, 
    3.178867, 3.153419, 3.132253, 3.113181, 3.105234, 3.10917, 3.110424, 
    3.101766, 3.092754, 3.100756, 3.126651, 3.14938, 3.143456,
  3.562569, 3.549218, 3.515377, 3.479601, 3.452511, 3.438695, 3.435607, 
    3.430646, 3.409761, 3.360414, 3.282638, 3.197111, 3.129217, 3.098085, 
    3.0795, 3.063821, 3.049386, 3.035381, 3.024231, 3.026223, 3.041991, 
    3.06223, 3.083314, 3.098104, 3.105911, 3.126867, 3.166875, 3.200305, 
    3.253996, 3.367849, 3.484998, 3.54791, 3.583717, 3.620326, 3.645271, 
    3.650466, 3.639058, 3.614861, 3.585426, 3.561666, 3.553077, 3.544076, 
    3.521257, 3.494943, 3.471929, 3.450369, 3.439025, 3.437721, 3.434158, 
    3.422975, 3.411841, 3.415423, 3.438992, 3.465777, 3.459034,
  4.027123, 4.011809, 3.979948, 3.946856, 3.921209, 3.906726, 3.901307, 
    3.893916, 3.87341, 3.829443, 3.761646, 3.687244, 3.62719, 3.590841, 
    3.568585, 3.549593, 3.531611, 3.514603, 3.501431, 3.503037, 3.521334, 
    3.54054, 3.556393, 3.56709, 3.572065, 3.587643, 3.618568, 3.643682, 
    3.685838, 3.797944, 3.941083, 4.017117, 4.059662, 4.102912, 4.132073, 
    4.1375, 4.123122, 4.093083, 4.056584, 4.026787, 4.01547, 4.003168, 
    3.973814, 3.940041, 3.909906, 3.88119, 3.865419, 3.861233, 3.854099, 
    3.83882, 3.823724, 3.825751, 3.845733, 3.863506, 3.854541,
  4.739353, 4.720115, 4.676747, 4.630809, 4.595498, 4.575374, 4.567377, 
    4.556464, 4.527824, 4.467808, 4.376022, 4.276075, 4.195912, 4.147911, 
    4.118397, 4.092996, 4.06836, 4.045627, 4.028408, 4.028679, 4.050037, 
    4.072623, 4.091862, 4.104654, 4.110441, 4.128227, 4.164603, 4.193951, 
    4.243067, 4.350407, 4.459471, 4.51447, 4.562629, 4.616679, 4.653052, 
    4.660084, 4.642945, 4.605944, 4.560754, 4.523882, 4.510604, 4.495391, 
    4.457856, 4.414558, 4.375206, 4.337066, 4.31597, 4.308618, 4.296809, 
    4.275917, 4.255067, 4.254225, 4.274409, 4.291321, 4.277235,
  5.667004, 5.638623, 5.570301, 5.497511, 5.441764, 5.410233, 5.39759, 
    5.380997, 5.336496, 5.24355, 5.102967, 4.951191, 4.843627, 4.795535, 
    4.761826, 4.731114, 4.699252, 4.670823, 4.648688, 4.637187, 4.644199, 
    4.653993, 4.677014, 4.693133, 4.699999, 4.720981, 4.76586, 4.801814, 
    4.861277, 4.993551, 5.127173, 5.191073, 5.221136, 5.252059, 5.2693, 
    5.265387, 5.244418, 5.206267, 5.16182, 5.124152, 5.107722, 5.086539, 
    5.044455, 4.997392, 4.949953, 4.899971, 4.867649, 4.844581, 4.816351, 
    4.784966, 4.753425, 4.737539, 4.740246, 4.741514, 4.719381,
  6.845986, 6.801805, 6.695018, 6.591485, 6.527524, 6.482353, 6.451823, 
    6.418143, 6.362002, 6.267405, 6.135569, 5.993139, 5.87354, 5.793712, 
    5.733973, 5.677314, 5.617938, 5.56438, 5.52061, 5.488142, 5.482305, 
    5.481596, 5.484124, 5.482198, 5.475596, 5.476721, 5.498257, 5.514639, 
    5.548364, 5.717415, 5.889119, 5.96724, 6.001755, 6.038151, 6.056448, 
    6.050922, 6.027283, 5.980328, 5.927202, 5.884532, 5.871164, 5.84931, 
    5.797775, 5.739374, 5.675829, 5.604451, 5.559418, 5.523191, 5.476704, 
    5.429265, 5.379512, 5.347299, 5.338785, 5.326406, 5.283937,
  8.706301, 8.626128, 8.501668, 8.375813, 8.268732, 8.191971, 8.138944, 
    8.084408, 7.993335, 7.841672, 7.636763, 7.414307, 7.225255, 7.09516, 
    6.993039, 6.893236, 6.789722, 6.694379, 6.612947, 6.545221, 6.516981, 
    6.497747, 6.484987, 6.468534, 6.448538, 6.436758, 6.454144, 6.46679, 
    6.500868, 6.608283, 6.761753, 6.846615, 6.879406, 6.915448, 6.927709, 
    6.916493, 6.889322, 6.832495, 6.771884, 6.726917, 6.718995, 6.698018, 
    6.638669, 6.570779, 6.490485, 6.394669, 6.335154, 6.282547, 6.213968, 
    6.148376, 6.077744, 6.026026, 6.003721, 5.975298, 5.909097,
  10.9433, 10.80951, 10.62635, 10.44802, 10.29209, 10.17676, 10.09359, 
    10.01018, 9.880295, 9.674184, 9.403767, 9.109703, 8.854716, 8.670988, 
    8.518481, 8.365427, 8.207639, 8.059644, 7.928638, 7.811977, 7.748458, 
    7.699871, 7.662011, 7.622371, 7.581148, 7.548729, 7.553849, 7.55434, 
    7.580985, 7.694857, 7.805526, 7.836843, 7.850939, 7.870021, 7.860864, 
    7.837819, 7.80925, 7.746197, 7.683877, 7.642712, 7.646112, 7.628692, 
    7.562409, 7.487982, 7.390248, 7.266051, 7.188338, 7.113422, 7.016668, 
    6.930462, 6.836664, 6.760279, 6.716149, 6.664035, 6.571085,
  13.26865, 13.07509, 12.84066, 12.61999, 12.42007, 12.26519, 12.14684, 
    12.03006, 11.864, 11.61874, 11.30941, 10.97314, 10.6731, 10.44435, 
    10.24193, 10.03403, 9.819605, 9.616706, 9.432354, 9.256017, 9.140244, 
    9.047395, 8.973229, 8.902094, 8.83368, 8.772907, 8.751916, 8.725544, 
    8.73089, 8.822315, 8.901583, 8.899631, 8.862402, 8.842679, 8.819265, 
    8.792333, 8.771431, 8.707089, 8.64598, 8.613842, 8.642436, 8.633844, 
    8.554989, 8.472848, 8.353091, 8.190833, 8.085912, 7.982127, 7.852509, 
    7.742188, 7.622602, 7.522756, 7.461221, 7.388158, 7.26522,
  15.5616, 15.32258, 15.04983, 14.79587, 14.55958, 14.37186, 14.225, 
    14.08207, 13.88396, 13.59936, 13.24811, 12.8624, 12.50864, 12.23157, 
    11.97725, 11.71271, 11.43611, 11.17698, 10.94271, 10.7086, 10.54764, 
    10.42098, 10.32485, 10.23517, 10.151, 10.07558, 10.03917, 9.989581, 
    9.987998, 10.07692, 10.14049, 10.12388, 10.06882, 10.02547, 9.968823, 
    9.939071, 9.93482, 9.882603, 9.832075, 9.810094, 9.853036, 9.833669, 
    9.728488, 9.61712, 9.46461, 9.268003, 9.123292, 8.980047, 8.815855, 
    8.679338, 8.533298, 8.397584, 8.292372, 8.178309, 8.026809,
  17.45164, 17.20202, 16.9417, 16.70185, 16.47468, 16.28368, 16.12532, 
    15.96964, 15.76724, 15.49426, 15.17101, 14.80704, 14.44951, 14.1501, 
    13.85591, 13.5423, 13.20722, 12.8945, 12.61135, 12.30782, 12.09742, 
    11.94065, 11.84059, 11.748, 11.66047, 11.57792, 11.51837, 11.42835, 
    11.40171, 11.45193, 11.47281, 11.4352, 11.36722, 11.30887, 11.21104, 
    11.1482, 11.12104, 11.05964, 10.9851, 10.91042, 10.85925, 10.74456, 
    10.5621, 10.34902, 10.13103, 9.907432, 9.717621, 9.548362, 9.398157, 
    9.253122, 9.104719, 8.94649, 8.778739, 8.613841, 8.46542,
  18.12847, 17.87702, 17.65426, 17.46062, 17.27352, 17.10526, 16.95605, 
    16.80029, 16.63478, 16.45506, 16.25115, 16.02111, 15.76817, 15.53481, 
    15.28542, 15.01665, 14.72431, 14.44996, 14.1962, 13.90305, 13.67755, 
    13.49745, 13.38827, 13.26801, 13.13335, 12.99823, 12.85083, 12.66079, 
    12.52878, 12.42788, 12.31502, 12.20275, 12.06905, 11.96567, 11.84418, 
    11.74228, 11.6608, 11.56792, 11.44511, 11.29308, 11.14594, 10.95944, 
    10.73176, 10.49677, 10.24677, 9.981548, 9.742962, 9.520123, 9.31158, 
    9.114863, 8.932801, 8.766032, 8.593534, 8.436359, 8.29427,
  18.13201, 17.87243, 17.64789, 17.45793, 17.27298, 17.11142, 16.97334, 
    16.82544, 16.67529, 16.52282, 16.34147, 16.14457, 15.93243, 15.75931, 
    15.57972, 15.39363, 15.16566, 14.97122, 14.81032, 14.60521, 14.41923, 
    14.25222, 14.13235, 13.98, 13.79439, 13.60292, 13.37799, 13.11518, 
    12.89862, 12.68302, 12.46021, 12.28361, 12.13736, 12.02599, 11.89517, 
    11.78699, 11.70151, 11.6103, 11.49297, 11.34962, 11.21048, 11.02648, 
    10.7974, 10.56106, 10.3093, 10.04195, 9.797045, 9.565816, 9.348311, 
    9.143609, 8.955969, 8.785471, 8.608732, 8.448646, 8.30487,
  18.12733, 17.86117, 17.634, 17.44563, 17.26245, 17.10291, 16.96708, 
    16.82262, 16.67463, 16.52306, 16.34275, 16.14631, 15.9338, 15.76281, 
    15.58657, 15.4051, 15.17987, 14.99236, 14.84254, 14.64799, 14.47562, 
    14.32547, 14.21244, 14.06301, 13.87715, 13.67966, 13.44525, 13.17383, 
    12.9434, 12.71025, 12.47424, 12.29455, 12.1475, 12.03304, 11.90152, 
    11.79271, 11.70667, 11.61563, 11.49751, 11.3524, 11.21855, 11.03677, 
    10.80695, 10.56438, 10.30925, 10.04152, 9.796665, 9.566337, 9.350468, 
    9.145797, 8.958586, 8.788885, 8.613728, 8.454757, 8.311923,
  18.13222, 17.85781, 17.6272, 17.44033, 17.25713, 17.09849, 16.96443, 
    16.82264, 16.67643, 16.52574, 16.34665, 16.15062, 15.93784, 15.76755, 
    15.59194, 15.41099, 15.18639, 14.99924, 14.84956, 14.65542, 14.48486, 
    14.33787, 14.22597, 14.07606, 13.88806, 13.69137, 13.45909, 13.19114, 
    12.95835, 12.72328, 12.48538, 12.30394, 12.15538, 12.03993, 11.90741, 
    11.79875, 11.714, 11.62333, 11.50598, 11.362, 11.22769, 11.04526, 
    10.81465, 10.57186, 10.31632, 10.04802, 9.80168, 9.570178, 9.353488, 
    9.148674, 8.961405, 8.791698, 8.616179, 8.456951, 8.313994,
  18.14363, 17.86458, 17.63183, 17.44537, 17.26223, 17.10408, 16.97092, 
    16.83057, 16.68502, 16.53426, 16.35586, 16.16009, 15.94699, 15.77688, 
    15.60134, 15.42034, 15.19559, 15.00832, 14.85855, 14.66438, 14.49471, 
    14.34953, 14.23874, 14.08862, 13.89915, 13.70332, 13.47216, 13.20562, 
    12.9708, 12.73397, 12.49502, 12.31202, 12.16229, 12.04586, 11.91211, 
    11.80307, 11.71872, 11.62804, 11.51085, 11.36716, 11.23351, 11.0513, 
    10.82055, 10.57799, 10.32191, 10.05232, 9.804834, 9.572553, 9.355474, 
    9.150363, 8.962881, 8.793028, 8.617417, 8.458148, 8.315222 ;

 temp_east =
  6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388 ;

 temp_south =
  1.137725, 1.138182, 1.138384, 1.136393, 1.132912, 1.130674, 1.131729, 
    1.135111, 1.136749, 1.135931, 1.13423, 1.133517, 1.13501, 1.138603, 
    1.141014, 1.14102, 1.142408, 1.147855, 1.154208, 1.156471, 1.154765, 
    1.152558, 1.151241, 1.152298, 1.15877, 1.16726, 1.171243, 1.1717, 
    1.172055, 1.173003, 1.174874, 1.179693, 1.190464, 1.203298, 1.212377, 
    1.214597, 1.2127, 1.211963, 1.214853, 1.22064, 1.229518, 1.244212, 
    1.262913, 1.281232, 1.307438, 1.367511, 1.513266, 1.82348, 2.432452, 
    3.342487, 4.408576, 5.487299, 6.471881, 7.264916, 7.799684, 6.362131,
  1.165706, 1.166017, 1.166233, 1.16366, 1.160465, 1.158746, 1.160367, 
    1.163443, 1.166066, 1.165927, 1.164781, 1.164565, 1.166388, 1.172419, 
    1.176946, 1.17766, 1.180942, 1.189933, 1.199712, 1.203487, 1.20188, 
    1.199713, 1.198539, 1.200451, 1.209043, 1.219753, 1.224864, 1.225704, 
    1.226549, 1.228102, 1.230737, 1.236525, 1.246943, 1.259243, 1.272308, 
    1.275871, 1.273141, 1.272226, 1.27723, 1.28681, 1.300559, 1.322339, 
    1.34958, 1.371653, 1.396605, 1.469587, 1.628767, 1.983219, 2.650853, 
    3.643325, 4.72141, 5.78198, 6.729449, 7.509469, 8.102378, 6.362131,
  1.209825, 1.210234, 1.210571, 1.207738, 1.202207, 1.19935, 1.202391, 
    1.207945, 1.211415, 1.211739, 1.210021, 1.209774, 1.212744, 1.219301, 
    1.223822, 1.224745, 1.227965, 1.236448, 1.248246, 1.254406, 1.251541, 
    1.247748, 1.245944, 1.248543, 1.262547, 1.27984, 1.287897, 1.288976, 
    1.29, 1.292193, 1.296133, 1.30512, 1.321401, 1.340503, 1.354006, 
    1.357679, 1.355576, 1.355158, 1.360166, 1.369371, 1.382349, 1.40276, 
    1.434402, 1.466192, 1.502232, 1.581819, 1.778316, 2.186081, 2.956237, 
    3.982757, 5.061129, 6.077973, 6.978192, 7.718756, 8.361522, 6.362131,
  1.26423, 1.264692, 1.265058, 1.259894, 1.250233, 1.245211, 1.250424, 
    1.260298, 1.265997, 1.265719, 1.262609, 1.261977, 1.26678, 1.277371, 
    1.284684, 1.286108, 1.291444, 1.305507, 1.320661, 1.326621, 1.324298, 
    1.321144, 1.31948, 1.322582, 1.335856, 1.352181, 1.360012, 1.361424, 
    1.362793, 1.365236, 1.369285, 1.377985, 1.393389, 1.418144, 1.438241, 
    1.443093, 1.439158, 1.438009, 1.44489, 1.457825, 1.476312, 1.505657, 
    1.54213, 1.571423, 1.604746, 1.695164, 1.923207, 2.392361, 3.218716, 
    4.274543, 5.353222, 6.337874, 7.214526, 7.969189, 8.584683, 6.362131,
  1.327183, 1.327663, 1.328074, 1.32339, 1.314465, 1.309901, 1.314873, 
    1.324059, 1.329634, 1.32993, 1.327284, 1.326972, 1.331728, 1.341991, 
    1.349106, 1.350658, 1.355819, 1.369097, 1.390156, 1.399619, 1.395064, 
    1.389111, 1.385681, 1.390132, 1.411254, 1.437095, 1.448828, 1.450038, 
    1.451148, 1.453962, 1.459299, 1.471947, 1.494994, 1.5218, 1.540275, 
    1.544628, 1.540832, 1.5396, 1.545844, 1.557736, 1.574737, 1.601812, 
    1.63551, 1.670751, 1.722917, 1.838474, 2.061069, 2.571187, 3.446288, 
    4.527568, 5.606569, 6.563367, 7.419657, 8.199811, 8.796298, 6.362131,
  1.405654, 1.406129, 1.40648, 1.397901, 1.3822, 1.373995, 1.382336, 
    1.398471, 1.407441, 1.406358, 1.401209, 1.400019, 1.407494, 1.423941, 
    1.435254, 1.437355, 1.445671, 1.467543, 1.49083, 1.49966, 1.495461, 
    1.489949, 1.48679, 1.490939, 1.51056, 1.534577, 1.545474, 1.546578, 
    1.547593, 1.550171, 1.555072, 1.566753, 1.588061, 1.612827, 1.629877, 
    1.633792, 1.630119, 1.628815, 1.634499, 1.645475, 1.671446, 1.713923, 
    1.766824, 1.809097, 1.857226, 1.964329, 2.255098, 2.793112, 3.704057, 
    4.787533, 5.835542, 6.761582, 7.600052, 8.402729, 9.075432, 6.362131,
  1.499188, 1.499637, 1.499991, 1.492049, 1.477425, 1.469839, 1.47772, 
    1.492809, 1.501397, 1.500795, 1.49618, 1.495268, 1.50244, 1.518072, 
    1.528814, 1.530868, 1.538694, 1.559143, 1.580907, 1.589173, 1.585291, 
    1.580175, 1.577258, 1.581137, 1.599414, 1.621801, 1.634639, 1.635241, 
    1.635659, 1.638647, 1.64545, 1.663382, 1.697106, 1.736448, 1.763034, 
    1.768153, 1.760943, 1.75774, 1.765713, 1.782043, 1.806092, 1.845159, 
    1.893921, 1.932888, 1.977405, 2.109954, 2.428721, 3.03058, 3.973792, 
    5.056771, 6.076018, 6.965693, 7.772936, 8.584635, 9.325778, 6.362131,
  1.58502, 1.585445, 1.585802, 1.578444, 1.564809, 1.557791, 1.565249, 
    1.579379, 1.587617, 1.587456, 1.583332, 1.582674, 1.589568, 1.604452, 
    1.615917, 1.618692, 1.631128, 1.66436, 1.699567, 1.712496, 1.705131, 
    1.695626, 1.689764, 1.695107, 1.724235, 1.760019, 1.775463, 1.775752, 
    1.775876, 1.778363, 1.784369, 1.800728, 1.831761, 1.867983, 1.892355, 
    1.896677, 1.889469, 1.885969, 1.892924, 1.907707, 1.929654, 1.965592, 
    2.010558, 2.057271, 2.129516, 2.29151, 2.588063, 3.248526, 4.221376, 
    5.303934, 6.29682, 7.169565, 7.99302, 8.785998, 9.555973, 6.362131,
  1.719404, 1.720013, 1.720471, 1.708207, 1.685907, 1.674212, 1.686169, 
    1.709665, 1.722464, 1.720356, 1.712921, 1.711074, 1.721604, 1.744812, 
    1.760733, 1.763491, 1.775244, 1.806302, 1.839136, 1.851188, 1.844278, 
    1.835314, 1.829754, 1.834581, 1.861509, 1.894648, 1.908798, 1.90879, 
    1.908637, 1.910647, 1.915899, 1.93077, 1.959256, 1.992523, 2.0148, 
    2.018367, 2.011161, 2.00738, 2.013371, 2.026688, 2.056901, 2.114935, 
    2.187974, 2.246457, 2.313216, 2.463415, 2.808861, 3.4549, 4.455829, 
    5.538011, 6.505959, 7.362701, 8.201565, 9.03666, 9.774223, 6.362131,
  1.859259, 1.86008, 1.860779, 1.849692, 1.829283, 1.818748, 1.830189, 
    1.852338, 1.864672, 1.863287, 1.856777, 1.855436, 1.865564, 1.887549, 
    1.902639, 1.90538, 1.916464, 1.945391, 1.9759, 1.987093, 1.980628, 
    1.972195, 1.966932, 1.971252, 1.996025, 2.026571, 2.043029, 2.042264, 
    2.041235, 2.043578, 2.051014, 2.073558, 2.117733, 2.169905, 2.205039, 
    2.210826, 2.199569, 2.193844, 2.203498, 2.224735, 2.257083, 2.310641, 
    2.377981, 2.431843, 2.493227, 2.631869, 3.05755, 3.719573, 4.701493, 
    5.767407, 6.710926, 7.551998, 8.405982, 9.28239, 10.04145, 6.362131,
  2.003505, 2.004563, 2.005414, 1.99286, 1.974366, 1.965004, 1.975923, 
    1.996709, 2.009722, 2.00792, 2.002346, 2.001517, 2.011237, 2.038685, 
    2.060117, 2.063778, 2.079874, 2.122417, 2.167399, 2.183944, 2.1741, 
    2.161202, 2.152963, 2.159129, 2.196303, 2.242378, 2.261855, 2.261346, 
    2.260591, 2.262924, 2.269928, 2.29083, 2.331614, 2.379722, 2.412181, 
    2.417554, 2.407174, 2.40185, 2.410625, 2.430005, 2.459647, 2.508676, 
    2.570248, 2.619435, 2.698372, 2.912108, 3.309196, 4.027651, 5.016097, 
    6.044277, 6.943497, 7.743524, 8.612796, 9.530982, 10.36816, 6.362131,
  2.230664, 2.232634, 2.234447, 2.220813, 2.195125, 2.182148, 2.197968, 
    2.228413, 2.245332, 2.243423, 2.235397, 2.234097, 2.247994, 2.277509, 
    2.298074, 2.30231, 2.317924, 2.357501, 2.399158, 2.414903, 2.406487, 
    2.395177, 2.388108, 2.394099, 2.428281, 2.470566, 2.488573, 2.488327, 
    2.487858, 2.49018, 2.496737, 2.515937, 2.553208, 2.597105, 2.626792, 
    2.631735, 2.622265, 2.617355, 2.62522, 2.642675, 2.684169, 2.757494, 
    2.850536, 2.925912, 3.012195, 3.207489, 3.587621, 4.346819, 5.342011, 
    6.335494, 7.213331, 8.040564, 8.912197, 9.805355, 10.70634, 6.362131,
  2.468373, 2.471299, 2.474118, 2.463098, 2.441331, 2.430979, 2.446493, 
    2.475259, 2.491886, 2.491608, 2.48573, 2.48585, 2.499577, 2.527426, 
    2.547083, 2.551922, 2.567031, 2.603503, 2.645837, 2.666411, 2.655546, 
    2.640774, 2.634174, 2.639982, 2.684534, 2.740911, 2.765347, 2.765538, 
    2.765361, 2.769047, 2.778631, 2.805741, 2.858286, 2.920892, 2.964169, 
    2.973288, 2.962248, 2.957805, 2.971434, 2.9989, 3.040442, 3.108072, 
    3.193079, 3.262126, 3.340585, 3.51658, 3.997321, 4.695258, 5.683018, 
    6.640173, 7.495608, 8.351404, 9.262537, 10.22426, 11.06809, 6.362131,
  2.775254, 2.779672, 2.784018, 2.77147, 2.745847, 2.734077, 2.754019, 
    2.790606, 2.811889, 2.811861, 2.805426, 2.806373, 2.824271, 2.859663, 
    2.88519, 2.892429, 2.912751, 2.960216, 3.010082, 3.030675, 3.02341, 
    3.012577, 3.006477, 3.015513, 3.057588, 3.109378, 3.133093, 3.135522, 
    3.137541, 3.143084, 3.153944, 3.180374, 3.22936, 3.287339, 3.328133, 
    3.338824, 3.331762, 3.330652, 3.345312, 3.372008, 3.411086, 3.47279, 
    3.558218, 3.650306, 3.755005, 3.988556, 4.423535, 5.165606, 6.09266, 
    6.996017, 7.815896, 8.674664, 9.626812, 10.65975, 11.66256, 6.362131,
  3.123553, 3.129791, 3.136136, 3.128056, 3.108782, 3.101575, 3.121865, 
    3.156694, 3.178366, 3.181692, 3.1794, 3.183481, 3.202199, 3.236127, 
    3.261395, 3.270723, 3.291454, 3.335423, 3.38126, 3.401871, 3.398275, 
    3.391456, 3.38866, 3.398934, 3.437741, 3.500865, 3.531155, 3.535822, 
    3.539897, 3.548445, 3.563721, 3.598422, 3.661511, 3.736429, 3.790205, 
    3.8067, 3.801041, 3.802887, 3.824474, 3.861236, 3.914239, 3.996464, 
    4.098387, 4.181884, 4.275257, 4.478927, 4.936018, 5.644892, 6.531266, 
    7.40376, 8.266735, 9.182453, 10.16327, 11.23174, 12.26808, 6.362131,
  3.559371, 3.566236, 3.573528, 3.564031, 3.541496, 3.533623, 3.558326, 
    3.600006, 3.626099, 3.630694, 3.629312, 3.635511, 3.658893, 3.69966, 
    3.730718, 3.743618, 3.769793, 3.823179, 3.878962, 3.905475, 3.903848, 
    3.898553, 3.897835, 3.912715, 3.961576, 4.020358, 4.05112, 4.060624, 
    4.06948, 4.082493, 4.101565, 4.137229, 4.197176, 4.26742, 4.319611, 
    4.34041, 4.342594, 4.351131, 4.375947, 4.413188, 4.464504, 4.539906, 
    4.638551, 4.736447, 4.845198, 5.079516, 5.515961, 6.190895, 7.00843, 
    7.845764, 8.71637, 9.697616, 10.75014, 11.92687, 13.15105, 6.362131,
  4.023047, 4.029872, 4.037664, 4.032213, 4.015967, 4.012455, 4.036463, 
    4.074482, 4.100077, 4.108368, 4.111835, 4.121824, 4.146258, 4.184961, 
    4.215768, 4.231707, 4.26323, 4.32759, 4.394132, 4.426051, 4.425545, 
    4.421236, 4.422199, 4.441267, 4.498895, 4.567091, 4.604054, 4.617737, 
    4.63056, 4.648496, 4.673636, 4.717285, 4.788167, 4.870829, 4.933372, 
    4.961412, 4.969079, 4.983637, 5.015996, 5.061903, 5.124087, 5.212988, 
    5.319801, 5.4075, 5.502632, 5.699885, 6.13031, 6.736045, 7.529856, 
    8.4266, 9.38745, 10.4462, 11.57716, 12.86807, 14.03904, 6.362131,
  4.731818, 4.729474, 4.728772, 4.710695, 4.679104, 4.665576, 4.68854, 
    4.728903, 4.753281, 4.75628, 4.754199, 4.760984, 4.785933, 4.827145, 
    4.859312, 4.874547, 4.902368, 4.956232, 5.012157, 5.040356, 5.042826, 
    5.042685, 5.046318, 5.065531, 5.116842, 5.176202, 5.211574, 5.229381, 
    5.246142, 5.26812, 5.297007, 5.341149, 5.408052, 5.485229, 5.555233, 
    5.589716, 5.603641, 5.624604, 5.663303, 5.715194, 5.78367, 5.878008, 
    5.989368, 6.080557, 6.178076, 6.37532, 6.739357, 7.351928, 8.156037, 
    9.103111, 10.12504, 11.30526, 12.54121, 13.8473, 14.78033, 6.362131,
  5.654085, 5.635841, 5.619353, 5.574149, 5.508645, 5.472019, 5.492241, 
    5.538878, 5.559791, 5.547891, 5.529426, 5.524851, 5.547047, 5.59123, 
    5.622309, 5.630002, 5.654542, 5.713303, 5.773098, 5.795901, 5.78617, 
    5.774291, 5.766546, 5.779283, 5.830976, 5.889112, 5.920285, 5.933342, 
    5.94409, 5.962238, 5.989429, 6.033558, 6.102273, 6.182201, 6.243049, 
    6.276548, 6.294965, 6.319735, 6.358727, 6.408343, 6.471225, 6.554618, 
    6.651519, 6.731448, 6.833633, 7.038347, 7.409668, 8.002745, 8.841807, 
    9.850951, 11.00345, 12.37914, 13.7103, 14.66776, 15.25131, 6.362131,
  6.825705, 6.784884, 6.745215, 6.657738, 6.551785, 6.500284, 6.493831, 
    6.536307, 6.552302, 6.514031, 6.465552, 6.439486, 6.456486, 6.508171, 
    6.538617, 6.531691, 6.551089, 6.623561, 6.696102, 6.710097, 6.67386, 
    6.634889, 6.601985, 6.600122, 6.654526, 6.714507, 6.735937, 6.733276, 
    6.726251, 6.730362, 6.74739, 6.786654, 6.8566, 6.940003, 6.996095, 
    7.020706, 7.029712, 7.048966, 7.085302, 7.134202, 7.193902, 7.275466, 
    7.370947, 7.450445, 7.533594, 7.695278, 8.136338, 8.724344, 9.722831, 
    10.88957, 12.28071, 13.77767, 14.58697, 15.10489, 15.33883, 6.362131,
  8.676331, 8.608376, 8.539832, 8.433104, 8.304549, 8.208417, 8.179864, 
    8.187611, 8.163034, 8.097162, 8.023645, 7.968942, 7.94891, 7.953301, 
    7.942251, 7.903368, 7.88291, 7.902439, 7.921252, 7.895268, 7.830635, 
    7.763826, 7.698774, 7.660699, 7.668969, 7.718703, 7.723687, 7.691364, 
    7.652077, 7.629579, 7.626449, 7.657026, 7.732832, 7.827184, 7.878469, 
    7.884169, 7.868409, 7.870127, 7.89729, 7.942814, 7.997199, 8.080375, 
    8.180965, 8.26543, 8.356091, 8.544676, 8.96311, 9.693784, 10.8238, 
    12.23919, 13.83795, 14.70637, 15.09966, 15.2543, 15.39415, 6.362131,
  10.92399, 10.83996, 10.75409, 10.61665, 10.45015, 10.32155, 10.28032, 
    10.29243, 10.25724, 10.16041, 10.05142, 9.965725, 9.926834, 9.92351, 
    9.895668, 9.824353, 9.778626, 9.790584, 9.800008, 9.739864, 9.61881, 
    9.491419, 9.369802, 9.284813, 9.26566, 9.250607, 9.194576, 9.114146, 
    9.027782, 8.958961, 8.909637, 8.887584, 8.905754, 8.968117, 9.005085, 
    8.978707, 8.921509, 8.889716, 8.895304, 8.92767, 8.967892, 9.048437, 
    9.152912, 9.239635, 9.336679, 9.561757, 9.948263, 10.8682, 12.25342, 
    13.91332, 14.9101, 15.25205, 15.28985, 15.31477, 15.39543, 6.362131,
  13.22495, 13.13683, 13.04867, 12.91038, 12.74402, 12.61235, 12.56806, 
    12.58444, 12.54989, 12.44701, 12.32939, 12.23364, 12.18714, 12.18177, 
    12.14537, 12.05451, 11.99357, 11.9972, 11.99448, 11.90833, 11.74232, 
    11.56244, 11.39048, 11.26031, 11.21018, 11.17085, 11.0746, 10.94132, 
    10.80877, 10.69739, 10.61003, 10.54954, 10.54184, 10.55937, 10.53547, 
    10.46308, 10.36661, 10.28895, 10.24202, 10.21789, 10.19721, 10.26381, 
    10.37122, 10.45297, 10.54988, 10.81393, 11.28141, 12.4463, 14.02154, 
    15.09322, 15.44468, 15.45423, 15.36075, 15.31665, 15.39645, 6.362131,
  15.41727, 15.33184, 15.24888, 15.12285, 14.97406, 14.8564, 14.81769, 
    14.83826, 14.81202, 14.72286, 14.6199, 14.53572, 14.49638, 14.49448, 
    14.45982, 14.3693, 14.30679, 14.30162, 14.2856, 14.18803, 14.00346, 
    13.79755, 13.5968, 13.43731, 13.36215, 13.30228, 13.17824, 13.00948, 
    12.84982, 12.7142, 12.60633, 12.51732, 12.49223, 12.4991, 12.47151, 
    12.37769, 12.24579, 12.1202, 12.02423, 11.94759, 11.89746, 11.91404, 
    12.02984, 12.09692, 12.18638, 12.50062, 13.13151, 14.41508, 15.25544, 
    15.59802, 15.5279, 15.53223, 15.36277, 15.31859, 15.39933, 6.362131,
  17.43805, 17.34934, 17.26926, 17.15983, 17.03227, 16.93411, 16.90556, 
    16.92876, 16.91301, 16.84423, 16.76402, 16.70317, 16.68408, 16.69323, 
    16.67365, 16.60501, 16.55723, 16.556, 16.54273, 16.45448, 16.27988, 
    16.07794, 15.87887, 15.71602, 15.63264, 15.56236, 15.42803, 15.24689, 
    15.07974, 14.94061, 14.83362, 14.73314, 14.70732, 14.72491, 14.72071, 
    14.64433, 14.52396, 14.39307, 14.2796, 14.17314, 14.14381, 14.19883, 
    14.29797, 14.31398, 14.35317, 14.63349, 15.32299, 15.51612, 15.70623, 
    15.61771, 15.55661, 15.53383, 15.36544, 15.32123, 15.40181, 6.362131,
  18.46674, 18.38478, 18.32462, 18.27884, 18.23628, 18.2035, 18.19345, 
    18.21174, 18.2217, 18.21494, 18.19625, 18.17925, 18.17432, 18.18985, 
    18.17809, 18.12812, 18.09666, 18.073, 18.0309, 17.96367, 17.85676, 
    17.7364, 17.61612, 17.51555, 17.46651, 17.44406, 17.36345, 17.22886, 
    17.12918, 17.04239, 16.97243, 16.89222, 16.87627, 16.862, 16.81468, 
    16.75378, 16.68421, 16.59544, 16.49002, 16.367, 16.28489, 16.20102, 
    16.11257, 15.982, 15.86, 15.7891, 15.81909, 15.78021, 15.72757, 15.62274, 
    15.55677, 15.53797, 15.36889, 15.32333, 15.40379, 6.362131,
  18.56439, 18.48776, 18.43825, 18.41583, 18.40644, 18.40457, 18.41039, 
    18.43452, 18.45905, 18.48383, 18.49822, 18.50162, 18.49413, 18.4998, 
    18.47771, 18.42782, 18.39054, 18.32838, 18.24127, 18.16463, 18.08672, 
    18.00745, 17.9195, 17.83784, 17.76353, 17.69782, 17.6235, 17.53977, 
    17.48783, 17.43656, 17.38659, 17.30225, 17.23205, 17.16429, 17.10471, 
    17.03232, 16.9475, 16.85597, 16.74913, 16.62687, 16.52385, 16.41378, 
    16.2966, 16.18176, 16.0742, 15.97372, 15.86683, 15.78596, 15.73092, 
    15.62228, 15.56341, 15.54358, 15.37166, 15.32503, 15.40507, 6.362131,
  18.56682, 18.4896, 18.43977, 18.41729, 18.40868, 18.40757, 18.41398, 
    18.4385, 18.46328, 18.4883, 18.50346, 18.50693, 18.49874, 18.50405, 
    18.48143, 18.43085, 18.39323, 18.33077, 18.24341, 18.16681, 18.08883, 
    18.00956, 17.92193, 17.84068, 17.76571, 17.70035, 17.63225, 17.56135, 
    17.51623, 17.46998, 17.42261, 17.33675, 17.25944, 17.19061, 17.13217, 
    17.05711, 16.96568, 16.8631, 16.7505, 16.62783, 16.52319, 16.41218, 
    16.29447, 16.17921, 16.07207, 15.97412, 15.86927, 15.7886, 15.73543, 
    15.63366, 15.57111, 15.54811, 15.37336, 15.32532, 15.40507, 6.362131,
  18.56869, 18.49128, 18.44132, 18.41879, 18.41065, 18.40975, 18.41612, 
    18.4408, 18.46564, 18.49062, 18.50571, 18.50919, 18.50107, 18.50633, 
    18.48349, 18.43256, 18.39487, 18.33225, 18.2447, 18.1678, 18.08956, 
    18.00998, 17.92256, 17.84109, 17.76559, 17.70078, 17.63503, 17.56833, 
    17.52598, 17.48238, 17.43756, 17.35431, 17.27978, 17.21395, 17.15663, 
    17.08309, 16.99341, 16.8905, 16.77555, 16.64847, 16.53767, 16.42376, 
    16.30647, 16.18832, 16.08139, 15.98657, 15.88291, 15.8047, 15.74949, 
    15.64337, 15.57577, 15.54919, 15.37336, 15.32532, 15.40507, 6.362131,
  18.57084, 18.49343, 18.44355, 18.42121, 18.41377, 18.41334, 18.41993, 
    18.44501, 18.46999, 18.49488, 18.50983, 18.5131, 18.50468, 18.50966, 
    18.48657, 18.43541, 18.39758, 18.335, 18.24765, 18.17071, 18.09252, 
    18.01309, 17.92582, 17.84477, 17.76995, 17.70571, 17.64106, 17.57603, 
    17.53505, 17.49298, 17.4498, 17.36823, 17.29499, 17.23006, 17.17284, 
    17.10078, 17.01387, 16.91422, 16.80184, 16.67673, 16.56829, 16.45516, 
    16.33733, 16.21971, 16.11059, 16.00998, 15.90179, 15.81669, 15.75466, 
    15.64426, 15.57577, 15.54919, 15.37336, 15.32532, 15.40507, 6.362131,
  1.137597, 1.138018, 1.138191, 1.136186, 1.132701, 1.130463, 1.131499, 
    1.134864, 1.136471, 1.135619, 1.133947, 1.133227, 1.13466, 1.138188, 
    1.140541, 1.140517, 1.141952, 1.147436, 1.153836, 1.156112, 1.154414, 
    1.152205, 1.150917, 1.151995, 1.158491, 1.167025, 1.171035, 1.171498, 
    1.171871, 1.172834, 1.174714, 1.179529, 1.190255, 1.203009, 1.21202, 
    1.214122, 1.212068, 1.211227, 1.214079, 1.219915, 1.228828, 1.243573, 
    1.262396, 1.281049, 1.307569, 1.368257, 1.517208, 1.832797, 2.444176, 
    3.363557, 4.442914, 5.527749, 6.504662, 7.282581, 7.80057, 6.262388,
  1.165555, 1.165814, 1.165973, 1.163343, 1.160117, 1.158357, 1.159909, 
    1.162962, 1.165497, 1.165211, 1.164087, 1.163853, 1.165602, 1.171562, 
    1.176048, 1.176759, 1.18024, 1.189355, 1.199199, 1.203006, 1.201438, 
    1.199297, 1.198188, 1.200136, 1.208732, 1.21947, 1.224604, 1.225458, 
    1.226341, 1.227916, 1.230556, 1.236311, 1.246657, 1.258842, 1.271813, 
    1.275193, 1.272192, 1.271127, 1.276131, 1.285872, 1.299766, 1.321747, 
    1.349313, 1.372066, 1.397585, 1.471955, 1.635584, 1.994388, 2.664046, 
    3.666072, 4.757276, 5.82129, 6.757092, 7.523089, 8.094893, 6.262388,
  1.209679, 1.210008, 1.210261, 1.207346, 1.201764, 1.198847, 1.201806, 
    1.20735, 1.210704, 1.210813, 1.20912, 1.208848, 1.211737, 1.218197, 
    1.222663, 1.22359, 1.227046, 1.235675, 1.247549, 1.253761, 1.250949, 
    1.247195, 1.245472, 1.248123, 1.262155, 1.279511, 1.287614, 1.288711, 
    1.289791, 1.292014, 1.295961, 1.304908, 1.321112, 1.340091, 1.353479, 
    1.356942, 1.354541, 1.353953, 1.358985, 1.368418, 1.381563, 1.40226, 
    1.434384, 1.467181, 1.504384, 1.586506, 1.787249, 2.197809, 2.970273, 
    4.00741, 5.095804, 6.112701, 7.001682, 7.728916, 8.34687, 6.262388,
  1.264199, 1.264554, 1.264809, 1.259522, 1.249771, 1.244661, 1.249794, 
    1.259688, 1.265245, 1.264664, 1.261569, 1.260897, 1.265596, 1.276049, 
    1.283286, 1.284717, 1.290332, 1.30457, 1.319812, 1.32585, 1.323602, 
    1.320504, 1.318947, 1.322123, 1.335441, 1.351855, 1.359744, 1.361181, 
    1.362622, 1.365103, 1.369157, 1.377804, 1.393114, 1.417739, 1.43771, 
    1.44233, 1.438069, 1.436737, 1.443674, 1.456918, 1.475602, 1.505327, 
    1.542415, 1.573003, 1.608085, 1.701705, 1.933848, 2.404075, 3.233474, 
    4.300835, 5.386873, 6.368226, 7.234628, 7.973103, 8.56386, 6.262388,
  1.327358, 1.327705, 1.327979, 1.323148, 1.31413, 1.309466, 1.314338, 
    1.323548, 1.328932, 1.328823, 1.326169, 1.325787, 1.330402, 1.340477, 
    1.347492, 1.349054, 1.354538, 1.368018, 1.389176, 1.39874, 1.39428, 
    1.388397, 1.385097, 1.389642, 1.410829, 1.436794, 1.448608, 1.449849, 
    1.451049, 1.453911, 1.459255, 1.471848, 1.494802, 1.521466, 1.53979, 
    1.543887, 1.539742, 1.538329, 1.544669, 1.556945, 1.574144, 1.601648, 
    1.636058, 1.672827, 1.727164, 1.846255, 2.072884, 2.582891, 3.461674, 
    4.55528, 5.639332, 6.589921, 7.436819, 8.197685, 8.769197, 6.262388,
  1.406091, 1.40641, 1.406605, 1.397844, 1.38202, 1.373689, 1.381931, 
    1.398125, 1.40687, 1.405275, 1.400083, 1.398788, 1.40609, 1.422307, 
    1.433499, 1.435604, 1.444272, 1.466361, 1.489738, 1.498692, 1.494608, 
    1.489188, 1.486181, 1.490447, 1.510155, 1.534322, 1.545317, 1.546462, 
    1.547588, 1.550224, 1.555131, 1.566747, 1.587948, 1.612555, 1.629433, 
    1.633071, 1.629028, 1.627544, 1.63336, 1.644787, 1.67094, 1.713857, 
    1.767523, 1.811513, 1.862147, 1.973199, 2.26612, 2.804435, 3.720417, 
    4.815454, 5.867069, 6.784798, 7.614628, 8.39529, 9.037982, 6.262388,
  1.49994, 1.500215, 1.500398, 1.492261, 1.477522, 1.46981, 1.477579, 
    1.492728, 1.50104, 1.499822, 1.495136, 1.49408, 1.501035, 1.516373, 
    1.526958, 1.529011, 1.537201, 1.55787, 1.579716, 1.588125, 1.584376, 
    1.579371, 1.576627, 1.580643, 1.599027, 1.621587, 1.634541, 1.635193, 
    1.635739, 1.638796, 1.64561, 1.663483, 1.697117, 1.736313, 1.762722, 
    1.767531, 1.759898, 1.756491, 1.764601, 1.781416, 1.805599, 1.845127, 
    1.894742, 1.935607, 1.982929, 2.119037, 2.439036, 3.041344, 3.991312, 
    5.083873, 6.10389, 6.985999, 7.784726, 8.572433, 9.279046, 6.262388,
  1.586061, 1.586297, 1.586467, 1.578904, 1.565161, 1.558015, 1.565351, 
    1.579542, 1.587456, 1.586584, 1.582361, 1.581526, 1.588162, 1.602693, 
    1.613969, 1.616733, 1.62954, 1.66297, 1.69822, 1.711301, 1.704098, 
    1.694739, 1.689075, 1.69458, 1.723839, 1.759833, 1.775432, 1.775806, 
    1.776103, 1.778688, 1.784721, 1.801027, 1.831958, 1.868008, 1.892178, 
    1.896154, 1.888475, 1.884743, 1.891838, 1.907136, 1.929173, 1.965593, 
    2.01149, 2.060178, 2.134985, 2.299688, 2.597727, 3.258776, 4.23996, 
    5.330285, 6.321336, 7.187245, 7.999654, 8.767658, 9.500708, 6.262388,
  1.720763, 1.721174, 1.721439, 1.708959, 1.68655, 1.674723, 1.686555, 
    1.710124, 1.72255, 1.719625, 1.712048, 1.709978, 1.720201, 1.742978, 
    1.75866, 1.761389, 1.773498, 1.804738, 1.837594, 1.849816, 1.843093, 
    1.834306, 1.82897, 1.833992, 1.861096, 1.894487, 1.90883, 1.90894, 
    1.909002, 1.911139, 1.916435, 1.931255, 1.959629, 1.9927, 2.01475, 
    2.017937, 2.010214, 2.006176, 2.012308, 2.02617, 2.056407, 2.114846, 
    2.188704, 2.248944, 2.318061, 2.470736, 2.817445, 3.464663, 4.475421, 
    5.56365, 6.527296, 7.377894, 8.203314, 9.009392, 9.710866, 6.262388,
  1.860936, 1.861552, 1.862052, 1.850747, 1.830245, 1.819583, 1.830892, 
    1.853107, 1.865013, 1.862703, 1.856009, 1.854397, 1.864164, 1.885641, 
    1.900443, 1.903138, 1.914563, 1.943656, 1.974166, 1.985547, 1.979294, 
    1.971068, 1.966053, 1.970603, 1.995594, 2.026435, 2.043119, 2.042509, 
    2.041735, 2.044236, 2.051734, 2.074246, 2.118328, 2.170315, 2.205235, 
    2.210612, 2.198771, 2.192724, 2.202458, 2.224158, 2.256403, 2.310298, 
    2.378441, 2.433919, 2.497459, 2.638349, 3.064867, 3.729048, 4.721726, 
    5.792349, 6.729147, 7.564753, 8.402943, 9.246367, 9.967228, 6.262388,
  2.005498, 2.006345, 2.006992, 1.994223, 1.975651, 1.966167, 1.976947, 
    1.997792, 2.010318, 2.007486, 2.001685, 2.000536, 2.009842, 2.036703, 
    2.057802, 2.061396, 2.077808, 2.120479, 2.16542, 2.182149, 2.172538, 
    2.159887, 2.151919, 2.158349, 2.195781, 2.242186, 2.261951, 2.261669, 
    2.261243, 2.263794, 2.270911, 2.291819, 2.332517, 2.380415, 2.412651, 
    2.417579, 2.406552, 2.400834, 2.409608, 2.429361, 2.45878, 2.508077, 
    2.570435, 2.621095, 2.701841, 2.91706, 3.315232, 4.036963, 5.03555, 
    6.065835, 6.958494, 7.753812, 8.604912, 9.486106, 10.27982, 6.262388,
  2.232812, 2.234587, 2.23621, 2.22238, 2.196642, 2.18356, 2.199239, 
    2.229708, 2.246103, 2.243121, 2.234832, 2.233176, 2.246622, 2.275488, 
    2.295671, 2.299805, 2.315662, 2.355312, 2.396892, 2.412817, 2.404646, 
    2.393615, 2.386831, 2.393127, 2.427637, 2.470312, 2.488674, 2.488732, 
    2.488666, 2.491271, 2.497993, 2.517238, 2.554429, 2.598091, 2.627546, 
    2.632007, 2.621824, 2.616447, 2.624227, 2.641963, 2.683071, 2.756485, 
    2.850081, 2.926522, 3.014261, 3.210829, 3.592354, 4.355962, 5.360657, 
    6.353284, 7.224905, 8.045053, 8.895041, 9.750486, 10.60339, 6.262388,
  2.470685, 2.473429, 2.476074, 2.464873, 2.44307, 2.432625, 2.448003, 
    2.476772, 2.49284, 2.491445, 2.485266, 2.484993, 2.498231, 2.525363, 
    2.544587, 2.549287, 2.564562, 2.601052, 2.643262, 2.663996, 2.653396, 
    2.638951, 2.632652, 2.638809, 2.683728, 2.740517, 2.765376, 2.765973, 
    2.766297, 2.770353, 2.780178, 2.807398, 2.859889, 2.922238, 2.965314, 
    2.973922, 2.962078, 2.957027, 2.970388, 2.9979, 3.038818, 3.106339, 
    3.19174, 3.261556, 3.341184, 3.518232, 4.000907, 4.703981, 5.700819, 
    6.65402, 7.503601, 8.349818, 9.233802, 10.15233, 10.95083, 6.262388,
  2.777702, 2.781951, 2.786133, 2.773421, 2.747775, 2.735923, 2.755733, 
    2.792271, 2.812954, 2.811778, 2.80501, 2.80553, 2.822903, 2.857494, 
    2.882518, 2.889563, 2.909917, 2.957285, 3.006957, 3.027658, 3.02064, 
    3.010153, 3.004359, 3.013792, 3.05634, 3.108633, 3.132889, 3.135875, 
    3.138536, 3.144582, 3.155809, 3.182442, 3.231398, 3.289078, 3.329697, 
    3.339845, 3.331885, 3.330011, 3.344204, 3.370705, 3.408915, 3.470305, 
    3.555932, 3.648391, 3.754011, 3.988972, 4.425929, 5.172126, 6.10708, 
    7.005608, 7.819336, 8.666759, 9.58604, 10.57008, 11.5552, 6.262388,
  3.126121, 3.1322, 3.138391, 3.130156, 3.110858, 3.103572, 3.123734, 
    3.158461, 3.179494, 3.181648, 3.178989, 3.18261, 3.200774, 3.23382, 
    3.258514, 3.267586, 3.288203, 3.331981, 3.377573, 3.398242, 3.394874, 
    3.388419, 3.385927, 3.396651, 3.436044, 3.499688, 3.530614, 3.536006, 
    3.540879, 3.550076, 3.565858, 3.600863, 3.663946, 3.738526, 3.7922, 
    3.808162, 3.801541, 3.802463, 3.823347, 3.859595, 3.911442, 3.993001, 
    4.09468, 4.178205, 4.272563, 4.47812, 4.936252, 5.649167, 6.541279, 
    7.40884, 8.261685, 9.159742, 10.10715, 11.14124, 12.1708, 6.262388,
  3.562569, 3.569246, 3.576355, 3.566655, 3.544049, 3.536062, 3.56063, 
    3.602159, 3.627555, 3.630917, 3.629089, 3.634759, 3.657525, 3.697295, 
    3.727661, 3.74019, 3.766024, 3.819041, 3.874451, 3.900846, 3.899343, 
    3.894371, 3.893909, 3.909257, 3.958758, 4.018147, 4.049705, 4.060171, 
    4.070033, 4.083913, 4.103719, 4.139878, 4.199914, 4.269825, 4.322034, 
    4.342344, 4.343531, 4.350992, 4.374842, 4.411198, 4.461064, 4.535445, 
    4.633432, 4.730927, 4.8405, 5.076531, 5.513181, 6.191139, 7.014067, 
    7.845285, 8.702718, 9.659621, 10.67775, 11.85297, 13.02817, 6.262388,
  4.027123, 4.033711, 4.041274, 4.035579, 4.019259, 4.015606, 4.039427, 
    4.07719, 4.102001, 4.108986, 4.111921, 4.121291, 4.14502, 4.182581, 
    4.21256, 4.227995, 4.258964, 4.322866, 4.388987, 4.420619, 4.420075, 
    4.415983, 4.417109, 4.436648, 4.495021, 4.563887, 4.601803, 4.616709, 
    4.63076, 4.649804, 4.675944, 4.720334, 4.79148, 4.873896, 4.936677, 
    4.964327, 4.970985, 4.984294, 5.01539, 5.059981, 5.120401, 5.207781, 
    5.313198, 5.399776, 5.495379, 5.694421, 6.124011, 6.731798, 7.531305, 
    8.416372, 9.354096, 10.40166, 11.52365, 12.78363, 13.85906, 6.262388,
  4.739353, 4.736605, 4.735537, 4.717043, 4.685232, 4.671457, 4.694231, 
    4.73434, 4.757846, 4.759343, 4.756516, 4.762458, 4.786486, 4.826399, 
    4.857512, 4.871931, 4.89887, 4.951952, 5.00715, 5.034749, 5.036915, 
    5.036772, 5.040344, 5.059937, 5.112045, 5.172077, 5.208554, 5.227889, 
    5.24612, 5.269487, 5.299685, 5.344851, 5.412172, 5.489141, 5.559755, 
    5.593998, 5.606876, 5.626409, 5.663593, 5.713832, 5.780399, 5.872961, 
    5.982463, 6.071897, 6.169232, 6.367417, 6.729352, 7.343995, 8.150097, 
    9.077673, 10.08037, 11.26898, 12.48716, 13.70742, 14.36202, 6.262388,
  5.667004, 5.648048, 5.630979, 5.585142, 5.519178, 5.482226, 5.502441, 
    5.549001, 5.569059, 5.555459, 5.536108, 5.53047, 5.551526, 5.594333, 
    5.624116, 5.630534, 5.653851, 5.711584, 5.770334, 5.792088, 5.781503, 
    5.769093, 5.760761, 5.773625, 5.826154, 5.8849, 5.917396, 5.932507, 
    5.945121, 5.96513, 5.994189, 6.039954, 6.109622, 6.189754, 6.25152, 
    6.284977, 6.302438, 6.325738, 6.362973, 6.410502, 6.471117, 6.552001, 
    6.645985, 6.723053, 6.824236, 7.029146, 7.397553, 7.989971, 8.82563, 
    9.806149, 10.96105, 12.38177, 13.59848, 14.31802, 14.66194, 6.262388,
  6.845986, 6.803929, 6.76335, 6.675097, 6.568592, 6.516914, 6.510757, 
    6.5533, 6.568557, 6.528468, 6.479133, 6.451841, 6.467539, 6.518003, 
    6.547027, 6.538234, 6.556142, 6.627532, 6.698659, 6.71094, 6.672799, 
    6.632189, 6.597595, 6.595252, 6.650338, 6.710574, 6.733641, 6.734084, 
    6.729829, 6.736887, 6.757089, 6.799382, 6.871575, 6.956177, 7.014411, 
    7.039359, 7.047072, 7.06441, 7.098553, 7.14487, 7.20177, 7.280066, 
    7.371525, 7.446836, 7.52686, 7.686341, 8.120902, 8.704581, 9.687585, 
    10.85786, 12.29615, 13.62948, 14.2852, 14.58595, 14.67079, 6.262388,
  8.706301, 8.635489, 8.565108, 8.457414, 8.328096, 8.232606, 8.206278, 
    8.215012, 8.190536, 8.123736, 8.051371, 7.996735, 7.975914, 7.979342, 
    7.96653, 7.924903, 7.902414, 7.919426, 7.934671, 7.905461, 7.837214, 
    7.766757, 7.697747, 7.65774, 7.66607, 7.714983, 7.721814, 7.694377, 
    7.659461, 7.641904, 7.64438, 7.680269, 7.760215, 7.857244, 7.913093, 
    7.920137, 7.90266, 7.901667, 7.925738, 7.967508, 8.017627, 8.095624, 
    8.189545, 8.267129, 8.351562, 8.534279, 8.941413, 9.656019, 10.8068, 
    12.26938, 13.70427, 14.38447, 14.61645, 14.60329, 14.67673, 6.262388,
  10.9433, 10.85271, 10.76232, 10.62292, 10.45532, 10.32845, 10.29111, 
    10.30368, 10.26944, 10.17415, 10.07123, 9.990081, 9.954312, 9.952505, 
    9.925642, 9.854568, 9.810038, 9.820988, 9.826689, 9.764466, 9.638773, 
    9.504656, 9.374514, 9.284109, 9.262474, 9.242562, 9.187706, 9.114756, 
    9.034769, 8.974702, 8.936585, 8.924655, 8.950351, 9.017918, 9.064445, 
    9.042062, 8.983212, 8.94769, 8.948771, 8.975309, 9.009264, 9.08214, 
    9.175738, 9.250498, 9.335622, 9.54838, 9.914434, 10.85448, 12.30261, 
    13.78666, 14.49002, 14.75512, 14.63902, 14.6112, 14.67805, 6.262388,
  13.26865, 13.1666, 13.06667, 12.91838, 12.74303, 12.60824, 12.56608, 
    12.58016, 12.54424, 12.44146, 12.33167, 12.2438, 12.2051, 12.20252, 
    12.17081, 12.08671, 12.03158, 12.03824, 12.03587, 11.95175, 11.78202, 
    11.59321, 11.40829, 11.26856, 11.21216, 11.15994, 11.06182, 10.9384, 
    10.81144, 10.71233, 10.64398, 10.60174, 10.6093, 10.63913, 10.63428, 
    10.57319, 10.4802, 10.4001, 10.34645, 10.31088, 10.27961, 10.33857, 
    10.43493, 10.50192, 10.58408, 10.83973, 11.29889, 12.49903, 13.8954, 
    14.62064, 14.78893, 14.77866, 14.6484, 14.61281, 14.6791, 6.262388,
  15.5616, 15.45212, 15.34839, 15.20205, 15.03238, 14.90344, 14.86545, 
    14.88464, 14.85534, 14.76074, 14.66308, 14.58744, 14.56122, 14.56497, 
    14.54067, 14.46437, 14.41311, 14.42144, 14.41804, 14.32889, 14.13981, 
    13.92034, 13.70124, 13.52678, 13.44186, 13.36147, 13.22938, 13.06699, 
    12.90467, 12.77928, 12.69467, 12.63091, 12.63068, 12.66143, 12.66652, 
    12.59613, 12.47896, 12.35671, 12.25768, 12.17105, 12.11829, 12.12187, 
    12.21153, 12.24886, 12.30803, 12.59807, 13.22473, 14.19771, 14.759, 
    14.85799, 14.79715, 14.78855, 14.65008, 14.61447, 14.68149, 6.262388,
  17.45164, 17.33763, 17.24136, 17.1328, 17.01126, 16.92144, 16.89837, 
    16.91749, 16.90403, 16.84352, 16.78717, 16.74694, 16.74432, 16.75379, 
    16.74323, 16.69303, 16.6559, 16.66158, 16.65525, 16.58029, 16.4161, 
    16.21827, 16.01841, 15.85181, 15.76322, 15.67975, 15.5467, 15.37984, 
    15.21722, 15.09352, 15.01311, 14.94371, 14.94608, 14.987, 15.01583, 
    14.96161, 14.85395, 14.72474, 14.61043, 14.50051, 14.45652, 14.43091, 
    14.41957, 14.34906, 14.30234, 14.44751, 14.90435, 14.9102, 14.96158, 
    14.85825, 14.8004, 14.78997, 14.65201, 14.61668, 14.68353, 6.262388,
  18.12847, 18.01842, 17.93835, 17.88674, 17.84173, 17.81504, 17.81018, 
    17.8139, 17.81645, 17.8148, 17.81823, 17.81829, 17.81849, 17.81686, 
    17.79679, 17.75339, 17.72352, 17.67727, 17.60417, 17.53641, 17.44536, 
    17.34006, 17.218, 17.1126, 17.04256, 16.97945, 16.90094, 16.80568, 
    16.72929, 16.67172, 16.636, 16.57844, 16.55952, 16.53228, 16.50419, 
    16.4524, 16.37827, 16.27213, 16.14913, 16.00877, 15.89535, 15.77133, 
    15.6351, 15.46906, 15.32083, 15.20582, 15.09438, 15.00554, 14.96251, 
    14.8584, 14.80099, 14.79222, 14.65429, 14.61843, 14.68517, 6.262388,
  18.13201, 18.02542, 17.95132, 17.9098, 17.87545, 17.86155, 17.86823, 
    17.87956, 17.89414, 17.91168, 17.92946, 17.93475, 17.92764, 17.92982, 
    17.90746, 17.86054, 17.83078, 17.76926, 17.67592, 17.60426, 17.52691, 
    17.44368, 17.33463, 17.2434, 17.16995, 17.08702, 17.01142, 16.9427, 
    16.89274, 16.85521, 16.83031, 16.76007, 16.69197, 16.62289, 16.59185, 
    16.53831, 16.4627, 16.35743, 16.23236, 16.08739, 15.97196, 15.84036, 
    15.69253, 15.53766, 15.39806, 15.27358, 15.10898, 15.00527, 14.96261, 
    14.85848, 14.80485, 14.79493, 14.65612, 14.61985, 14.68621, 6.262388,
  18.12733, 18.02046, 17.94744, 17.90826, 17.8772, 17.86592, 17.87464, 
    17.88956, 17.90705, 17.92694, 17.94617, 17.95103, 17.94163, 17.94267, 
    17.91852, 17.86916, 17.83633, 17.77234, 17.67705, 17.60527, 17.52744, 
    17.44362, 17.33255, 17.23961, 17.16467, 17.08205, 17.01192, 16.95426, 
    16.90949, 16.87496, 16.8507, 16.78439, 16.71602, 16.64528, 16.61064, 
    16.55471, 16.47774, 16.36185, 16.23105, 16.08527, 15.97025, 15.83871, 
    15.69061, 15.53555, 15.39593, 15.27161, 15.10774, 15.00459, 14.96578, 
    14.86565, 14.80918, 14.79713, 14.65724, 14.6201, 14.68621, 6.262388,
  18.13222, 18.02454, 17.95127, 17.91236, 17.88393, 17.87457, 17.88442, 
    17.90185, 17.92061, 17.94062, 17.96073, 17.96693, 17.95931, 17.95914, 
    17.93371, 17.88297, 17.85378, 17.79075, 17.6935, 17.62229, 17.5445, 
    17.46034, 17.34999, 17.25754, 17.18319, 17.10089, 17.03044, 16.97192, 
    16.92716, 16.89421, 16.87309, 16.80853, 16.74173, 16.6726, 16.63876, 
    16.58343, 16.50673, 16.38755, 16.25198, 16.09988, 15.97467, 15.83854, 
    15.69115, 15.53661, 15.39749, 15.27486, 15.11418, 15.01483, 14.97561, 
    14.87177, 14.8118, 14.79764, 14.65724, 14.6201, 14.68621, 6.262388,
  18.14363, 18.03578, 17.96225, 17.92302, 17.89565, 17.8868, 17.89651, 
    17.91446, 17.93315, 17.95256, 17.97298, 17.97948, 17.97208, 17.97134, 
    17.94492, 17.89278, 17.86407, 17.80091, 17.7033, 17.63271, 17.55551, 
    17.47173, 17.36205, 17.27086, 17.19822, 17.11613, 17.04762, 16.99273, 
    16.95018, 16.91881, 16.89862, 16.83256, 16.76501, 16.69596, 16.66158, 
    16.60649, 16.53068, 16.41279, 16.27823, 16.127, 16.00248, 15.86557, 
    15.71629, 15.55689, 15.41522, 15.29129, 15.12689, 15.02287, 14.97923, 
    14.87233, 14.8118, 14.79764, 14.65724, 14.6201, 14.68621, 6.262388 ;

 temp_north =
  1.245957, 1.24621, 1.267426, 1.304018, 1.338612, 1.357394, 1.372541, 
    1.397368, 1.41785, 1.430443, 1.446943, 1.465768, 1.483243, 1.503218, 
    1.522053, 1.529888, 1.524523, 1.514423, 1.511968, 1.528278, 1.612276, 
    1.826295, 2.329157, 3.138641, 4.067322, 5.069591, 5.968559, 6.746574, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  1.310103, 1.310213, 1.329811, 1.374272, 1.428578, 1.45329, 1.467158, 
    1.489659, 1.508684, 1.521006, 1.536775, 1.565065, 1.591098, 1.62052, 
    1.647983, 1.659136, 1.650975, 1.635939, 1.632116, 1.655813, 1.742854, 
    2.009727, 2.558835, 3.372389, 4.294739, 5.256949, 6.13126, 6.880507, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  1.377501, 1.377518, 1.409097, 1.463014, 1.512623, 1.537435, 1.559012, 
    1.594257, 1.62365, 1.641751, 1.664916, 1.690865, 1.714546, 1.741395, 
    1.766508, 1.776754, 1.769624, 1.756016, 1.752481, 1.77442, 1.864749, 
    2.176995, 2.755141, 3.572209, 4.489198, 5.437089, 6.270554, 6.995317, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  1.460587, 1.460584, 1.489643, 1.544857, 1.622458, 1.657959, 1.677989, 
    1.710521, 1.737544, 1.754053, 1.77523, 1.798974, 1.820634, 1.85375, 
    1.893084, 1.909121, 1.897205, 1.875021, 1.869172, 1.904536, 2.033986, 
    2.325309, 2.923874, 3.761423, 4.690339, 5.598116, 6.390507, 7.186949, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  1.534149, 1.534139, 1.579539, 1.657368, 1.729393, 1.762435, 1.781124, 
    1.811304, 1.841269, 1.8658, 1.898082, 1.934951, 1.969192, 2.008378, 
    2.045478, 2.061001, 2.051019, 2.031293, 2.026429, 2.060542, 2.180697, 
    2.51515, 3.122961, 3.97482, 4.87116, 5.737887, 6.500329, 7.36262, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  1.640938, 1.641171, 1.683602, 1.756175, 1.823305, 1.871377, 1.899736, 
    1.946168, 1.98476, 2.00835, 2.039188, 2.07433, 2.107075, 2.144179, 
    2.179319, 2.194391, 2.186108, 2.16854, 2.164541, 2.197555, 2.309551, 
    2.681892, 3.307418, 4.162317, 5.03009, 5.860807, 6.6256, 7.517515, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  1.736491, 1.736943, 1.776718, 1.856634, 1.958109, 2.005298, 2.032446, 
    2.07645, 2.113161, 2.13591, 2.165456, 2.199053, 2.23046, 2.265703, 
    2.302195, 2.322878, 2.310505, 2.291356, 2.288132, 2.325265, 2.481927, 
    2.831116, 3.472515, 4.330171, 5.172417, 5.980026, 6.737951, 7.656651, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  1.825388, 1.826054, 1.885706, 1.987958, 2.083417, 2.128201, 2.154239, 
    2.196015, 2.231, 2.252976, 2.281904, 2.328182, 2.37163, 2.420518, 
    2.466939, 2.48728, 2.477153, 2.455009, 2.45067, 2.494319, 2.641438, 
    2.978266, 3.62406, 4.484274, 5.310036, 6.101804, 6.841259, 7.897038, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  1.958394, 1.959854, 2.016243, 2.112302, 2.202066, 2.244572, 2.270417, 
    2.327812, 2.375901, 2.405959, 2.445134, 2.489796, 2.531869, 2.578575, 
    2.622933, 2.64295, 2.634949, 2.615603, 2.612685, 2.654394, 2.792478, 
    3.163711, 3.798753, 4.655183, 5.456071, 6.2172, 6.939206, 8.169513, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  2.088728, 2.090967, 2.144159, 2.234148, 2.344714, 2.40263, 2.436994, 
    2.491786, 2.537869, 2.567149, 2.605088, 2.648166, 2.688891, 2.733459, 
    2.775796, 2.795495, 2.789578, 2.772973, 2.771448, 2.811256, 2.940488, 
    3.345437, 4.000491, 4.830882, 5.599199, 6.330312, 7.076134, 8.436745, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  2.220614, 2.223639, 2.282341, 2.403226, 2.517056, 2.572176, 2.605552, 
    2.657709, 2.701763, 2.730256, 2.766943, 2.808419, 2.847781, 2.890186, 
    2.942712, 2.967615, 2.958703, 2.936357, 2.933973, 2.984316, 3.152753, 
    3.529321, 4.204621, 5.00866, 5.744015, 6.44475, 7.257391, 8.70702, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  2.406135, 2.410783, 2.477599, 2.589825, 2.695608, 2.74783, 2.780183, 
    2.829611, 2.877982, 2.914063, 2.960737, 3.0135, 3.0634, 3.117434, 
    3.168739, 3.193139, 3.18709, 3.168755, 3.168573, 3.216375, 3.372772, 
    3.735641, 4.416087, 5.192811, 5.894259, 6.603612, 7.445015, 8.985534, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  2.612982, 2.619536, 2.681922, 2.785084, 2.905399, 2.971439, 3.012515, 
    3.075431, 3.128769, 3.16384, 3.208602, 3.258782, 3.306335, 3.357081, 
    3.405249, 3.429123, 3.42607, 3.411933, 3.414054, 3.459198, 3.602993, 
    4.020767, 4.665866, 5.406788, 6.087566, 6.773714, 7.653823, 9.276009, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  2.842401, 2.851133, 2.928805, 3.05707, 3.178497, 3.240421, 3.280207, 
    3.339285, 3.389665, 3.423684, 3.466458, 3.513949, 3.559061, 3.612216, 
    3.670419, 3.699097, 3.694571, 3.676779, 3.679224, 3.734251, 3.914425, 
    4.317374, 4.947594, 5.641399, 6.288604, 6.95058, 8.189198, 9.57774, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  3.148876, 3.160818, 3.232316, 3.347522, 3.456789, 3.524746, 3.572603, 
    3.64359, 3.704033, 3.744807, 3.795814, 3.852399, 3.906152, 3.962761, 
    4.01661, 4.044854, 4.045604, 4.034829, 4.041473, 4.0949, 4.2595, 
    4.650807, 5.234666, 5.880734, 6.514492, 7.241356, 8.734527, 9.747207, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  3.465548, 3.480754, 3.565494, 3.701151, 3.829767, 3.898143, 3.943992, 
    4.009625, 4.06598, 4.10535, 4.153403, 4.2062, 4.256636, 4.308633, 
    4.364947, 4.396713, 4.398715, 4.388611, 4.398893, 4.457904, 4.636822, 
    5.018706, 5.565107, 6.170244, 6.78921, 7.54401, 9.230739, 9.90495, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  3.862947, 3.881897, 3.958332, 4.076886, 4.20312, 4.28111, 4.333273, 
    4.407238, 4.470118, 4.513614, 4.566523, 4.624382, 4.679407, 4.735268, 
    4.787935, 4.816738, 4.822724, 4.818359, 4.829559, 4.883456, 5.039683, 
    5.395751, 5.885077, 6.45725, 7.098429, 8.312657, 9.657565, 9.969707, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  4.287123, 4.309016, 4.395475, 4.528418, 4.652891, 4.721354, 4.769054, 
    4.834115, 4.889766, 4.929307, 4.979548, 5.041674, 5.099886, 5.156789, 
    5.20893, 5.235512, 5.240201, 5.234764, 5.244898, 5.29633, 5.449494, 
    5.772014, 6.239637, 6.797163, 7.465186, 9.033981, 9.785495, 9.962668, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  4.730273, 4.754196, 4.847495, 5.002749, 5.143881, 5.217457, 5.266278, 
    5.332232, 5.385851, 5.420258, 5.465323, 5.514446, 5.560974, 5.601872, 
    5.638994, 5.655868, 5.659083, 5.65366, 5.659953, 5.699368, 5.841367, 
    6.1702, 6.606461, 7.201584, 8.309376, 9.605104, 9.858678, 9.956853, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  5.297616, 5.319724, 5.401657, 5.524809, 5.671625, 5.751658, 5.800555, 
    5.86771, 5.918239, 5.944163, 5.984531, 6.028951, 6.069735, 6.098689, 
    6.12224, 6.123118, 6.113697, 6.095208, 6.088432, 6.116451, 6.242064, 
    6.570706, 6.996988, 7.762683, 9.085742, 9.66643, 9.852953, 9.95568, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  5.933947, 5.953869, 6.045378, 6.184854, 6.305823, 6.360886, 6.393981, 
    6.45084, 6.489282, 6.500584, 6.530526, 6.565409, 6.597153, 6.611278, 
    6.61827, 6.599247, 6.575433, 6.540245, 6.515649, 6.532207, 6.660822, 
    6.991693, 7.481159, 8.570871, 9.475721, 9.689924, 9.848933, 9.954707, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  6.601238, 6.620006, 6.708712, 6.844537, 6.96105, 7.009423, 7.030231, 
    7.062696, 7.077682, 7.0717, 7.097851, 7.131819, 7.163863, 7.174197, 
    7.171784, 7.130533, 7.087871, 7.027197, 6.97697, 6.987247, 7.138068, 
    7.496853, 8.273354, 9.282553, 9.466999, 9.686647, 9.847492, 9.954126, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  7.280087, 7.298243, 7.39325, 7.540055, 7.665428, 7.714491, 7.732381, 
    7.769241, 7.787574, 7.779332, 7.79004, 7.828151, 7.874927, 7.896694, 
    7.891066, 7.820716, 7.749943, 7.65168, 7.564209, 7.573371, 7.780179, 
    8.314257, 9.049097, 9.314894, 9.466215, 9.684662, 9.846343, 9.953871, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  8.053718, 8.069534, 8.174252, 8.342855, 8.498165, 8.565199, 8.593062, 
    8.662016, 8.712484, 8.732795, 8.760833, 8.782416, 8.793197, 8.785297, 
    8.738009, 8.628796, 8.542135, 8.431669, 8.324265, 8.33378, 8.561695, 
    9.094908, 9.198695, 9.322967, 9.465496, 9.683416, 9.845759, 9.953666, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  8.775131, 8.802241, 8.847577, 8.914437, 8.986495, 9.035107, 9.071488, 
    9.134012, 9.192887, 9.242589, 9.273397, 9.271971, 9.247445, 9.225661, 
    9.159841, 9.050269, 8.981463, 8.91772, 8.857529, 8.882457, 8.975542, 
    9.136733, 9.213281, 9.32319, 9.464646, 9.682498, 9.845327, 9.9535, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  8.885454, 8.932167, 8.979181, 9.026379, 9.069717, 9.107424, 9.139755, 
    9.183731, 9.224627, 9.262288, 9.282115, 9.275706, 9.242622, 9.221846, 
    9.159096, 9.054259, 8.968754, 8.890588, 8.819575, 8.87495, 8.980664, 
    9.136898, 9.213085, 9.322563, 9.463881, 9.681834, 9.844982, 9.953402, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  8.890863, 8.936971, 8.983357, 9.030029, 9.072984, 9.110579, 9.142873, 
    9.186733, 9.227396, 9.264832, 9.284437, 9.277658, 9.244469, 9.2239, 
    9.160919, 9.05545, 8.967244, 8.887074, 8.814813, 8.870517, 8.977069, 
    9.135388, 9.212781, 9.321939, 9.463029, 9.681302, 9.844759, 9.953402, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  8.893392, 8.9387, 8.984726, 9.031461, 9.074368, 9.111878, 9.144028, 
    9.18796, 9.228607, 9.265952, 9.28569, 9.278975, 9.245792, 9.225298, 
    9.162257, 9.05664, 8.967952, 8.887297, 8.814701, 8.870156, 8.977078, 
    9.135494, 9.212236, 9.321132, 9.462341, 9.680987, 9.844759, 9.953402, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  8.894401, 8.939698, 8.985659, 9.03229, 9.075052, 9.112443, 9.14445, 
    9.188402, 9.228995, 9.266229, 9.285987, 9.279239, 9.245988, 9.22549, 
    9.162396, 9.056715, 8.96814, 8.887542, 8.814918, 8.870014, 8.976653, 
    9.134772, 9.211488, 9.320496, 9.462088, 9.680987, 9.844759, 9.953402, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  8.894047, 8.939241, 8.985186, 9.031881, 9.074703, 9.112122, 9.144136, 
    9.188128, 9.228708, 9.265879, 9.285584, 9.278778, 9.245461, 9.22501, 
    9.161934, 9.056231, 8.967778, 8.887237, 8.814606, 8.869612, 8.976202, 
    9.134377, 9.211259, 9.320496, 9.462088, 9.680987, 9.844759, 9.953402, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 
    6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131, 6.362131,
  1.2455, 1.245733, 1.266942, 1.303443, 1.33789, 1.356524, 1.371479, 
    1.396243, 1.416652, 1.429175, 1.445899, 1.46496, 1.48269, 1.502868, 
    1.521868, 1.529759, 1.524101, 1.513778, 1.511183, 1.527096, 1.61017, 
    1.823348, 2.326532, 3.145936, 4.08553, 5.100328, 6.021739, 6.852392, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  1.309547, 1.309707, 1.329278, 1.373518, 1.427586, 1.452053, 1.465614, 
    1.488099, 1.507111, 1.519439, 1.535604, 1.564232, 1.590597, 1.6202, 
    1.647761, 1.658929, 1.650082, 1.634692, 1.630673, 1.653107, 1.738968, 
    2.006618, 2.559304, 3.382565, 4.316866, 5.292053, 6.189271, 7.006361, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  1.376846, 1.376954, 1.40844, 1.462026, 1.511379, 1.53588, 1.557044, 
    1.592281, 1.621671, 1.639798, 1.663376, 1.689728, 1.713831, 1.740911, 
    1.766147, 1.776407, 1.76814, 1.753905, 1.750094, 1.770091, 1.859436, 
    2.173849, 2.758254, 3.584847, 4.514678, 5.477215, 6.3327, 7.138349, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  1.459817, 1.459904, 1.488839, 1.54365, 1.620889, 1.656024, 1.675608, 
    1.708143, 1.735183, 1.751743, 1.773371, 1.797576, 1.819735, 1.853125, 
    1.892644, 1.908769, 1.89544, 1.872357, 1.866147, 1.8991, 2.028026, 
    2.322327, 2.92926, 3.776638, 4.719925, 5.642956, 6.456213, 7.367796, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  1.533274, 1.533352, 1.578541, 1.655846, 1.72751, 1.76017, 1.778386, 
    1.808578, 1.838575, 1.863192, 1.895966, 1.93333, 1.968062, 2.007632, 
    2.045042, 2.060781, 2.049392, 2.028784, 2.023585, 2.054578, 2.174177, 
    2.514892, 3.131134, 3.993565, 4.90454, 5.786819, 6.571452, 7.578598, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  1.639819, 1.640143, 1.682352, 1.754376, 1.821146, 1.868784, 1.896662, 
    1.943118, 1.981785, 2.005517, 2.036876, 2.072517, 2.105733, 2.143329, 
    2.178888, 2.194288, 2.184601, 2.166166, 2.161856, 2.191128, 2.302538, 
    2.684028, 3.318184, 4.184164, 5.066804, 5.913338, 6.713408, 7.764469, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  1.735154, 1.735699, 1.775242, 1.854548, 1.955555, 2.002336, 2.029053, 
    2.073109, 2.109935, 2.132875, 2.162968, 2.197068, 2.228928, 2.264759, 
    2.30177, 2.322922, 2.309153, 2.289104, 2.285589, 2.318658, 2.477391, 
    2.835394, 3.485602, 4.354794, 5.212117, 6.035927, 6.840723, 7.93143, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  1.823844, 1.824606, 1.883933, 1.985492, 2.080497, 2.124899, 2.150553, 
    2.192406, 2.227543, 2.249757, 2.279249, 2.325992, 2.36988, 2.419464, 
    2.46661, 2.487696, 2.476624, 2.453852, 2.449433, 2.489878, 2.63924, 
    2.984723, 3.639278, 4.511446, 5.352926, 6.161009, 6.95779, 8.151769, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  1.95647, 1.958018, 2.014091, 2.109476, 2.198799, 2.24095, 2.26645, 
    2.323891, 2.372112, 2.402423, 2.442135, 2.487299, 2.529876, 2.577414, 
    2.622694, 2.643716, 2.635198, 2.615588, 2.612875, 2.652004, 2.792492, 
    3.173172, 3.816633, 4.685387, 5.503007, 6.279536, 7.068783, 8.387207, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  2.086432, 2.08875, 2.141633, 2.23097, 2.341042, 2.398584, 2.432616, 
    2.487455, 2.533693, 2.563267, 2.60175, 2.645368, 2.686661, 2.732193, 
    2.775646, 2.796606, 2.790591, 2.774078, 2.773037, 2.810875, 2.942671, 
    3.357842, 4.021594, 4.864256, 5.650101, 6.395718, 7.232646, 8.618114, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  2.217941, 2.221037, 2.279411, 2.399576, 2.512909, 2.567679, 2.60076, 
    2.652964, 2.697195, 2.726024, 2.763264, 2.805316, 2.84531, 2.888813, 
    2.942698, 2.969236, 2.960728, 2.938708, 2.937041, 2.986638, 3.159759, 
    3.544706, 4.228987, 5.045242, 5.798929, 6.513262, 7.456049, 8.851652, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  2.402938, 2.407643, 2.474117, 2.58566, 2.690969, 2.742867, 2.774961, 
    2.824436, 2.872961, 2.909364, 2.956511, 3.009865, 3.060595, 3.115976, 
    3.169084, 3.195725, 3.191168, 3.174069, 3.175293, 3.223932, 3.384772, 
    3.754342, 4.443832, 5.232717, 5.953322, 6.689865, 7.687301, 9.008857, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  2.609205, 2.615802, 2.677861, 2.780381, 2.900139, 2.965792, 3.006558, 
    3.069392, 3.122842, 3.158272, 3.203489, 3.254429, 3.303159, 3.355539, 
    3.405971, 3.43272, 3.432297, 3.420347, 3.424597, 3.472231, 3.620218, 
    4.043904, 4.697464, 5.451077, 6.151078, 6.879975, 7.936086, 9.139157, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  2.837958, 2.846715, 2.923985, 3.051483, 3.172349, 3.233892, 3.273342, 
    3.332299, 3.382796, 3.417213, 3.460422, 3.508849, 3.555498, 3.610574, 
    3.671577, 3.703927, 3.703215, 3.68857, 3.693923, 3.753302, 3.938009, 
    4.345125, 4.983426, 5.690755, 6.356743, 7.077646, 8.37468, 9.274508, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  3.143456, 3.155388, 3.226492, 3.340973, 3.449736, 3.51721, 3.564603, 
    3.635251, 3.695663, 3.736794, 3.78815, 3.845928, 3.901878, 3.960926, 
    4.018413, 4.051475, 4.057413, 4.051156, 4.062014, 4.121174, 4.289903, 
    4.68316, 5.274814, 5.935258, 6.594157, 7.444654, 8.821426, 9.281816, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  3.459034, 3.474185, 3.558341, 3.692973, 3.820843, 3.888692, 3.934019, 
    3.999243, 4.055565, 4.095347, 4.14381, 4.198231, 4.251642, 4.306607, 
    4.367339, 4.405052, 4.413615, 4.409416, 4.425198, 4.491298, 4.673801, 
    5.055458, 5.610755, 6.23001, 6.897085, 7.830447, 9.037585, 9.279936, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  3.854541, 3.873326, 3.949164, 4.06676, 4.192363, 4.26983, 4.321373, 
    4.394754, 4.457452, 4.501256, 4.554517, 4.614347, 4.673112, 4.73236, 
    4.790318, 4.826348, 4.840105, 4.843112, 4.861496, 4.923382, 5.082692, 
    5.437228, 5.935996, 6.527196, 7.269145, 8.469343, 9.176283, 9.26673, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  4.277235, 4.298769, 4.384559, 4.516523, 4.640506, 4.708406, 4.755311, 
    4.819527, 4.874803, 4.914507, 4.965041, 5.029413, 5.092142, 5.152842, 
    5.211209, 5.246536, 5.260462, 5.263991, 5.283147, 5.343765, 5.500137, 
    5.818426, 6.295386, 6.909492, 7.756647, 8.922326, 9.15218, 9.245784, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  4.719381, 4.742665, 4.834918, 4.988655, 5.12948, 5.202552, 5.250181, 
    5.314982, 5.367848, 5.401946, 5.447012, 5.498933, 5.551254, 5.596487, 
    5.641043, 5.668519, 5.682921, 5.688692, 5.706445, 5.755907, 5.900147, 
    6.220753, 6.69159, 7.414134, 8.493544, 9.074056, 9.118957, 9.227711, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  5.283937, 5.305204, 5.385936, 5.507582, 5.653279, 5.73208, 5.778859, 
    5.843968, 5.892894, 5.917742, 5.957554, 6.005213, 6.053413, 6.08672, 
    6.118748, 6.132558, 6.138668, 6.135108, 6.142914, 6.183603, 6.310002, 
    6.644467, 7.145537, 8.042947, 8.885116, 9.004281, 9.069715, 9.21582, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  5.909097, 5.928159, 6.017141, 6.152972, 6.274635, 6.329611, 6.360882, 
    6.41781, 6.455679, 6.465568, 6.49519, 6.534958, 6.577274, 6.595447, 
    6.612441, 6.60986, 6.609645, 6.595407, 6.590385, 6.627825, 6.768495, 
    7.124302, 7.767109, 8.704806, 8.917662, 8.937886, 9.029695, 9.205968, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  6.571085, 6.588748, 6.677146, 6.812906, 6.936154, 6.986323, 7.003834, 
    7.035451, 7.047778, 7.037532, 7.063308, 7.103855, 7.149562, 7.162134, 
    7.172574, 7.155423, 7.147761, 7.118564, 7.098998, 7.144939, 7.334332, 
    7.76004, 8.51723, 8.890981, 8.790522, 8.876978, 8.998861, 9.198643, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  7.26522, 7.282465, 7.380837, 7.534199, 7.677644, 7.733049, 7.746973, 
    7.785235, 7.800112, 7.782821, 7.784188, 7.812715, 7.855638, 7.861645, 
    7.86367, 7.830834, 7.81505, 7.775656, 7.746192, 7.801632, 8.026665, 
    8.5189, 8.787936, 8.713651, 8.72548, 8.827675, 8.974268, 9.193447, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  8.026809, 8.045335, 8.126633, 8.254253, 8.379496, 8.432811, 8.451886, 
    8.500279, 8.532369, 8.539518, 8.549438, 8.547565, 8.540124, 8.516006, 
    8.480927, 8.426221, 8.414773, 8.396402, 8.37838, 8.424245, 8.545591, 
    8.738806, 8.663361, 8.644545, 8.672573, 8.788335, 8.955485, 9.189279, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  8.46542, 8.498246, 8.505643, 8.500601, 8.505439, 8.522048, 8.539491, 
    8.560914, 8.582428, 8.603366, 8.617355, 8.619307, 8.609044, 8.607809, 
    8.581034, 8.53019, 8.518718, 8.514446, 8.513552, 8.562596, 8.595395, 
    8.602793, 8.585411, 8.615152, 8.625932, 8.757768, 8.94064, 9.185922, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  8.29427, 8.340991, 8.385525, 8.427224, 8.467234, 8.499536, 8.524328, 
    8.556134, 8.584125, 8.608197, 8.615553, 8.60854, 8.587181, 8.58257, 
    8.554281, 8.502302, 8.464011, 8.426552, 8.389888, 8.428865, 8.486185, 
    8.554317, 8.56803, 8.595769, 8.589727, 8.733973, 8.928759, 9.183905, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  8.30487, 8.350659, 8.393442, 8.432896, 8.471384, 8.502049, 8.525118, 
    8.557068, 8.585025, 8.608995, 8.615446, 8.608089, 8.586941, 8.582458, 
    8.554212, 8.502192, 8.462961, 8.423017, 8.382333, 8.419756, 8.471973, 
    8.539445, 8.56514, 8.580795, 8.562089, 8.714919, 8.921031, 9.183905, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  8.311923, 8.355963, 8.397163, 8.435447, 8.473177, 8.503417, 8.526216, 
    8.558029, 8.585896, 8.609814, 8.616069, 8.608389, 8.586743, 8.58217, 
    8.55372, 8.501399, 8.461893, 8.421409, 8.379916, 8.417391, 8.469882, 
    8.536789, 8.563216, 8.569563, 8.539781, 8.703568, 8.921031, 9.183905, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  8.313994, 8.357833, 8.398724, 8.436629, 8.474208, 8.504337, 8.527034, 
    8.55875, 8.58656, 8.610467, 8.616557, 8.608436, 8.586082, 8.581421, 
    8.552763, 8.500118, 8.460227, 8.419559, 8.378067, 8.416103, 8.468533, 
    8.535147, 8.56203, 8.56073, 8.531516, 8.703568, 8.921031, 9.183905, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388,
  8.315222, 8.358829, 8.399449, 8.437082, 8.474545, 8.504587, 8.527208, 
    8.558853, 8.586631, 8.61054, 8.616548, 8.608116, 8.585246, 8.580614, 
    8.55187, 8.499016, 8.458711, 8.417808, 8.376307, 8.415048, 8.467724, 
    8.534336, 8.56167, 8.56073, 8.531516, 8.703568, 8.921031, 9.183905, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 
    6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388, 6.262388 ;

 salt_west =
  34.68758, 34.68752, 34.68773, 34.688, 34.68818, 34.68819, 34.68806, 
    34.68793, 34.68801, 34.68829, 34.68863, 34.68903, 34.68933, 34.68948, 
    34.68953, 34.68957, 34.6896, 34.68964, 34.68967, 34.68954, 34.68928, 
    34.68903, 34.6888, 34.68864, 34.68854, 34.68827, 34.6878, 34.68737, 
    34.68641, 34.68388, 34.68103, 34.6786, 34.67691, 34.67513, 34.67365, 
    34.67284, 34.67256, 34.67258, 34.67274, 34.67279, 34.67245, 34.6721, 
    34.67212, 34.67223, 34.67226, 34.67223, 34.67197, 34.67142, 34.67092, 
    34.6707, 34.67055, 34.66994, 34.66881, 34.66777, 34.66766,
  34.6845, 34.68444, 34.6847, 34.68489, 34.68499, 34.68494, 34.68478, 
    34.68462, 34.68465, 34.68506, 34.68584, 34.68676, 34.68747, 34.6878, 
    34.68789, 34.68787, 34.68781, 34.68777, 34.68774, 34.68756, 34.68713, 
    34.68655, 34.68605, 34.68564, 34.68535, 34.6848, 34.68392, 34.68315, 
    34.68194, 34.67876, 34.67508, 34.6729, 34.67097, 34.66873, 34.6669, 
    34.66589, 34.66558, 34.66574, 34.66611, 34.66626, 34.66578, 34.66529, 
    34.66541, 34.66569, 34.66582, 34.66586, 34.66549, 34.66462, 34.66386, 
    34.66357, 34.66336, 34.6625, 34.66089, 34.65948, 34.65937,
  34.67997, 34.6799, 34.68021, 34.68055, 34.68074, 34.68069, 34.68046, 
    34.68024, 34.68033, 34.68097, 34.68216, 34.68352, 34.68419, 34.68445, 
    34.6845, 34.68449, 34.68442, 34.68439, 34.68434, 34.68399, 34.68339, 
    34.6828, 34.68229, 34.68176, 34.68132, 34.68055, 34.67933, 34.67826, 
    34.67664, 34.67345, 34.66885, 34.66602, 34.66404, 34.66194, 34.66023, 
    34.65921, 34.65881, 34.659, 34.65928, 34.65934, 34.65881, 34.65828, 
    34.6583, 34.65848, 34.65852, 34.6585, 34.65808, 34.65724, 34.65651, 
    34.65622, 34.656, 34.65519, 34.65291, 34.65061, 34.65049,
  34.6751, 34.67502, 34.67548, 34.676, 34.6763, 34.67626, 34.67596, 34.67568, 
    34.67583, 34.67675, 34.67786, 34.6791, 34.68003, 34.68044, 34.68052, 
    34.68053, 34.68047, 34.68043, 34.68037, 34.6799, 34.67907, 34.67825, 
    34.67754, 34.67693, 34.67646, 34.67569, 34.6745, 34.67341, 34.67128, 
    34.66708, 34.66262, 34.65947, 34.6563, 34.65289, 34.6501, 34.64854, 
    34.64806, 34.64833, 34.64897, 34.64923, 34.64852, 34.64779, 34.648, 
    34.64847, 34.64869, 34.64878, 34.64825, 34.64698, 34.64588, 34.64553, 
    34.64529, 34.644, 34.64157, 34.63943, 34.63929,
  34.66994, 34.66985, 34.67025, 34.67072, 34.67096, 34.67089, 34.67059, 
    34.67031, 34.67042, 34.67125, 34.67279, 34.67456, 34.67589, 34.67645, 
    34.67649, 34.67646, 34.67636, 34.67628, 34.67618, 34.6757, 34.67487, 
    34.67377, 34.67281, 34.672, 34.67137, 34.67036, 34.66877, 34.66735, 
    34.66531, 34.66138, 34.65427, 34.64987, 34.64681, 34.64354, 34.64084, 
    34.63929, 34.63874, 34.63889, 34.63937, 34.63952, 34.63874, 34.63797, 
    34.63809, 34.63844, 34.63858, 34.63863, 34.63809, 34.63687, 34.63582, 
    34.63547, 34.63522, 34.63401, 34.63174, 34.62946, 34.62931,
  34.66393, 34.66383, 34.66452, 34.6653, 34.66576, 34.66573, 34.6653, 
    34.66492, 34.66517, 34.66642, 34.66783, 34.66945, 34.67068, 34.6712, 
    34.67131, 34.67133, 34.67125, 34.6712, 34.6711, 34.67049, 34.66941, 
    34.66835, 34.6674, 34.66659, 34.66594, 34.66494, 34.6634, 34.66203, 
    34.65899, 34.65253, 34.64563, 34.64144, 34.63848, 34.63324, 34.62866, 
    34.62613, 34.6254, 34.62593, 34.62707, 34.62762, 34.62657, 34.62551, 
    34.626, 34.6269, 34.62738, 34.62767, 34.62693, 34.62498, 34.62331, 
    34.62286, 34.62256, 34.62052, 34.61658, 34.61311, 34.61296,
  34.65708, 34.65696, 34.65756, 34.65826, 34.65863, 34.65856, 34.65811, 
    34.65771, 34.65789, 34.65914, 34.66146, 34.66412, 34.66601, 34.66647, 
    34.66655, 34.66652, 34.66641, 34.66633, 34.66619, 34.66558, 34.66453, 
    34.66344, 34.66199, 34.66078, 34.65985, 34.65832, 34.6559, 34.65371, 
    34.65057, 34.64444, 34.63675, 34.62943, 34.62437, 34.619, 34.61458, 
    34.61208, 34.61125, 34.6116, 34.61253, 34.61291, 34.61178, 34.61066, 
    34.61102, 34.61175, 34.61212, 34.61233, 34.61158, 34.60971, 34.60812, 
    34.60765, 34.60735, 34.60543, 34.60174, 34.59849, 34.59832,
  34.65079, 34.65065, 34.65118, 34.65179, 34.6521, 34.65197, 34.65151, 
    34.65109, 34.65122, 34.65234, 34.65446, 34.6569, 34.65876, 34.65958, 
    34.65979, 34.65985, 34.65981, 34.65979, 34.65968, 34.6588, 34.65718, 
    34.65556, 34.65412, 34.6529, 34.65193, 34.65039, 34.64803, 34.64589, 
    34.64284, 34.63452, 34.62296, 34.61598, 34.61111, 34.60593, 34.60166, 
    34.59918, 34.59826, 34.59845, 34.59919, 34.59941, 34.59821, 34.59704, 
    34.59728, 34.59785, 34.59811, 34.59825, 34.59749, 34.5957, 34.59418, 
    34.5937, 34.59339, 34.59159, 34.58812, 34.58481, 34.58464,
  34.64055, 34.64035, 34.64132, 34.64244, 34.64309, 34.643, 34.6423, 
    34.64166, 34.64198, 34.64405, 34.64783, 34.65006, 34.65174, 34.65246, 
    34.6526, 34.65259, 34.65247, 34.65238, 34.65219, 34.65129, 34.6497, 
    34.6481, 34.64667, 34.64544, 34.64442, 34.64288, 34.63994, 34.63632, 
    34.63109, 34.62085, 34.60992, 34.60324, 34.59855, 34.59119, 34.58433, 
    34.5805, 34.57932, 34.58003, 34.58167, 34.58245, 34.58088, 34.5793, 
    34.58003, 34.58137, 34.58213, 34.5826, 34.58156, 34.57873, 34.57636, 
    34.57575, 34.57537, 34.57243, 34.56662, 34.56154, 34.56137,
  34.62986, 34.62959, 34.63039, 34.63132, 34.63181, 34.63161, 34.63083, 
    34.63012, 34.63029, 34.6321, 34.63557, 34.63958, 34.64267, 34.64409, 
    34.64451, 34.64469, 34.64471, 34.64479, 34.64469, 34.6433, 34.64064, 
    34.63797, 34.63561, 34.63363, 34.63209, 34.6296, 34.62569, 34.62217, 
    34.61713, 34.60744, 34.59549, 34.58455, 34.57701, 34.56902, 34.56242, 
    34.55862, 34.55729, 34.55771, 34.55899, 34.55949, 34.55779, 34.55612, 
    34.55663, 34.55769, 34.55826, 34.55862, 34.55754, 34.55484, 34.55262, 
    34.55199, 34.55161, 34.54888, 34.54347, 34.53874, 34.53857,
  34.61873, 34.61839, 34.61934, 34.62007, 34.6204, 34.62008, 34.61923, 
    34.61843, 34.61846, 34.62, 34.62306, 34.62663, 34.62933, 34.6305, 
    34.63074, 34.63076, 34.63061, 34.63051, 34.63025, 34.6288, 34.62618, 
    34.62355, 34.6212, 34.61919, 34.61757, 34.61507, 34.61128, 34.60784, 
    34.603, 34.58877, 34.57175, 34.56142, 34.55421, 34.54658, 34.54024, 
    34.53648, 34.535, 34.53513, 34.53605, 34.53626, 34.53444, 34.53266, 
    34.53294, 34.53372, 34.53411, 34.53435, 34.53323, 34.53068, 34.5286, 
    34.52796, 34.52758, 34.52506, 34.52004, 34.51566, 34.51549,
  34.59831, 34.59771, 34.5988, 34.6001, 34.60078, 34.60039, 34.5991, 
    34.59787, 34.59806, 34.60083, 34.60621, 34.61247, 34.61552, 34.61643, 
    34.61649, 34.61633, 34.616, 34.61572, 34.6153, 34.61378, 34.6112, 
    34.6086, 34.60622, 34.60316, 34.6008, 34.59698, 34.59099, 34.58557, 
    34.57785, 34.56298, 34.54716, 34.53745, 34.53058, 34.52055, 34.51167, 
    34.50657, 34.50476, 34.50529, 34.50697, 34.5076, 34.50534, 34.50311, 
    34.50377, 34.5052, 34.506, 34.50653, 34.50512, 34.50161, 34.49879, 
    34.49803, 34.4976, 34.49411, 34.48704, 34.48091, 34.48081,
  34.57694, 34.57608, 34.57672, 34.57755, 34.57782, 34.57714, 34.57566, 
    34.57422, 34.57407, 34.57626, 34.58078, 34.5861, 34.59011, 34.59181, 
    34.5921, 34.59206, 34.59179, 34.5916, 34.59116, 34.58891, 34.58489, 
    34.58084, 34.57723, 34.57415, 34.57168, 34.56792, 34.56219, 34.55697, 
    34.54969, 34.53598, 34.51475, 34.50105, 34.49154, 34.48153, 34.47318, 
    34.4682, 34.46618, 34.46623, 34.46733, 34.46747, 34.465, 34.46262, 
    34.4629, 34.46388, 34.46439, 34.46477, 34.46335, 34.46014, 34.45764, 
    34.45691, 34.45656, 34.45351, 34.44719, 34.44173, 34.44171,
  34.54314, 34.54183, 34.54301, 34.54457, 34.54527, 34.54446, 34.54239, 
    34.54037, 34.54042, 34.54417, 34.55154, 34.55867, 34.56186, 34.56302, 
    34.56293, 34.56256, 34.56197, 34.56145, 34.56073, 34.55841, 34.55452, 
    34.55061, 34.54706, 34.54396, 34.54138, 34.53651, 34.52851, 34.52127, 
    34.51114, 34.49185, 34.47144, 34.45895, 34.45016, 34.44093, 34.43313, 
    34.42829, 34.42603, 34.4256, 34.42608, 34.42571, 34.42303, 34.42049, 
    34.42038, 34.42089, 34.4211, 34.42133, 34.41989, 34.41699, 34.41483, 
    34.41414, 34.41386, 34.41128, 34.40484, 34.39811, 34.39823,
  34.5018, 34.49992, 34.50024, 34.50095, 34.50093, 34.49967, 34.49738, 
    34.49513, 34.49472, 34.49759, 34.50356, 34.51057, 34.51577, 34.51784, 
    34.51804, 34.51785, 34.51736, 34.51698, 34.51628, 34.51329, 34.50802, 
    34.50275, 34.49801, 34.49395, 34.49065, 34.48582, 34.47849, 34.47174, 
    34.46255, 34.44542, 34.42246, 34.40649, 34.39546, 34.38394, 34.3743, 
    34.36846, 34.36589, 34.36565, 34.3665, 34.36623, 34.36304, 34.36001, 
    34.36005, 34.36088, 34.36137, 34.3619, 34.36031, 34.35693, 34.35456, 
    34.35398, 34.35394, 34.35109, 34.34455, 34.33907, 34.33959,
  34.43709, 34.43472, 34.436, 34.43795, 34.43866, 34.43744, 34.43467, 34.432, 
    34.43212, 34.43712, 34.44666, 34.45756, 34.46562, 34.4671, 34.4669, 
    34.46639, 34.46566, 34.46501, 34.4641, 34.46131, 34.45659, 34.45102, 
    34.44497, 34.4399, 34.43589, 34.42992, 34.42066, 34.4122, 34.40068, 
    34.37897, 34.35615, 34.3424, 34.33279, 34.32271, 34.31418, 34.30876, 
    34.30599, 34.30519, 34.30527, 34.30432, 34.30088, 34.29771, 34.29725, 
    34.29746, 34.29764, 34.29809, 34.29663, 34.2939, 34.29223, 34.2919, 
    34.29219, 34.29026, 34.28421, 34.27821, 34.2792,
  34.36266, 34.35987, 34.36029, 34.36144, 34.36157, 34.36024, 34.3578, 
    34.35542, 34.35545, 34.35962, 34.36751, 34.37656, 34.38331, 34.38619, 
    34.38686, 34.3871, 34.38707, 34.38713, 34.38683, 34.38404, 34.37866, 
    34.37327, 34.36836, 34.36412, 34.36063, 34.35566, 34.34782, 34.34048, 
    34.33072, 34.30904, 34.28169, 34.26564, 34.2547, 34.24327, 34.2338, 
    34.22791, 34.22501, 34.22448, 34.22484, 34.22387, 34.21994, 34.21637, 
    34.21602, 34.21643, 34.2169, 34.21782, 34.2165, 34.2138, 34.21244, 
    34.21258, 34.2135, 34.21199, 34.20674, 34.20274, 34.20464,
  34.24461, 34.24247, 34.24482, 34.2481, 34.2499, 34.24958, 34.24766, 
    34.24577, 34.24714, 34.25404, 34.2658, 34.27899, 34.28899, 34.29382, 
    34.29573, 34.2971, 34.29811, 34.29927, 34.29993, 34.29747, 34.29171, 
    34.28596, 34.28085, 34.27655, 34.27312, 34.26797, 34.25926, 34.25113, 
    34.24019, 34.21917, 34.19719, 34.18443, 34.17298, 34.16026, 34.1499, 
    34.14359, 34.14059, 34.14038, 34.14113, 34.14023, 34.13591, 34.1321, 
    34.13208, 34.13288, 34.13383, 34.13536, 34.13438, 34.13194, 34.13104, 
    34.13178, 34.13341, 34.1324, 34.12734, 34.12371, 34.12656,
  34.1222, 34.12083, 34.12425, 34.12863, 34.13154, 34.13214, 34.13096, 
    34.12967, 34.13204, 34.14058, 34.15446, 34.17004, 34.18124, 34.18603, 
    34.18861, 34.19086, 34.19284, 34.195, 34.19686, 34.19635, 34.19311, 
    34.18976, 34.18529, 34.18139, 34.17836, 34.17336, 34.16412, 34.15549, 
    34.14358, 34.12006, 34.09563, 34.08174, 34.07253, 34.06279, 34.05499, 
    34.04993, 34.04702, 34.04637, 34.04633, 34.04483, 34.04063, 34.03733, 
    34.03751, 34.03843, 34.03987, 34.04219, 34.04239, 34.04155, 34.04203, 
    34.04376, 34.04627, 34.04678, 34.04411, 34.04266, 34.04645,
  34.00139, 34.00056, 34.00294, 34.00633, 34.00923, 34.01035, 34.01011, 
    34.00951, 34.012, 34.01954, 34.03099, 34.04391, 34.05425, 34.06042, 
    34.06429, 34.06792, 34.07108, 34.07459, 34.0779, 34.07838, 34.07568, 
    34.07274, 34.07029, 34.06815, 34.06639, 34.06311, 34.05643, 34.05011, 
    34.04116, 34.01411, 33.9856, 33.96902, 33.95795, 33.94613, 33.9367, 
    33.9304, 33.92657, 33.9254, 33.92569, 33.92477, 33.92084, 33.9189, 
    33.9222, 33.9267, 33.93148, 33.93703, 33.94013, 33.94128, 33.94313, 
    33.94679, 33.95062, 33.95159, 33.94969, 33.94875, 33.95308,
  33.92289, 33.91837, 33.91647, 33.91542, 33.91459, 33.913, 33.91084, 
    33.90807, 33.90845, 33.91372, 33.92237, 33.93279, 33.94151, 33.9469, 
    33.95042, 33.95386, 33.95668, 33.95992, 33.96305, 33.96313, 33.95977, 
    33.9558, 33.95234, 33.94912, 33.9463, 33.94133, 33.93296, 33.92548, 
    33.91397, 33.89251, 33.86334, 33.84093, 33.82548, 33.80889, 33.79521, 
    33.78562, 33.77946, 33.77655, 33.77714, 33.77733, 33.7737, 33.77407, 
    33.78301, 33.79387, 33.80454, 33.81572, 33.8236, 33.8277, 33.83149, 
    33.83813, 33.84398, 33.8452, 33.84356, 33.84259, 33.84758,
  33.92331, 33.90643, 33.89128, 33.87834, 33.86725, 33.85801, 33.85031, 
    33.84176, 33.8367, 33.8365, 33.83887, 33.8436, 33.84813, 33.85064, 
    33.85183, 33.85296, 33.8535, 33.85423, 33.85471, 33.85211, 33.84566, 
    33.83799, 33.83055, 33.82351, 33.81721, 33.80758, 33.79481, 33.7841, 
    33.7665, 33.73709, 33.70829, 33.68719, 33.66666, 33.64487, 33.62616, 
    33.61201, 33.60177, 33.59489, 33.59433, 33.59521, 33.59163, 33.59509, 
    33.61146, 33.63031, 33.6489, 33.66804, 33.68269, 33.69103, 33.69769, 
    33.70825, 33.71682, 33.71832, 33.71645, 33.71515, 33.72155,
  33.99631, 33.95935, 33.92434, 33.89379, 33.86636, 33.84441, 33.82714, 
    33.80901, 33.79541, 33.7874, 33.78128, 33.77829, 33.77668, 33.77424, 
    33.7707, 33.76693, 33.76275, 33.75812, 33.75261, 33.74448, 33.73198, 
    33.71762, 33.70279, 33.68901, 33.67675, 33.65981, 33.641, 33.62611, 
    33.60071, 33.56314, 33.52752, 33.50014, 33.47957, 33.45748, 33.43392, 
    33.41426, 33.39798, 33.38453, 33.38055, 33.38079, 33.3758, 33.38168, 
    33.40536, 33.43116, 33.45784, 33.48613, 33.50818, 33.52076, 33.53041, 
    33.54487, 33.55642, 33.55755, 33.55325, 33.55056, 33.56034,
  34.13303, 34.0731, 34.01531, 33.96374, 33.91568, 33.87708, 33.84686, 
    33.81636, 33.79094, 33.77111, 33.75206, 33.73684, 33.72511, 33.71479, 
    33.7039, 33.69268, 33.68105, 33.66835, 33.65417, 33.63851, 33.61801, 
    33.59501, 33.57016, 33.54763, 33.52802, 33.50229, 33.4771, 33.45821, 
    33.42498, 33.38151, 33.34154, 33.30777, 33.28136, 33.25509, 33.2271, 
    33.20052, 33.1762, 33.15354, 33.14271, 33.13873, 33.12806, 33.13127, 
    33.15535, 33.17673, 33.20188, 33.23268, 33.25894, 33.2773, 33.28921, 
    33.30568, 33.31937, 33.31887, 33.30792, 33.30148, 33.31736,
  34.32937, 34.25089, 34.17238, 34.0991, 34.03009, 33.97298, 33.92657, 
    33.88124, 33.8401, 33.80319, 33.76613, 33.73307, 33.70506, 33.68171, 
    33.65881, 33.63594, 33.61159, 33.58669, 33.56086, 33.53441, 33.50376, 
    33.471, 33.43528, 33.40416, 33.37813, 33.34385, 33.31306, 33.29053, 
    33.25026, 33.20224, 33.15749, 33.1165, 33.08328, 33.05042, 33.015, 
    32.98298, 32.95462, 32.92561, 32.909, 32.90129, 32.88645, 32.88266, 
    32.89293, 32.89162, 32.89595, 32.907, 32.91954, 32.92974, 32.94051, 
    32.94865, 32.9558, 32.95344, 32.94054, 32.93188, 32.94391,
  34.45667, 34.36971, 34.28521, 34.20415, 34.12684, 34.05975, 34.0027, 
    33.94899, 33.89865, 33.85156, 33.80499, 33.75872, 33.71383, 33.67323, 
    33.63382, 33.5954, 33.55415, 33.51432, 33.47557, 33.4361, 33.39445, 
    33.35275, 33.309, 33.2724, 33.24319, 33.2028, 33.16763, 33.14093, 
    33.09695, 33.04628, 32.99461, 32.94804, 32.91692, 32.88907, 32.8552, 
    32.82768, 32.80669, 32.78162, 32.76944, 32.77005, 32.77024, 32.77508, 
    32.78465, 32.79096, 32.78986, 32.78136, 32.77874, 32.76873, 32.75139, 
    32.73983, 32.7269, 32.71246, 32.6991, 32.68863, 32.68126,
  34.47111, 34.38123, 34.29589, 34.21503, 34.13678, 34.06878, 34.01099, 
    33.95726, 33.90652, 33.85883, 33.81294, 33.76471, 33.71416, 33.664, 
    33.61371, 33.56335, 33.5111, 33.46045, 33.41142, 33.36197, 33.31533, 
    33.27194, 33.22969, 33.19601, 33.17094, 33.1342, 33.10456, 33.08218, 
    33.046, 33.0116, 32.97892, 32.94334, 32.91118, 32.88224, 32.84669, 
    32.81888, 32.7988, 32.77494, 32.7636, 32.76474, 32.76573, 32.77114, 
    32.78098, 32.78788, 32.78705, 32.77848, 32.77588, 32.76565, 32.7478, 
    32.73604, 32.72283, 32.70813, 32.69493, 32.68428, 32.67618,
  34.47064, 34.37995, 34.29424, 34.21351, 34.13506, 34.06686, 34.00892, 
    33.95497, 33.90419, 33.85656, 33.81095, 33.76272, 33.71188, 33.66126, 
    33.6097, 33.55723, 33.50448, 33.45195, 33.39963, 33.34869, 33.30154, 
    33.25816, 33.21759, 33.18615, 33.16385, 33.12933, 33.10136, 33.07995, 
    33.04421, 33.01004, 32.9775, 32.94222, 32.91009, 32.88105, 32.84549, 
    32.81775, 32.79781, 32.774, 32.76276, 32.76407, 32.76501, 32.77039, 
    32.78022, 32.78711, 32.78625, 32.77765, 32.77498, 32.76471, 32.74681, 
    32.7351, 32.72198, 32.70747, 32.69439, 32.68378, 32.67564,
  34.46987, 34.37873, 34.29281, 34.2121, 34.13366, 34.06553, 34.00773, 
    33.95391, 33.90318, 33.85553, 33.81, 33.7618, 33.71093, 33.66036, 
    33.6088, 33.55627, 33.50349, 33.45094, 33.3986, 33.34768, 33.30051, 
    33.2571, 33.21655, 33.18517, 33.16294, 33.12846, 33.10045, 33.07893, 
    33.04316, 33.00904, 32.9766, 32.94132, 32.90908, 32.87984, 32.84396, 
    32.81614, 32.79639, 32.77264, 32.76156, 32.76313, 32.76423, 32.76976, 
    32.77971, 32.78664, 32.7858, 32.7772, 32.77454, 32.76426, 32.74639, 
    32.73471, 32.72163, 32.70715, 32.69409, 32.68349, 32.67534,
  34.46923, 34.37754, 34.29137, 34.21074, 34.13223, 34.06419, 34.00662, 
    33.95303, 33.90239, 33.85471, 33.80918, 33.76094, 33.71001, 33.6594, 
    33.60778, 33.55517, 33.50237, 33.4497, 33.39716, 33.34621, 33.29897, 
    33.25544, 33.21487, 33.18349, 33.16127, 33.12683, 33.09893, 33.07757, 
    33.04193, 33.00797, 32.9757, 32.94049, 32.9082, 32.87884, 32.84282, 
    32.81494, 32.79519, 32.77139, 32.76038, 32.76217, 32.76346, 32.76912, 
    32.77915, 32.78615, 32.78534, 32.77673, 32.7741, 32.76386, 32.74601, 
    32.73438, 32.72134, 32.70689, 32.69385, 32.68325, 32.6751,
  34.68758, 34.68752, 34.68773, 34.688, 34.68818, 34.68819, 34.68806, 
    34.68793, 34.68803, 34.68833, 34.68867, 34.68906, 34.68935, 34.68949, 
    34.68953, 34.68957, 34.68959, 34.68963, 34.68966, 34.68953, 34.68927, 
    34.68902, 34.6888, 34.68864, 34.68855, 34.68827, 34.6878, 34.68737, 
    34.68641, 34.68388, 34.68106, 34.67865, 34.67698, 34.67522, 34.67374, 
    34.67294, 34.67267, 34.67268, 34.67285, 34.67289, 34.67255, 34.6722, 
    34.67221, 34.67233, 34.67235, 34.67232, 34.67207, 34.67151, 34.67102, 
    34.6708, 34.67064, 34.67002, 34.66889, 34.66785, 34.66774,
  34.6845, 34.68443, 34.68469, 34.68489, 34.68498, 34.68494, 34.68478, 
    34.68462, 34.68468, 34.68512, 34.68591, 34.68682, 34.68753, 34.68785, 
    34.68791, 34.68788, 34.68781, 34.68776, 34.68773, 34.68755, 34.68711, 
    34.68655, 34.68605, 34.68565, 34.68536, 34.68481, 34.68394, 34.68317, 
    34.68196, 34.67879, 34.67515, 34.67299, 34.67109, 34.66887, 34.66705, 
    34.66604, 34.66574, 34.66589, 34.66627, 34.6664, 34.66592, 34.66544, 
    34.66556, 34.66584, 34.66596, 34.66601, 34.66564, 34.66479, 34.66402, 
    34.66373, 34.66351, 34.66264, 34.66102, 34.6596, 34.65948,
  34.67998, 34.6799, 34.68021, 34.68056, 34.68074, 34.6807, 34.68047, 
    34.68026, 34.68037, 34.68105, 34.68225, 34.68362, 34.68428, 34.68452, 
    34.68454, 34.68451, 34.68443, 34.68438, 34.68433, 34.68398, 34.68338, 
    34.68281, 34.6823, 34.68178, 34.68135, 34.68058, 34.67938, 34.67831, 
    34.67669, 34.67352, 34.66895, 34.66615, 34.6642, 34.66212, 34.66042, 
    34.65941, 34.65903, 34.65921, 34.65949, 34.65954, 34.65901, 34.65849, 
    34.65852, 34.65869, 34.65873, 34.65872, 34.65832, 34.65749, 34.65675, 
    34.65644, 34.65622, 34.6554, 34.65309, 34.65077, 34.65063,
  34.67511, 34.67502, 34.67548, 34.676, 34.6763, 34.67627, 34.67598, 34.6757, 
    34.67588, 34.67684, 34.67798, 34.67921, 34.68014, 34.68052, 34.68058, 
    34.68057, 34.68048, 34.68044, 34.68037, 34.6799, 34.67907, 34.67828, 
    34.67758, 34.67699, 34.67652, 34.67575, 34.67457, 34.67347, 34.67135, 
    34.66716, 34.66275, 34.65964, 34.65649, 34.65311, 34.65034, 34.64879, 
    34.64833, 34.64861, 34.64924, 34.6495, 34.64879, 34.64808, 34.6483, 
    34.64876, 34.64898, 34.64908, 34.64856, 34.6473, 34.6462, 34.64583, 
    34.64556, 34.64426, 34.64179, 34.63962, 34.63947,
  34.66994, 34.66985, 34.67025, 34.67072, 34.67096, 34.6709, 34.6706, 
    34.67033, 34.67048, 34.67135, 34.67292, 34.67469, 34.67602, 34.67655, 
    34.67657, 34.67651, 34.67639, 34.6763, 34.6762, 34.67572, 34.6749, 
    34.67382, 34.67287, 34.67207, 34.67145, 34.67044, 34.66887, 34.66744, 
    34.66541, 34.66149, 34.65442, 34.65006, 34.64703, 34.64379, 34.64111, 
    34.63958, 34.63906, 34.63922, 34.63971, 34.63985, 34.63908, 34.63832, 
    34.63846, 34.63881, 34.63895, 34.63899, 34.63847, 34.63726, 34.6362, 
    34.63582, 34.63554, 34.63431, 34.632, 34.62969, 34.62951,
  34.66392, 34.66381, 34.6645, 34.66529, 34.66576, 34.66573, 34.66532, 
    34.66495, 34.66523, 34.66653, 34.66798, 34.66961, 34.67082, 34.67133, 
    34.67142, 34.6714, 34.6713, 34.67125, 34.67115, 34.67053, 34.66945, 
    34.6684, 34.66747, 34.66668, 34.66604, 34.66505, 34.66352, 34.66214, 
    34.6591, 34.65266, 34.6458, 34.64165, 34.63873, 34.63353, 34.62897, 
    34.62647, 34.62578, 34.62632, 34.62747, 34.62803, 34.627, 34.62595, 
    34.62646, 34.62735, 34.62783, 34.62812, 34.6274, 34.62545, 34.62377, 
    34.62329, 34.62295, 34.62088, 34.6169, 34.6134, 34.61321,
  34.65704, 34.65691, 34.65752, 34.65822, 34.65861, 34.65854, 34.6581, 
    34.65772, 34.65794, 34.65925, 34.66161, 34.6643, 34.66617, 34.66662, 
    34.66667, 34.66661, 34.66648, 34.66639, 34.66625, 34.66563, 34.66459, 
    34.66351, 34.66208, 34.66088, 34.65997, 34.65845, 34.65603, 34.65384, 
    34.65068, 34.64458, 34.63693, 34.62965, 34.62465, 34.61933, 34.61494, 
    34.61247, 34.61169, 34.61206, 34.61301, 34.61341, 34.61231, 34.61122, 
    34.6116, 34.61232, 34.61269, 34.6129, 34.61216, 34.61029, 34.60868, 
    34.60817, 34.60782, 34.60587, 34.60212, 34.59882, 34.59862,
  34.65073, 34.65059, 34.65112, 34.65173, 34.65205, 34.65194, 34.65149, 
    34.65109, 34.65126, 34.65244, 34.65461, 34.65707, 34.65892, 34.65973, 
    34.65992, 34.65995, 34.65989, 34.65987, 34.65975, 34.65886, 34.65724, 
    34.65564, 34.65422, 34.65301, 34.65205, 34.65053, 34.64817, 34.64602, 
    34.64296, 34.63466, 34.62316, 34.61623, 34.61141, 34.6063, 34.60206, 
    34.59962, 34.59876, 34.59898, 34.59974, 34.6, 34.59883, 34.5977, 
    34.59796, 34.59853, 34.5988, 34.59893, 34.59818, 34.59638, 34.59483, 
    34.5943, 34.59393, 34.59209, 34.58855, 34.58519, 34.58497,
  34.64046, 34.64025, 34.64122, 34.64235, 34.64301, 34.64294, 34.64225, 
    34.64164, 34.642, 34.64415, 34.64798, 34.65023, 34.65191, 34.65262, 
    34.65273, 34.65269, 34.65256, 34.65246, 34.65227, 34.65135, 34.64976, 
    34.64818, 34.64677, 34.64555, 34.64455, 34.64303, 34.64009, 34.63646, 
    34.63122, 34.62099, 34.61013, 34.60351, 34.59887, 34.59159, 34.58477, 
    34.58101, 34.57991, 34.58065, 34.58232, 34.58315, 34.58162, 34.58009, 
    34.58085, 34.58219, 34.58294, 34.5834, 34.58237, 34.57953, 34.57713, 
    34.57645, 34.576, 34.57301, 34.56715, 34.56202, 34.56178,
  34.62974, 34.62946, 34.63026, 34.6312, 34.63169, 34.6315, 34.63075, 
    34.63006, 34.63028, 34.63217, 34.6357, 34.63975, 34.64283, 34.64425, 
    34.64465, 34.6448, 34.64481, 34.64487, 34.64476, 34.64336, 34.64071, 
    34.63804, 34.63571, 34.63375, 34.63222, 34.62975, 34.62585, 34.62231, 
    34.61726, 34.6076, 34.59571, 34.58485, 34.57738, 34.56948, 34.56293, 
    34.55921, 34.55797, 34.55844, 34.55978, 34.56034, 34.5587, 34.55708, 
    34.55762, 34.55869, 34.55926, 34.5596, 34.55853, 34.55581, 34.55354, 
    34.55283, 34.55237, 34.54958, 34.54409, 34.5393, 34.53906,
  34.61858, 34.61821, 34.61916, 34.6199, 34.62024, 34.61994, 34.61911, 
    34.61834, 34.61843, 34.62005, 34.62318, 34.62677, 34.62947, 34.63064, 
    34.63087, 34.63085, 34.6307, 34.63058, 34.63032, 34.62885, 34.62624, 
    34.62362, 34.62129, 34.6193, 34.6177, 34.61523, 34.61145, 34.60799, 
    34.60314, 34.58895, 34.57202, 34.56176, 34.55463, 34.54711, 34.54082, 
    34.53715, 34.53578, 34.53597, 34.53697, 34.53726, 34.5355, 34.53379, 
    34.53411, 34.53491, 34.53529, 34.53551, 34.53439, 34.53181, 34.52967, 
    34.52893, 34.52845, 34.52587, 34.52077, 34.51631, 34.51607,
  34.59812, 34.5975, 34.59858, 34.59989, 34.60058, 34.6002, 34.59894, 
    34.59774, 34.59798, 34.60084, 34.6063, 34.61259, 34.61563, 34.61655, 
    34.61659, 34.6164, 34.61607, 34.61578, 34.61536, 34.61382, 34.61125, 
    34.60867, 34.60631, 34.60328, 34.60094, 34.59716, 34.59118, 34.58574, 
    34.57802, 34.56319, 34.54747, 34.53783, 34.53106, 34.52114, 34.51234, 
    34.50735, 34.50568, 34.50629, 34.50807, 34.5088, 34.50663, 34.50447, 
    34.50518, 34.50662, 34.50741, 34.50791, 34.50649, 34.50294, 34.50005, 
    34.49917, 34.49864, 34.49506, 34.48791, 34.4817, 34.4815,
  34.57671, 34.57582, 34.57645, 34.57729, 34.57758, 34.57692, 34.57545, 
    34.57405, 34.57396, 34.57623, 34.58082, 34.58616, 34.59016, 34.59187, 
    34.59215, 34.59209, 34.59182, 34.59163, 34.59119, 34.58894, 34.58492, 
    34.58089, 34.57733, 34.57428, 34.57185, 34.56812, 34.56241, 34.55718, 
    34.5499, 34.53624, 34.51513, 34.50153, 34.49213, 34.48226, 34.47399, 
    34.46914, 34.46729, 34.46746, 34.46868, 34.46896, 34.4666, 34.46431, 
    34.46465, 34.46564, 34.46615, 34.46649, 34.46503, 34.46177, 34.45917, 
    34.4583, 34.45781, 34.45465, 34.44822, 34.44267, 34.44254,
  34.54284, 34.5415, 34.54269, 34.54427, 34.54499, 34.54419, 34.54214, 
    34.54017, 34.54027, 34.54408, 34.55151, 34.55867, 34.56183, 34.563, 
    34.56291, 34.56253, 34.56194, 34.56143, 34.56072, 34.55841, 34.55455, 
    34.55067, 34.54717, 34.54411, 34.54158, 34.53675, 34.52878, 34.52155, 
    34.51143, 34.49223, 34.47193, 34.45955, 34.45088, 34.4418, 34.43409, 
    34.4294, 34.42735, 34.42706, 34.4277, 34.42751, 34.42496, 34.42253, 
    34.42248, 34.42302, 34.42323, 34.4234, 34.42191, 34.41893, 34.41665, 
    34.41578, 34.41534, 34.41262, 34.40606, 34.39921, 34.39921,
  34.50141, 34.49951, 34.49985, 34.5006, 34.50061, 34.49937, 34.4971, 
    34.4949, 34.49453, 34.49742, 34.50342, 34.51042, 34.51557, 34.51765, 
    34.51786, 34.51768, 34.51722, 34.51687, 34.5162, 34.51325, 34.50803, 
    34.50282, 34.49816, 34.49416, 34.49093, 34.48616, 34.47887, 34.47215, 
    34.46297, 34.44592, 34.4231, 34.40724, 34.39635, 34.385, 34.37547, 
    34.36981, 34.36749, 34.36745, 34.36852, 34.36848, 34.36547, 34.36258, 
    34.36269, 34.36355, 34.36402, 34.36448, 34.3628, 34.35931, 34.35677, 
    34.35596, 34.35571, 34.35268, 34.34598, 34.34036, 34.34073,
  34.43657, 34.43421, 34.43554, 34.43755, 34.43831, 34.43711, 34.43435, 
    34.43171, 34.43184, 34.43682, 34.44636, 34.45724, 34.46524, 34.46672, 
    34.46654, 34.46606, 34.46537, 34.46478, 34.46393, 34.46122, 34.45659, 
    34.45111, 34.44517, 34.4402, 34.43627, 34.43039, 34.42121, 34.41278, 
    34.40131, 34.37971, 34.35702, 34.34336, 34.33387, 34.32398, 34.31555, 
    34.31034, 34.30789, 34.30735, 34.3077, 34.30706, 34.30383, 34.30082, 
    34.30046, 34.30071, 34.30085, 34.30122, 34.29963, 34.29674, 34.29486, 
    34.29424, 34.29426, 34.2921, 34.28587, 34.2797, 34.2805,
  34.36198, 34.35925, 34.35974, 34.36099, 34.36119, 34.35989, 34.35742, 
    34.35506, 34.35505, 34.35912, 34.36692, 34.37589, 34.38252, 34.38539, 
    34.3861, 34.38644, 34.38649, 34.38666, 34.38648, 34.38385, 34.37863, 
    34.37341, 34.36866, 34.36456, 34.36119, 34.35636, 34.34861, 34.34132, 
    34.33161, 34.31004, 34.28282, 34.26683, 34.25602, 34.24479, 34.2354, 
    34.22978, 34.2273, 34.22715, 34.22791, 34.22738, 34.22374, 34.22039, 
    34.22017, 34.22061, 34.22104, 34.22183, 34.22032, 34.2174, 34.21577, 
    34.2155, 34.21605, 34.21422, 34.20872, 34.20448, 34.20614,
  34.24387, 34.2418, 34.24423, 34.24759, 34.24943, 34.24909, 34.24708, 
    34.24517, 34.24645, 34.25317, 34.26481, 34.27789, 34.28776, 34.29258, 
    34.29457, 34.29612, 34.29727, 34.29858, 34.29945, 34.29724, 34.29173, 
    34.28624, 34.28134, 34.27723, 34.27398, 34.269, 34.26042, 34.25235, 
    34.24147, 34.22055, 34.19863, 34.18587, 34.17451, 34.162, 34.1517, 
    34.14572, 34.1433, 34.14364, 34.14496, 34.14469, 34.14077, 34.13725, 
    34.13736, 34.13819, 34.13906, 34.14042, 34.13917, 34.13646, 34.13525, 
    34.13545, 34.1366, 34.13519, 34.12984, 34.12592, 34.12845,
  34.12169, 34.12035, 34.1238, 34.12821, 34.1311, 34.13161, 34.13029, 
    34.12896, 34.13119, 34.13949, 34.15316, 34.16853, 34.17955, 34.18435, 
    34.18708, 34.18963, 34.19181, 34.1942, 34.19634, 34.19618, 34.19327, 
    34.19024, 34.18605, 34.18239, 34.17958, 34.17478, 34.16569, 34.15712, 
    34.14524, 34.12172, 34.0972, 34.08322, 34.0741, 34.06464, 34.0569, 
    34.05228, 34.05021, 34.0504, 34.05124, 34.05071, 34.04708, 34.04416, 
    34.04449, 34.04543, 34.04678, 34.04889, 34.04868, 34.04745, 34.04756, 
    34.0486, 34.0505, 34.05047, 34.0474, 34.04556, 34.04892,
  34.00134, 34.00043, 34.00281, 34.00621, 34.009, 34.00996, 34.00953, 
    34.0089, 34.01128, 34.01862, 34.02995, 34.04277, 34.05305, 34.05933, 
    34.06345, 34.06747, 34.07087, 34.07462, 34.07818, 34.079, 34.07663, 
    34.07398, 34.07173, 34.06978, 34.0682, 34.06506, 34.05846, 34.05214, 
    34.04314, 34.01575, 33.98671, 33.9699, 33.95903, 33.94785, 33.93866, 
    33.93333, 33.9312, 33.93186, 33.93393, 33.93481, 33.93193, 33.93059, 
    33.93388, 33.93817, 33.94262, 33.94769, 33.94999, 33.95051, 33.9518, 
    33.95438, 33.95725, 33.95748, 33.95502, 33.95353, 33.95723,
  33.92232, 33.91744, 33.91543, 33.91449, 33.91358, 33.91198, 33.90988, 
    33.90739, 33.90797, 33.91334, 33.92212, 33.93259, 33.94135, 33.94703, 
    33.95094, 33.95481, 33.95786, 33.96126, 33.96451, 33.96482, 33.96165, 
    33.95778, 33.9543, 33.9511, 33.94834, 33.94327, 33.93472, 33.92698, 
    33.91521, 33.89328, 33.86343, 33.84103, 33.82634, 33.81131, 33.79848, 
    33.7909, 33.78785, 33.78849, 33.79226, 33.79551, 33.79368, 33.79493, 
    33.80347, 33.81364, 33.8235, 33.83372, 33.84015, 33.8432, 33.84609, 
    33.85101, 33.85532, 33.8554, 33.85296, 33.85114, 33.85509,
  33.9174, 33.9003, 33.88559, 33.87356, 33.86316, 33.8547, 33.84792, 
    33.84043, 33.83631, 33.83687, 33.83978, 33.84473, 33.84932, 33.85237, 
    33.85406, 33.85566, 33.85624, 33.85698, 33.85743, 33.85487, 33.8484, 
    33.84063, 33.833, 33.82582, 33.81941, 33.80953, 33.79635, 33.78505, 
    33.76731, 33.73742, 33.70768, 33.6872, 33.66859, 33.64992, 33.63306, 
    33.6223, 33.61699, 33.61604, 33.62061, 33.62618, 33.62499, 33.62937, 
    33.64476, 33.66216, 33.67943, 33.69726, 33.70963, 33.71636, 33.72179, 
    33.72982, 33.73609, 33.73583, 33.73278, 33.73027, 33.73506,
  33.98709, 33.9506, 33.91687, 33.88834, 33.86295, 33.84318, 33.8283, 
    33.81231, 33.8003, 33.79313, 33.78684, 33.78313, 33.78065, 33.77865, 
    33.77555, 33.7721, 33.76734, 33.76238, 33.75678, 33.74847, 33.73589, 
    33.72149, 33.70656, 33.69261, 33.68008, 33.66293, 33.6436, 33.62774, 
    33.60275, 33.56517, 33.52875, 33.50332, 33.48591, 33.46816, 33.4465, 
    33.43106, 33.42128, 33.41674, 33.42039, 33.42709, 33.42381, 33.42962, 
    33.45168, 33.47489, 33.5002, 33.5282, 33.54729, 33.55761, 33.56611, 
    33.57738, 33.58585, 33.58386, 33.57664, 33.57113, 33.57859,
  34.13664, 34.07759, 34.02061, 33.97049, 33.92485, 33.88913, 33.86214, 
    33.83368, 33.80939, 33.78962, 33.76847, 33.75075, 33.73646, 33.72611, 
    33.71526, 33.70397, 33.6904, 33.6767, 33.66248, 33.64605, 33.62516, 
    33.60204, 33.57709, 33.55408, 33.5336, 33.50724, 33.48055, 33.45929, 
    33.42593, 33.38074, 33.33777, 33.30602, 33.28345, 33.26265, 33.23636, 
    33.21398, 33.19655, 33.18562, 33.18418, 33.18705, 33.17422, 33.17416, 
    33.19446, 33.2094, 33.23204, 33.26442, 33.28793, 33.30638, 33.32102, 
    33.33442, 33.34469, 33.34, 33.32467, 33.31378, 33.32598,
  34.33096, 34.25303, 34.17707, 34.10738, 34.04207, 33.98875, 33.94643, 
    33.90327, 33.86402, 33.82874, 33.78993, 33.75399, 33.72195, 33.69807, 
    33.67468, 33.65165, 33.62433, 33.59803, 33.57236, 33.54472, 33.51274, 
    33.47873, 33.4416, 33.4082, 33.37904, 33.34228, 33.30716, 33.279, 
    33.23647, 33.18302, 33.13168, 33.09303, 33.06459, 33.0376, 33.00483, 
    32.97723, 32.95464, 32.93915, 32.93277, 32.93118, 32.91155, 32.90282, 
    32.90864, 32.90376, 32.90702, 32.91959, 32.93072, 32.94129, 32.95494, 
    32.96152, 32.96661, 32.96123, 32.94411, 32.93177, 32.94015,
  34.41564, 34.32846, 34.24817, 34.1746, 34.10335, 34.04344, 33.99494, 
    33.9463, 33.90174, 33.86112, 33.81639, 33.76884, 33.71932, 33.6792, 
    33.63991, 33.60136, 33.55721, 33.51549, 33.4758, 33.43389, 33.38964, 
    33.34574, 33.29905, 33.25747, 33.22123, 33.17663, 33.13444, 33.09858, 
    33.05162, 32.99555, 32.9389, 32.89831, 32.87431, 32.85277, 32.8244, 
    32.80099, 32.78272, 32.76619, 32.76054, 32.76555, 32.76531, 32.76863, 
    32.77588, 32.77827, 32.77528, 32.76704, 32.76294, 32.75411, 32.7406, 
    32.73006, 32.71892, 32.70693, 32.69558, 32.68758, 32.68339,
  34.41077, 34.32056, 34.23909, 34.16618, 34.09525, 34.03664, 33.9904, 
    33.94404, 33.90057, 33.86008, 33.81776, 33.77123, 33.72054, 33.67418, 
    33.6253, 33.57401, 33.51389, 33.45827, 33.40708, 33.34946, 33.29705, 
    33.25015, 33.20437, 33.16413, 33.12948, 33.0876, 33.05013, 33.01751, 
    32.98124, 32.94556, 32.9105, 32.88231, 32.85691, 32.83351, 32.804, 
    32.78141, 32.76575, 32.75033, 32.74437, 32.74786, 32.74888, 32.75365, 
    32.76221, 32.76756, 32.76651, 32.75906, 32.7569, 32.74832, 32.73335, 
    32.72388, 32.71242, 32.69896, 32.68774, 32.6787, 32.67185,
  34.40595, 34.31359, 34.23145, 34.15941, 34.08914, 34.03116, 33.9855, 
    33.94035, 33.89724, 33.85619, 33.81394, 33.76669, 33.71442, 33.66722, 
    33.61696, 33.5637, 33.50187, 33.4446, 33.39187, 33.33371, 33.28041, 
    33.23202, 33.18804, 33.15012, 33.11826, 33.0784, 33.04274, 33.01125, 
    32.97676, 32.94268, 32.90903, 32.88137, 32.85577, 32.83221, 32.80251, 
    32.77982, 32.76418, 32.7488, 32.74287, 32.74639, 32.74695, 32.75146, 
    32.75995, 32.76602, 32.76535, 32.75795, 32.75583, 32.74731, 32.73243, 
    32.72299, 32.71156, 32.69813, 32.6871, 32.67815, 32.67131,
  34.40304, 34.30877, 34.22594, 34.15447, 34.08439, 34.02679, 33.98167, 
    33.93755, 33.89489, 33.85372, 33.8116, 33.76412, 33.71129, 33.66394, 
    33.6137, 33.56057, 33.49834, 33.44101, 33.38855, 33.33065, 33.27771, 
    33.22976, 33.18639, 33.14898, 33.11749, 33.07817, 33.04284, 33.01147, 
    32.97693, 32.94282, 32.9091, 32.8811, 32.85519, 32.83138, 32.80132, 
    32.77834, 32.76242, 32.74707, 32.74086, 32.74376, 32.74423, 32.74862, 
    32.75695, 32.76313, 32.76264, 32.75547, 32.75377, 32.74561, 32.73098, 
    32.72183, 32.71059, 32.69725, 32.68639, 32.67756, 32.67076,
  34.40163, 34.30633, 34.22304, 34.15175, 34.08188, 34.02453, 33.9797, 
    33.93613, 33.89362, 33.85217, 33.80995, 33.76218, 33.70883, 33.66071, 
    33.61006, 33.55687, 33.49448, 33.43718, 33.38499, 33.3274, 33.27485, 
    33.22734, 33.18469, 33.14791, 33.117, 33.07812, 33.04307, 33.01184, 
    32.97722, 32.94296, 32.90907, 32.88084, 32.85469, 32.8306, 32.80037, 
    32.77716, 32.76099, 32.74557, 32.73926, 32.74204, 32.74245, 32.74662, 
    32.75455, 32.76033, 32.75992, 32.75333, 32.75178, 32.74389, 32.72968, 
    32.72075, 32.70966, 32.6964, 32.68584, 32.67718, 32.67041 ;

 salt_east =
  33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647 ;

 salt_south =
  34.68758, 34.6876, 34.68762, 34.68786, 34.68828, 34.68855, 34.68845, 
    34.68811, 34.68796, 34.68806, 34.68829, 34.68839, 34.68825, 34.68789, 
    34.68766, 34.68767, 34.68752, 34.68697, 34.68634, 34.68613, 34.68631, 
    34.68652, 34.68665, 34.68656, 34.68597, 34.68522, 34.68488, 34.68486, 
    34.68483, 34.68476, 34.6846, 34.68422, 34.68344, 34.68255, 34.68195, 
    34.68182, 34.68198, 34.68206, 34.68188, 34.68151, 34.68095, 34.68005, 
    34.67893, 34.67787, 34.67635, 34.67298, 34.6637, 34.64002, 34.59103, 
    34.52918, 34.47678, 34.42651, 34.35043, 34.24358, 34.15375, 33.97319,
  34.6845, 34.68452, 34.68455, 34.68486, 34.68526, 34.6855, 34.68536, 
    34.68507, 34.68484, 34.68489, 34.68505, 34.68511, 34.68496, 34.68442, 
    34.68404, 34.68401, 34.68376, 34.68299, 34.68217, 34.68189, 34.68209, 
    34.68234, 34.68249, 34.68238, 34.68172, 34.68092, 34.68058, 34.68058, 
    34.68059, 34.68055, 34.68042, 34.68006, 34.67938, 34.67859, 34.67781, 
    34.67767, 34.67793, 34.67807, 34.67783, 34.6773, 34.67654, 34.67531, 
    34.67379, 34.6726, 34.67128, 34.6666, 34.65553, 34.62691, 34.57379, 
    34.51165, 34.46203, 34.41224, 34.32589, 34.20141, 34.09222, 33.97319,
  34.67997, 34.68001, 34.68005, 34.68041, 34.68104, 34.6814, 34.68116, 
    34.68068, 34.68041, 34.68045, 34.68069, 34.68078, 34.68057, 34.68004, 
    34.6797, 34.67969, 34.67949, 34.67881, 34.67792, 34.67754, 34.67786, 
    34.67825, 34.67849, 34.67838, 34.67744, 34.67628, 34.67582, 34.67587, 
    34.67593, 34.67591, 34.67577, 34.67528, 34.67431, 34.67318, 34.67245, 
    34.67237, 34.67266, 34.67284, 34.67266, 34.67223, 34.67158, 34.6705, 
    34.66856, 34.66646, 34.66408, 34.65862, 34.64353, 34.61053, 34.55389, 
    34.49565, 34.44513, 34.3849, 34.29059, 34.16533, 34.03954, 33.97319,
  34.6751, 34.67514, 34.67519, 34.6757, 34.67657, 34.67706, 34.67672, 
    34.67599, 34.67561, 34.6757, 34.67604, 34.67618, 34.67588, 34.67512, 
    34.67464, 34.67463, 34.67432, 34.67332, 34.67226, 34.67193, 34.67226, 
    34.67265, 34.67292, 34.67283, 34.672, 34.67097, 34.67059, 34.67068, 
    34.67078, 34.6708, 34.67072, 34.67031, 34.66947, 34.66788, 34.66661, 
    34.66648, 34.66699, 34.66729, 34.667, 34.66626, 34.66512, 34.6632, 
    34.66079, 34.65891, 34.65676, 34.6501, 34.6316, 34.59396, 34.53679, 
    34.48189, 34.4306, 34.35955, 34.24897, 34.11459, 33.99417, 33.97319,
  34.66994, 34.66998, 34.67002, 34.67049, 34.6713, 34.67176, 34.67144, 
    34.67076, 34.6704, 34.67048, 34.67079, 34.67091, 34.67064, 34.66993, 
    34.66949, 34.66949, 34.66922, 34.66832, 34.66685, 34.66628, 34.6668, 
    34.66745, 34.6679, 34.66775, 34.66634, 34.66456, 34.66389, 34.66403, 
    34.66419, 34.66422, 34.66406, 34.66335, 34.66186, 34.6601, 34.65898, 
    34.65892, 34.65945, 34.65979, 34.65958, 34.65895, 34.65796, 34.65623, 
    34.65405, 34.65156, 34.64751, 34.63829, 34.6203, 34.57959, 34.52196, 
    34.46996, 34.418, 34.33756, 34.21285, 34.06684, 33.95291, 33.97319,
  34.66393, 34.66395, 34.66399, 34.66469, 34.66592, 34.66661, 34.66607, 
    34.66492, 34.66432, 34.66448, 34.66496, 34.66516, 34.6647, 34.66355, 
    34.6628, 34.66277, 34.66226, 34.66071, 34.65907, 34.65854, 34.65904, 
    34.65966, 34.66009, 34.65997, 34.65869, 34.65707, 34.65647, 34.65664, 
    34.65683, 34.65689, 34.65679, 34.65618, 34.65485, 34.65327, 34.65228, 
    34.65228, 34.65283, 34.65321, 34.65307, 34.65253, 34.65065, 34.64738, 
    34.64325, 34.64004, 34.63638, 34.62791, 34.60469, 34.56413, 34.50814, 
    34.45712, 34.40476, 34.31823, 34.18109, 34.02483, 33.90691, 33.97319,
  34.65708, 34.65707, 34.65707, 34.6577, 34.65881, 34.65942, 34.65889, 
    34.65779, 34.65719, 34.6573, 34.65772, 34.65787, 34.65742, 34.65631, 
    34.6556, 34.65556, 34.65508, 34.65364, 34.65211, 34.65162, 34.6521, 
    34.65269, 34.6531, 34.65302, 34.65184, 34.65036, 34.6496, 34.64983, 
    34.65008, 34.65012, 34.64986, 34.64867, 34.64617, 34.6432, 34.64127, 
    34.64112, 34.64201, 34.64257, 34.64219, 34.64113, 34.6394, 34.63642, 
    34.63264, 34.62973, 34.62641, 34.61605, 34.59073, 34.5486, 34.49523, 
    34.44334, 34.38086, 34.28752, 34.14951, 33.98718, 33.86566, 33.97319,
  34.65079, 34.65075, 34.65072, 34.65128, 34.65229, 34.65283, 34.6523, 
    34.65125, 34.65066, 34.65071, 34.65107, 34.65119, 34.65074, 34.64968, 
    34.64889, 34.64878, 34.64791, 34.64539, 34.64271, 34.64181, 34.64256, 
    34.64351, 34.64416, 34.64394, 34.6418, 34.6391, 34.63807, 34.6383, 
    34.63854, 34.63859, 34.63837, 34.63729, 34.63499, 34.63226, 34.63049, 
    34.6304, 34.63126, 34.63184, 34.63156, 34.63063, 34.62907, 34.62635, 
    34.6229, 34.61943, 34.61401, 34.60144, 34.57791, 34.53434, 34.48338, 
    34.43068, 34.35891, 34.25105, 34.10357, 33.94864, 33.82772, 33.97319,
  34.64055, 34.64048, 34.64042, 34.64135, 34.64304, 34.64394, 34.64302, 
    34.64119, 34.64019, 34.64038, 34.64098, 34.64116, 34.64039, 34.63863, 
    34.63743, 34.63729, 34.63644, 34.63406, 34.63153, 34.63068, 34.63136, 
    34.63224, 34.63283, 34.63261, 34.63062, 34.6281, 34.62715, 34.62738, 
    34.62761, 34.62768, 34.62749, 34.62651, 34.6244, 34.6219, 34.62029, 
    34.62024, 34.62109, 34.62169, 34.62148, 34.62068, 34.6185, 34.61409, 
    34.60848, 34.60414, 34.59919, 34.58761, 34.5627, 34.52084, 34.47216, 
    34.4187, 34.33813, 34.2165, 34.06004, 33.90525, 33.79176, 33.97319,
  34.62986, 34.62975, 34.62966, 34.63047, 34.632, 34.63278, 34.63187, 
    34.63012, 34.62914, 34.62923, 34.62973, 34.62984, 34.62907, 34.62737, 
    34.62621, 34.62603, 34.62521, 34.62297, 34.62059, 34.61977, 34.62039, 
    34.62119, 34.62172, 34.62151, 34.61967, 34.61733, 34.61617, 34.61644, 
    34.61671, 34.61673, 34.61634, 34.61477, 34.61145, 34.6075, 34.60489, 
    34.60465, 34.6058, 34.60654, 34.60605, 34.60465, 34.6023, 34.59824, 
    34.5931, 34.58915, 34.58466, 34.57405, 34.54637, 34.50666, 34.46011, 
    34.40696, 34.31775, 34.18263, 34.01736, 33.86271, 33.75369, 33.97319,
  34.61873, 34.6186, 34.61847, 34.61946, 34.62083, 34.62149, 34.62059, 
    34.61892, 34.61784, 34.61795, 34.61835, 34.61839, 34.61761, 34.61538, 
    34.61363, 34.61335, 34.61209, 34.60868, 34.60508, 34.60384, 34.60476, 
    34.60594, 34.6067, 34.60635, 34.60353, 34.59998, 34.59859, 34.59884, 
    34.59909, 34.59909, 34.59874, 34.59728, 34.59423, 34.5906, 34.58818, 
    34.58796, 34.58902, 34.58971, 34.58929, 34.58805, 34.58591, 34.58221, 
    34.57753, 34.57398, 34.56896, 34.55549, 34.52985, 34.49169, 34.4435, 
    34.3798, 34.28461, 34.14837, 33.97419, 33.81967, 33.71222, 33.97319,
  34.59831, 34.59826, 34.59822, 34.59952, 34.60187, 34.60307, 34.60176, 
    34.59923, 34.59789, 34.59814, 34.59888, 34.59906, 34.59797, 34.59564, 
    34.59404, 34.59378, 34.59263, 34.58952, 34.58624, 34.58512, 34.58597, 
    34.58705, 34.58775, 34.58743, 34.58487, 34.58163, 34.58038, 34.58061, 
    34.58083, 34.58083, 34.58049, 34.57917, 34.57639, 34.57308, 34.57087, 
    34.57066, 34.57163, 34.57228, 34.57194, 34.57086, 34.56827, 34.56367, 
    34.55784, 34.55336, 34.54825, 34.53604, 34.51244, 34.47619, 34.4263, 
    34.35015, 34.23588, 34.0865, 33.9193, 33.77405, 33.66929, 33.97319,
  34.57694, 34.57699, 34.57702, 34.57825, 34.58044, 34.58158, 34.58042, 
    34.5782, 34.57701, 34.57725, 34.57791, 34.57806, 34.57707, 34.57498, 
    34.57354, 34.5733, 34.57227, 34.56948, 34.56614, 34.56465, 34.5658, 
    34.56723, 34.56792, 34.56763, 34.56438, 34.56027, 34.5587, 34.55901, 
    34.5593, 34.5593, 34.55886, 34.55723, 34.55382, 34.54976, 34.54707, 
    34.54679, 34.5479, 34.54863, 34.54815, 34.54677, 34.54437, 34.54027, 
    34.53507, 34.53111, 34.52658, 34.51568, 34.49222, 34.45895, 34.40831, 
    34.31914, 34.1849, 34.02174, 33.85744, 33.71812, 33.62437, 33.97319,
  34.54314, 34.54359, 34.54402, 34.54631, 34.55004, 34.55208, 34.55063, 
    34.54759, 34.54622, 34.547, 34.5483, 34.54882, 34.54771, 34.54512, 
    34.54345, 34.54339, 34.54229, 34.53882, 34.53519, 34.53422, 34.53555, 
    34.53712, 34.5382, 34.53808, 34.53542, 34.53205, 34.53089, 34.53135, 
    34.5318, 34.53196, 34.5317, 34.53038, 34.52747, 34.52396, 34.52165, 
    34.52146, 34.52247, 34.52314, 34.52277, 34.5216, 34.5195, 34.51592, 
    34.51115, 34.50707, 34.50253, 34.49169, 34.47118, 34.43338, 34.37047, 
    34.26778, 34.12487, 33.9544, 33.79312, 33.65998, 33.57653, 33.97319,
  34.5018, 34.50283, 34.50381, 34.50638, 34.51023, 34.51255, 34.51182, 
    34.50974, 34.50906, 34.51022, 34.51178, 34.51265, 34.5121, 34.5103, 
    34.50926, 34.50959, 34.50906, 34.50645, 34.50366, 34.50321, 34.50473, 
    34.50644, 34.5077, 34.50791, 34.50592, 34.50165, 34.50031, 34.50109, 
    34.50186, 34.50223, 34.50207, 34.50063, 34.49733, 34.4934, 34.49104, 
    34.49111, 34.4925, 34.49348, 34.49329, 34.49228, 34.49031, 34.48686, 
    34.48251, 34.47944, 34.47598, 34.46707, 34.44386, 34.40732, 34.32453, 
    34.19328, 34.031, 33.86501, 33.71645, 33.5997, 33.5278, 33.97319,
  34.43709, 34.43912, 34.44115, 34.44579, 34.45237, 34.45657, 34.45596, 
    34.45317, 34.45273, 34.45524, 34.45834, 34.46035, 34.46017, 34.45816, 
    34.45731, 34.45853, 34.45845, 34.45541, 34.45224, 34.45245, 34.45544, 
    34.45863, 34.46123, 34.46235, 34.46051, 34.458, 34.45797, 34.45964, 
    34.46133, 34.46259, 34.46333, 34.46296, 34.46093, 34.4583, 34.45702, 
    34.45774, 34.45952, 34.46093, 34.46133, 34.46099, 34.45987, 34.45745, 
    34.45356, 34.44948, 34.44496, 34.43338, 34.41131, 34.35573, 34.25775, 
    34.1097, 33.93783, 33.77517, 33.63691, 33.53913, 33.50425, 33.97319,
  34.36266, 34.36588, 34.36913, 34.37455, 34.38155, 34.38658, 34.38764, 
    34.38689, 34.38803, 34.3916, 34.39565, 34.39878, 34.40008, 34.39988, 
    34.40063, 34.40307, 34.40332, 34.3985, 34.39352, 34.39397, 34.39902, 
    34.40444, 34.40892, 34.41096, 34.4082, 34.40444, 34.40474, 34.4078, 
    34.41092, 34.41338, 34.41501, 34.41491, 34.4123, 34.40887, 34.40767, 
    34.4095, 34.41287, 34.41555, 34.41673, 34.41684, 34.41606, 34.41354, 
    34.41005, 34.40801, 34.4056, 34.39734, 34.35727, 34.29716, 34.16117, 
    33.98938, 33.82123, 33.67222, 33.55999, 33.50066, 33.49156, 33.97319,
  34.24461, 34.24866, 34.2529, 34.26057, 34.27051, 34.27781, 34.27932, 
    34.27787, 34.27944, 34.28492, 34.29123, 34.29622, 34.29842, 34.29812, 
    34.29944, 34.30355, 34.30587, 34.30441, 34.30292, 34.30581, 34.3125, 
    34.31957, 34.32593, 34.33031, 34.33078, 34.33053, 34.33344, 34.33848, 
    34.34363, 34.34812, 34.35182, 34.35403, 34.35407, 34.3533, 34.35102, 
    34.35398, 34.35978, 34.36426, 34.36595, 34.36564, 34.36377, 34.35854, 
    34.35133, 34.3465, 34.34081, 34.32372, 34.29003, 34.1866, 34.03656, 
    33.86312, 33.70612, 33.57545, 33.49996, 33.48138, 33.51398, 33.97319,
  34.1222, 34.12582, 34.12982, 34.13791, 34.14881, 34.15699, 34.15846, 
    34.15611, 34.15749, 34.16393, 34.1715, 34.17754, 34.18002, 34.17901, 
    34.18016, 34.18521, 34.18769, 34.18478, 34.18172, 34.18492, 34.19391, 
    34.2037, 34.21246, 34.21837, 34.21831, 34.21685, 34.22052, 34.22783, 
    34.23524, 34.24176, 34.24714, 34.25002, 34.24925, 34.24711, 34.2482, 
    34.25355, 34.26112, 34.26734, 34.27124, 34.27347, 34.27484, 34.27346, 
    34.27043, 34.26889, 34.25842, 34.22738, 34.16679, 34.05983, 33.90025, 
    33.73526, 33.58892, 33.49141, 33.47034, 33.49822, 33.5295, 33.97319,
  34.00139, 34.00306, 34.00526, 34.01066, 34.01855, 34.02489, 34.02625, 
    34.0244, 34.02556, 34.03128, 34.03807, 34.04379, 34.0463, 34.04525, 
    34.04627, 34.05133, 34.05373, 34.05023, 34.04633, 34.04934, 34.05924, 
    34.07046, 34.08034, 34.08714, 34.08677, 34.08404, 34.0879, 34.09679, 
    34.10546, 34.1131, 34.11933, 34.12233, 34.12013, 34.11581, 34.11552, 
    34.12159, 34.13125, 34.13924, 34.14376, 34.14572, 34.14597, 34.14172, 
    34.13463, 34.12976, 34.12358, 34.1019, 34.02359, 33.91216, 33.7518, 
    33.59795, 33.48885, 33.46653, 33.48154, 33.51027, 33.53548, 33.97319,
  33.92289, 33.91921, 33.91602, 33.91533, 33.91732, 33.91802, 33.91477, 
    33.90956, 33.90701, 33.90825, 33.90987, 33.91114, 33.9104, 33.9073, 
    33.90609, 33.90829, 33.90886, 33.90522, 33.90158, 33.9038, 33.9119, 
    33.92161, 33.92966, 33.93613, 33.93788, 33.93532, 33.93893, 33.94813, 
    33.95636, 33.96366, 33.96955, 33.9725, 33.96947, 33.96388, 33.96176, 
    33.96727, 33.97745, 33.98648, 33.99151, 33.99359, 33.99277, 33.9864, 
    33.97646, 33.96971, 33.96111, 33.93244, 33.86426, 33.74912, 33.60287, 
    33.48509, 33.45364, 33.46853, 33.49271, 33.51839, 33.53928, 33.97319,
  33.92331, 33.91288, 33.90282, 33.89315, 33.88619, 33.87867, 33.86981, 
    33.86208, 33.85489, 33.84892, 33.84181, 33.83518, 33.82803, 33.82041, 
    33.81354, 33.80855, 33.80327, 33.79498, 33.78632, 33.7826, 33.78435, 
    33.78839, 33.79018, 33.79182, 33.79013, 33.78453, 33.78537, 33.79181, 
    33.79582, 33.79943, 33.80227, 33.80487, 33.80322, 33.7989, 33.79428, 
    33.79725, 33.80545, 33.81454, 33.82005, 33.82303, 33.82101, 33.81334, 
    33.80224, 33.79631, 33.78868, 33.76059, 33.70129, 33.58842, 33.47945, 
    33.44241, 33.46198, 33.47801, 33.50238, 33.52171, 33.53947, 33.97319,
  33.99631, 33.97913, 33.96267, 33.94501, 33.93001, 33.9149, 33.90115, 
    33.89241, 33.88158, 33.86848, 33.85217, 33.83658, 33.82188, 33.80993, 
    33.7963, 33.78115, 33.7682, 33.75423, 33.73883, 33.72612, 33.71671, 
    33.70987, 33.70042, 33.69322, 33.68585, 33.67389, 33.66778, 33.66744, 
    33.66365, 33.6599, 33.65582, 33.6537, 33.64798, 33.64076, 33.63075, 
    33.62723, 33.62843, 33.63466, 33.64004, 33.64535, 33.64224, 33.63332, 
    33.62143, 33.61801, 33.61339, 33.58936, 33.53117, 33.45555, 33.4329, 
    33.4538, 33.47751, 33.48825, 33.506, 33.52185, 33.53962, 33.97319,
  34.13303, 34.10936, 34.08702, 34.06275, 34.04167, 34.0208, 34.00304, 
    33.99345, 33.9797, 33.96109, 33.93744, 33.91397, 33.8918, 33.8751, 
    33.85414, 33.82825, 33.8066, 33.78524, 33.76139, 33.73783, 33.71483, 
    33.69398, 33.67076, 33.65175, 33.63568, 33.61578, 33.60017, 33.58947, 
    33.57585, 33.56281, 33.55005, 33.54064, 33.52884, 33.51586, 33.49691, 
    33.48286, 33.47266, 33.4718, 33.47265, 33.47574, 33.46435, 33.45303, 
    33.44404, 33.44746, 33.45132, 33.4433, 33.4049, 33.41793, 33.44546, 
    33.47193, 33.48176, 33.49222, 33.50611, 33.52192, 33.53958, 33.97319,
  34.32937, 34.29786, 34.26839, 34.23699, 34.21014, 34.18361, 34.16081, 
    34.14817, 34.12993, 34.10535, 34.07455, 34.04388, 34.01457, 33.99113, 
    33.96244, 33.92774, 33.89682, 33.86663, 33.83408, 33.80007, 33.76511, 
    33.7316, 33.69677, 33.66637, 33.6403, 33.61281, 33.58747, 33.56509, 
    33.54217, 33.52052, 33.49998, 33.48263, 33.46526, 33.44825, 33.42371, 
    33.40165, 33.38173, 33.37339, 33.36878, 33.368, 33.35246, 33.34753, 
    33.34904, 33.36243, 33.37877, 33.40004, 33.41382, 33.43714, 33.46096, 
    33.47292, 33.48331, 33.49232, 33.50616, 33.52186, 33.53954, 33.97319,
  34.45667, 34.42141, 34.38903, 34.35859, 34.33643, 34.31074, 34.28281, 
    34.26471, 34.2428, 34.21651, 34.18394, 34.15014, 34.11579, 34.08504, 
    34.05039, 34.01142, 33.97348, 33.93622, 33.8983, 33.8592, 33.82027, 
    33.78283, 33.74577, 33.71166, 33.68124, 33.65199, 33.62212, 33.59204, 
    33.56408, 33.53868, 33.51587, 33.49524, 33.47846, 33.4658, 33.44594, 
    33.4268, 33.4089, 33.40184, 33.39893, 33.39991, 33.38961, 33.38437, 
    33.38386, 33.39354, 33.40626, 33.42435, 33.43756, 33.44928, 33.46191, 
    33.47332, 33.48345, 33.49237, 33.50613, 33.52182, 33.53951, 33.97319,
  34.47111, 34.43566, 34.40356, 34.37484, 34.35606, 34.33239, 34.3038, 
    34.28457, 34.26215, 34.23658, 34.20539, 34.17199, 34.13635, 34.10255, 
    34.06575, 34.02598, 33.98621, 33.94601, 33.90543, 33.86522, 33.82669, 
    33.78978, 33.75347, 33.72001, 33.68948, 33.66022, 33.63305, 33.60784, 
    33.5845, 33.56307, 33.54363, 33.52639, 33.51251, 33.50072, 33.48059, 
    33.46048, 33.44046, 33.43207, 33.42711, 33.42559, 33.41172, 33.40271, 
    33.39856, 33.40741, 33.4195, 33.43485, 33.44065, 33.44983, 33.46224, 
    33.47348, 33.48349, 33.49239, 33.50611, 33.52179, 33.53948, 33.97319,
  34.47064, 34.43496, 34.40276, 34.37405, 34.35544, 34.3318, 34.30314, 
    34.28392, 34.26149, 34.23585, 34.20448, 34.17099, 34.13538, 34.10153, 
    34.0647, 34.02488, 33.98521, 33.94516, 33.90474, 33.86455, 33.82573, 
    33.7883, 33.75201, 33.71843, 33.68751, 33.65844, 33.63291, 33.6109, 
    33.58891, 33.5684, 33.54938, 33.53175, 33.5169, 33.50482, 33.48481, 
    33.46415, 33.44286, 33.43291, 33.42722, 33.4258, 33.41172, 33.40264, 
    33.39852, 33.40747, 33.41964, 33.43504, 33.44085, 33.44994, 33.46249, 
    33.47359, 33.48349, 33.4924, 33.5061, 33.52179, 33.53948, 33.97319,
  34.46987, 34.43404, 34.40176, 34.37301, 34.35455, 34.33101, 34.30237, 
    34.28321, 34.26083, 34.23521, 34.20386, 34.17039, 34.1348, 34.10104, 
    34.06417, 34.02419, 33.98443, 33.94432, 33.90387, 33.86362, 33.82472, 
    33.78714, 33.75091, 33.71723, 33.6861, 33.65716, 33.63224, 33.61132, 
    33.59, 33.57009, 33.55159, 33.53442, 33.51995, 33.50821, 33.48844, 
    33.46795, 33.44672, 33.43631, 33.43013, 33.42816, 33.41314, 33.40355, 
    33.39935, 33.40807, 33.42008, 33.43544, 33.44119, 33.4503, 33.46286, 
    33.47368, 33.4835, 33.49241, 33.5061, 33.52179, 33.53948, 33.97319,
  34.46923, 34.43326, 34.40086, 34.37204, 34.35368, 34.33012, 34.30134, 
    34.28218, 34.25978, 34.23413, 34.20279, 34.1693, 34.13369, 34.09998, 
    34.06318, 34.02328, 33.98355, 33.94351, 33.90318, 33.86298, 33.8241, 
    33.78655, 33.75038, 33.71678, 33.68576, 33.65692, 33.63223, 33.61166, 
    33.59059, 33.57099, 33.55287, 33.53609, 33.52189, 33.51025, 33.49059, 
    33.47031, 33.44942, 33.43913, 33.43293, 33.43082, 33.41588, 33.40614, 
    33.4016, 33.40976, 33.42135, 33.43636, 33.44168, 33.45056, 33.46299, 
    33.47369, 33.4835, 33.49241, 33.5061, 33.52179, 33.53948, 33.97319,
  34.68758, 34.6876, 34.68762, 34.68786, 34.68828, 34.68855, 34.68845, 
    34.68812, 34.68797, 34.68808, 34.6883, 34.68841, 34.68827, 34.68792, 
    34.68769, 34.68771, 34.68755, 34.687, 34.68636, 34.68615, 34.68633, 
    34.68653, 34.68666, 34.68657, 34.68599, 34.68523, 34.68489, 34.68486, 
    34.68484, 34.68476, 34.68461, 34.68422, 34.68345, 34.68256, 34.68196, 
    34.68185, 34.68202, 34.6821, 34.68192, 34.68155, 34.68098, 34.68008, 
    34.67894, 34.67786, 34.67631, 34.67289, 34.66336, 34.63921, 34.59017, 
    34.52825, 34.47561, 34.42394, 34.34577, 34.23838, 34.15038, 33.96647,
  34.6845, 34.68452, 34.68456, 34.68488, 34.68528, 34.68552, 34.68539, 
    34.6851, 34.68488, 34.68495, 34.6851, 34.68516, 34.68501, 34.68448, 
    34.6841, 34.68407, 34.6838, 34.68302, 34.68219, 34.68192, 34.68212, 
    34.68236, 34.6825, 34.68239, 34.68174, 34.68093, 34.68059, 34.68059, 
    34.6806, 34.68055, 34.68042, 34.68007, 34.67939, 34.6786, 34.67783, 
    34.6777, 34.67797, 34.67812, 34.67787, 34.67734, 34.67656, 34.67532, 
    34.67377, 34.67254, 34.67117, 34.66639, 34.65493, 34.62595, 34.5729, 
    34.51078, 34.46076, 34.40929, 34.32071, 34.19622, 34.09034, 33.96647,
  34.67998, 34.68002, 34.68007, 34.68044, 34.68107, 34.68142, 34.68119, 
    34.68071, 34.68045, 34.68052, 34.68075, 34.68084, 34.68064, 34.68011, 
    34.67978, 34.67977, 34.67954, 34.67885, 34.67795, 34.67757, 34.67789, 
    34.67828, 34.67851, 34.6784, 34.67746, 34.6763, 34.67583, 34.67588, 
    34.67593, 34.67591, 34.67577, 34.67528, 34.67432, 34.67319, 34.67246, 
    34.67239, 34.6727, 34.67288, 34.6727, 34.67225, 34.67159, 34.67048, 
    34.66851, 34.66634, 34.66387, 34.6582, 34.64275, 34.60958, 34.5531, 
    34.49476, 34.4435, 34.38139, 34.28511, 34.16015, 34.03893, 33.96647,
  34.67511, 34.67516, 34.67521, 34.67573, 34.6766, 34.6771, 34.67675, 
    34.67603, 34.67565, 34.67577, 34.67611, 34.67624, 34.67595, 34.6752, 
    34.67472, 34.67471, 34.67438, 34.67337, 34.6723, 34.67197, 34.67229, 
    34.67268, 34.67294, 34.67285, 34.67202, 34.67099, 34.67059, 34.67068, 
    34.67078, 34.6708, 34.67071, 34.67031, 34.66946, 34.66788, 34.66661, 
    34.66648, 34.66702, 34.66733, 34.66703, 34.66627, 34.66511, 34.66316, 
    34.66069, 34.65872, 34.65644, 34.64952, 34.63068, 34.59307, 34.53609, 
    34.48098, 34.42865, 34.35553, 34.24336, 34.11045, 33.99467, 33.96647,
  34.66994, 34.66999, 34.67004, 34.67052, 34.67133, 34.67179, 34.67147, 
    34.67079, 34.67044, 34.67054, 34.67085, 34.67098, 34.67072, 34.67002, 
    34.66958, 34.66959, 34.66929, 34.66837, 34.66689, 34.66632, 34.66684, 
    34.66748, 34.66792, 34.66777, 34.66635, 34.66457, 34.66389, 34.66403, 
    34.66418, 34.6642, 34.66404, 34.66333, 34.66184, 34.66008, 34.65896, 
    34.65891, 34.65946, 34.65982, 34.6596, 34.65894, 34.65792, 34.65616, 
    34.65392, 34.65132, 34.64711, 34.63759, 34.61929, 34.57877, 34.52134, 
    34.46904, 34.41578, 34.3331, 34.20712, 34.06381, 33.95432, 33.96647,
  34.66392, 34.66395, 34.66399, 34.6647, 34.66594, 34.66663, 34.66609, 
    34.66493, 34.66434, 34.66454, 34.66502, 34.66522, 34.66476, 34.66363, 
    34.66289, 34.66286, 34.66233, 34.66077, 34.65911, 34.65858, 34.65907, 
    34.65969, 34.66011, 34.65999, 34.65869, 34.65706, 34.65646, 34.65662, 
    34.6568, 34.65686, 34.65675, 34.65614, 34.65481, 34.65323, 34.65225, 
    34.65225, 34.65283, 34.65322, 34.65307, 34.6525, 34.6506, 34.6473, 
    34.64311, 34.63977, 34.63591, 34.62712, 34.6038, 34.56342, 34.50752, 
    34.45604, 34.40228, 34.31338, 34.17525, 34.02277, 33.90891, 33.96647,
  34.65704, 34.65704, 34.65705, 34.65768, 34.65881, 34.65942, 34.65889, 
    34.65778, 34.65719, 34.65734, 34.65776, 34.65792, 34.65748, 34.6564, 
    34.65569, 34.65565, 34.65515, 34.65369, 34.65215, 34.65166, 34.65213, 
    34.65271, 34.65312, 34.65302, 34.65184, 34.65034, 34.64957, 34.6498, 
    34.65004, 34.65007, 34.6498, 34.64862, 34.64612, 34.64315, 34.64122, 
    34.64109, 34.642, 34.64257, 34.64219, 34.64109, 34.63934, 34.63633, 
    34.63248, 34.62943, 34.62589, 34.61526, 34.58994, 34.54802, 34.49458, 
    34.44199, 34.37799, 34.28244, 34.14375, 33.98598, 33.86819, 33.96647,
  34.65073, 34.6507, 34.65068, 34.65125, 34.65226, 34.65281, 34.65228, 
    34.65121, 34.65063, 34.65073, 34.6511, 34.65123, 34.6508, 34.64976, 
    34.64898, 34.64888, 34.64798, 34.64545, 34.64277, 34.64186, 34.6426, 
    34.64354, 34.64418, 34.64394, 34.6418, 34.63908, 34.63804, 34.63826, 
    34.63848, 34.63853, 34.6383, 34.63721, 34.63492, 34.63219, 34.63043, 
    34.63035, 34.63125, 34.63184, 34.63155, 34.63058, 34.62901, 34.62626, 
    34.62273, 34.61912, 34.61351, 34.60077, 34.57722, 34.53389, 34.48269, 
    34.42909, 34.3557, 34.24582, 34.09872, 33.94818, 33.83074, 33.96647,
  34.64046, 34.6404, 34.64035, 34.64129, 34.64299, 34.64388, 34.64296, 
    34.64112, 34.64015, 34.64038, 34.641, 34.64119, 34.64044, 34.63871, 
    34.63754, 34.63739, 34.63652, 34.63413, 34.63161, 34.63074, 34.63142, 
    34.63229, 34.63286, 34.63263, 34.63063, 34.62809, 34.62712, 34.62734, 
    34.62755, 34.62761, 34.6274, 34.62642, 34.62432, 34.62182, 34.62022, 
    34.62019, 34.62107, 34.62169, 34.62147, 34.62063, 34.61844, 34.61401, 
    34.60835, 34.60389, 34.59877, 34.58704, 34.56216, 34.52051, 34.47144, 
    34.41687, 34.33458, 34.21112, 34.05606, 33.90536, 33.79524, 33.96647,
  34.62974, 34.62965, 34.62956, 34.63038, 34.63191, 34.63269, 34.63178, 
    34.63002, 34.62906, 34.62922, 34.62973, 34.62986, 34.62911, 34.62745, 
    34.62632, 34.62614, 34.6253, 34.62305, 34.62068, 34.61985, 34.62046, 
    34.62125, 34.62177, 34.62154, 34.61969, 34.61732, 34.61615, 34.6164, 
    34.61665, 34.61664, 34.61625, 34.61467, 34.61136, 34.60742, 34.60482, 
    34.6046, 34.60579, 34.60654, 34.60604, 34.60462, 34.60227, 34.5982, 
    34.59301, 34.58896, 34.58433, 34.57359, 34.54599, 34.50638, 34.45929, 
    34.4049, 34.31388, 34.17712, 34.01425, 33.86338, 33.75711, 33.96647,
  34.61858, 34.61845, 34.61834, 34.61934, 34.6207, 34.62137, 34.62047, 
    34.61879, 34.61774, 34.61793, 34.61833, 34.61839, 34.61765, 34.61546, 
    34.61375, 34.61348, 34.61219, 34.60878, 34.60519, 34.60395, 34.60486, 
    34.60603, 34.60678, 34.6064, 34.60357, 34.60001, 34.5986, 34.59883, 
    34.59905, 34.59903, 34.59866, 34.5972, 34.59415, 34.59053, 34.58812, 
    34.58792, 34.58901, 34.58973, 34.58931, 34.58804, 34.58591, 34.58221, 
    34.57749, 34.57385, 34.56872, 34.55519, 34.52964, 34.49141, 34.44236, 
    34.37735, 34.28053, 34.14272, 33.97194, 33.82091, 33.71504, 33.96647,
  34.59812, 34.59809, 34.59805, 34.59936, 34.60171, 34.60291, 34.6016, 
    34.59906, 34.59776, 34.5981, 34.59885, 34.59905, 34.598, 34.59572, 
    34.59416, 34.59391, 34.59275, 34.58965, 34.58638, 34.58526, 34.58611, 
    34.58718, 34.58787, 34.58753, 34.58496, 34.5817, 34.58042, 34.58062, 
    34.58081, 34.58079, 34.58044, 34.5791, 34.57632, 34.57302, 34.57082, 
    34.57063, 34.57163, 34.5723, 34.57197, 34.57087, 34.56831, 34.56371, 
    34.55785, 34.55333, 34.54815, 34.5359, 34.51237, 34.47591, 34.42482, 
    34.34729, 34.23173, 34.08178, 33.91771, 33.77574, 33.67149, 33.96647,
  34.57671, 34.57677, 34.57682, 34.57806, 34.58025, 34.58138, 34.58023, 
    34.57799, 34.57685, 34.57719, 34.57787, 34.57804, 34.57709, 34.57507, 
    34.57367, 34.57344, 34.57241, 34.56963, 34.56631, 34.56483, 34.56598, 
    34.5674, 34.56808, 34.56778, 34.56451, 34.56038, 34.55878, 34.55906, 
    34.55931, 34.55928, 34.55883, 34.55717, 34.55376, 34.54971, 34.54702, 
    34.54676, 34.5479, 34.54865, 34.54818, 34.54681, 34.54444, 34.54034, 
    34.53514, 34.53117, 34.52662, 34.51573, 34.49216, 34.45862, 34.40646, 
    34.31583, 34.18068, 34.01801, 33.85645, 33.71918, 33.62599, 33.96647,
  34.54284, 34.54331, 34.54375, 34.54605, 34.54977, 34.55181, 34.55036, 
    34.54731, 34.54598, 34.54688, 34.5482, 34.54876, 34.54768, 34.54516, 
    34.54353, 34.5435, 34.5424, 34.53895, 34.53534, 34.53439, 34.53573, 
    34.5373, 34.53838, 34.53826, 34.53558, 34.53219, 34.53101, 34.53143, 
    34.53185, 34.53197, 34.53168, 34.53034, 34.52742, 34.52391, 34.5216, 
    34.52142, 34.52245, 34.52316, 34.52281, 34.52167, 34.5196, 34.51604, 
    34.51128, 34.50719, 34.50262, 34.4917, 34.47113, 34.4327, 34.36805, 
    34.26421, 34.12081, 33.9517, 33.79275, 33.66039, 33.57925, 33.96647,
  34.50141, 34.50246, 34.50345, 34.50603, 34.50986, 34.51218, 34.51144, 
    34.50935, 34.50873, 34.51, 34.5116, 34.5125, 34.51199, 34.51027, 
    34.50928, 34.50964, 34.50912, 34.50654, 34.5038, 34.50337, 34.50491, 
    34.50663, 34.50791, 34.50812, 34.5061, 34.5018, 34.50043, 34.50117, 
    34.5019, 34.50224, 34.50204, 34.50056, 34.49722, 34.49326, 34.49085, 
    34.49092, 34.49234, 34.49336, 34.4932, 34.49221, 34.49028, 34.48683, 
    34.48248, 34.47946, 34.476, 34.46704, 34.44362, 34.4063, 34.32145, 
    34.18965, 34.02824, 33.86258, 33.7156, 33.60035, 33.53165, 33.96647,
  34.43657, 34.43862, 34.44065, 34.4453, 34.45185, 34.45604, 34.45541, 
    34.4526, 34.4522, 34.45483, 34.45795, 34.46, 34.45986, 34.4579, 34.4571, 
    34.45834, 34.45827, 34.45524, 34.45211, 34.45234, 34.45537, 34.45861, 
    34.46124, 34.46236, 34.4605, 34.45798, 34.45791, 34.45953, 34.46118, 
    34.46241, 34.4631, 34.46267, 34.46059, 34.45793, 34.4566, 34.4573, 
    34.45909, 34.46054, 34.46099, 34.46072, 34.45961, 34.45722, 34.45335, 
    34.44931, 34.44476, 34.43299, 34.4107, 34.35418, 34.25418, 34.1063, 
    33.93631, 33.77294, 33.6352, 33.54096, 33.51435, 33.96647,
  34.36198, 34.36522, 34.36847, 34.37389, 34.38084, 34.38584, 34.38687, 
    34.38608, 34.38726, 34.39093, 34.39499, 34.39815, 34.39948, 34.39933, 
    34.40012, 34.40259, 34.40285, 34.39803, 34.39307, 34.39356, 34.39867, 
    34.40414, 34.40869, 34.41074, 34.40794, 34.40416, 34.4044, 34.40738, 
    34.41046, 34.41287, 34.41443, 34.41421, 34.41148, 34.40794, 34.40662, 
    34.4084, 34.41177, 34.4145, 34.41574, 34.41594, 34.41515, 34.41263, 
    34.40915, 34.40725, 34.40488, 34.3965, 34.35618, 34.29504, 34.15742, 
    33.98733, 33.81947, 33.6689, 33.5601, 33.50854, 33.50694, 33.96647,
  34.24387, 34.24794, 34.25219, 34.25983, 34.26971, 34.27694, 34.27838, 
    34.27687, 34.27845, 34.284, 34.29027, 34.29523, 34.29742, 34.29714, 
    34.29847, 34.30259, 34.3049, 34.30344, 34.302, 34.30493, 34.31168, 
    34.31882, 34.32527, 34.32967, 34.3301, 34.32985, 34.33268, 34.33757, 
    34.34266, 34.34707, 34.35065, 34.35267, 34.35255, 34.35163, 34.34919, 
    34.35205, 34.35783, 34.36236, 34.36413, 34.36393, 34.36202, 34.35677, 
    34.34956, 34.34493, 34.33934, 34.32215, 34.28839, 34.18439, 34.03342, 
    33.86137, 33.70345, 33.57274, 33.50426, 33.49497, 33.52157, 33.96647,
  34.12169, 34.12535, 34.12936, 34.13741, 34.14822, 34.15628, 34.15764, 
    34.15523, 34.15659, 34.16304, 34.17046, 34.17638, 34.17876, 34.17773, 
    34.17884, 34.18385, 34.18629, 34.18338, 34.18037, 34.18362, 34.19271, 
    34.20264, 34.21154, 34.21751, 34.21746, 34.21608, 34.21965, 34.22671, 
    34.23401, 34.24035, 34.24549, 34.24801, 34.24693, 34.2445, 34.24529, 
    34.25043, 34.25788, 34.26411, 34.26809, 34.27047, 34.2718, 34.27045, 
    34.26752, 34.26635, 34.25613, 34.22525, 34.16505, 34.05779, 33.89782, 
    33.73278, 33.58419, 33.49384, 33.48254, 33.50681, 33.53043, 33.96647,
  34.00134, 34.00309, 34.00534, 34.01074, 34.01858, 34.02478, 34.02596, 
    34.02403, 34.02514, 34.03075, 34.03726, 34.04271, 34.04501, 34.04389, 
    34.0448, 34.04971, 34.05201, 34.04846, 34.04453, 34.04753, 34.05754, 
    34.06898, 34.07906, 34.08597, 34.08564, 34.08304, 34.08681, 34.09536, 
    34.1039, 34.11129, 34.11712, 34.11955, 34.11681, 34.11202, 34.11121, 
    34.11691, 34.12636, 34.13431, 34.13893, 34.14111, 34.14134, 34.1372, 
    34.13039, 34.12618, 34.12061, 34.09945, 34.02177, 33.91056, 33.74823, 
    33.59341, 33.49155, 33.47544, 33.49057, 33.51268, 33.53103, 33.96647,
  33.92232, 33.91882, 33.91587, 33.91551, 33.91769, 33.91853, 33.91541, 
    33.91038, 33.90794, 33.90919, 33.91058, 33.91148, 33.91025, 33.90696, 
    33.90536, 33.90698, 33.90719, 33.90319, 33.8992, 33.9012, 33.90929, 
    33.9192, 33.92743, 33.93407, 33.93599, 33.9337, 33.93725, 33.94608, 
    33.95428, 33.96131, 33.9667, 33.96889, 33.96519, 33.95898, 33.95618, 
    33.96112, 33.97083, 33.97971, 33.9848, 33.98714, 33.9862, 33.97992, 
    33.97038, 33.96458, 33.95699, 33.92938, 33.86185, 33.7456, 33.59838, 
    33.48812, 33.4655, 33.47618, 33.49596, 33.51412, 33.53145, 33.96647,
  33.9174, 33.90679, 33.897, 33.88823, 33.8819, 33.87525, 33.86741, 33.86026, 
    33.85374, 33.8485, 33.84222, 33.83596, 33.82877, 33.82148, 33.81437, 
    33.80852, 33.80301, 33.7941, 33.78427, 33.77998, 33.78134, 33.78519, 
    33.78645, 33.78793, 33.78641, 33.78115, 33.78209, 33.7884, 33.79292, 
    33.79668, 33.79933, 33.80116, 33.79869, 33.79361, 33.78841, 33.7906, 
    33.79781, 33.80636, 33.81173, 33.8149, 33.81242, 33.80468, 33.79385, 
    33.7889, 33.78246, 33.75561, 33.69661, 33.58419, 33.48298, 33.45445, 
    33.46765, 33.48036, 33.49789, 33.51477, 33.5316, 33.96647,
  33.98709, 33.96806, 33.9507, 33.93326, 33.91821, 33.90402, 33.89189, 
    33.88362, 33.87366, 33.86194, 33.84792, 33.83408, 33.82061, 33.80977, 
    33.79661, 33.78124, 33.76891, 33.75446, 33.73738, 33.72437, 33.71446, 
    33.70697, 33.69568, 33.6876, 33.6802, 33.66797, 33.66188, 33.6619, 
    33.65948, 33.65702, 33.65417, 33.65197, 33.64601, 33.63833, 33.62862, 
    33.62454, 33.62432, 33.62936, 33.63371, 33.63808, 33.63314, 33.62387, 
    33.61228, 33.60999, 33.60689, 33.58516, 33.52743, 33.46133, 33.44331, 
    33.45824, 33.47301, 33.48238, 33.49869, 33.51491, 33.53172, 33.96647,
  34.13664, 34.10793, 34.0822, 34.0558, 34.03195, 34.01048, 33.99446, 
    33.98539, 33.97216, 33.95407, 33.93303, 33.91215, 33.8926, 33.87753, 
    33.85769, 33.83239, 33.81218, 33.79066, 33.76471, 33.74128, 33.7176, 
    33.69546, 33.6682, 33.64697, 33.63044, 33.60865, 33.59243, 33.58255, 
    33.57074, 33.56035, 33.55111, 33.54305, 33.53254, 33.52083, 33.50525, 
    33.49283, 33.48251, 33.48071, 33.48001, 33.48082, 33.46707, 33.45413, 
    33.44497, 33.44922, 33.45478, 33.45143, 33.41817, 33.42957, 33.44821, 
    33.464, 33.47401, 33.48323, 33.49882, 33.51497, 33.53166, 33.96647,
  34.33096, 34.2934, 34.26087, 34.22988, 34.2023, 34.17693, 34.15723, 
    34.14608, 34.1295, 34.1064, 34.08059, 34.05431, 34.02912, 34.0078, 
    33.98063, 33.94659, 33.9173, 33.88637, 33.84993, 33.81546, 33.77903, 
    33.74345, 33.70168, 33.66747, 33.6408, 33.60975, 33.58334, 33.56258, 
    33.54174, 33.52426, 33.51001, 33.49609, 33.48252, 33.46962, 33.45286, 
    33.43583, 33.41823, 33.41027, 33.4048, 33.40184, 33.38436, 33.37521, 
    33.37086, 33.38128, 33.39574, 33.41639, 33.4267, 33.43579, 33.45326, 
    33.46443, 33.47448, 33.48334, 33.49887, 33.51492, 33.5316, 33.96647,
  34.41564, 34.37495, 34.3409, 34.31345, 34.29168, 34.26983, 34.24804, 
    34.23204, 34.21403, 34.1938, 34.1702, 34.14385, 34.11503, 34.08929, 
    34.05782, 34.02017, 33.98614, 33.9481, 33.90536, 33.86613, 33.82642, 
    33.78707, 33.74409, 33.70658, 33.67514, 33.64215, 33.61309, 33.58812, 
    33.56505, 33.54651, 33.53256, 33.5177, 33.50608, 33.49709, 33.48497, 
    33.46976, 33.4517, 33.44333, 33.43732, 33.43355, 33.41646, 33.40356, 
    33.39463, 33.40086, 33.41151, 33.4269, 33.42899, 33.43766, 33.45366, 
    33.46471, 33.47466, 33.48342, 33.49885, 33.51487, 33.53155, 33.96647,
  34.41077, 34.36985, 34.3359, 34.30904, 34.28764, 34.26645, 34.24535, 
    34.22935, 34.21235, 34.19439, 34.17234, 34.14724, 34.11905, 34.09358, 
    34.06188, 34.02401, 33.98876, 33.94822, 33.90246, 33.86212, 33.8226, 
    33.78366, 33.73899, 33.70115, 33.66998, 33.6367, 33.60977, 33.589, 
    33.56993, 33.55519, 33.54486, 33.53214, 33.52113, 33.5113, 33.49855, 
    33.48273, 33.46391, 33.45444, 33.44689, 33.44126, 33.42329, 33.40903, 
    33.3985, 33.40368, 33.41363, 33.42837, 33.42947, 33.43801, 33.45394, 
    33.46492, 33.47471, 33.48346, 33.49883, 33.51484, 33.53152, 33.96647,
  34.40595, 34.36478, 34.3307, 34.30378, 34.28304, 34.26193, 34.24045, 
    34.22444, 34.20735, 34.1892, 34.16724, 34.14221, 34.11409, 34.08798, 
    34.05547, 34.01661, 33.98077, 33.93974, 33.89365, 33.85366, 33.8144, 
    33.77574, 33.73103, 33.69306, 33.66173, 33.62917, 33.60453, 33.58775, 
    33.57099, 33.5577, 33.54788, 33.5363, 33.52523, 33.5146, 33.501, 
    33.48468, 33.46569, 33.45461, 33.44631, 33.44077, 33.42297, 33.40887, 
    33.39848, 33.40374, 33.41378, 33.42863, 33.42978, 33.4383, 33.45417, 
    33.46501, 33.47473, 33.48349, 33.49883, 33.51483, 33.53152, 33.96647,
  34.40304, 34.36176, 34.32753, 34.30039, 34.28017, 34.25915, 34.23732, 
    34.22137, 34.20416, 34.18571, 34.16368, 34.13847, 34.11008, 34.08351, 
    34.05073, 34.01176, 33.97617, 33.93542, 33.88956, 33.85009, 33.81114, 
    33.77266, 33.7284, 33.69083, 33.65995, 33.62767, 33.60322, 33.58659, 
    33.57014, 33.55742, 33.54842, 33.53738, 33.52686, 33.51686, 33.50356, 
    33.48754, 33.4688, 33.45741, 33.44872, 33.44272, 33.42362, 33.40898, 
    33.39876, 33.40405, 33.41412, 33.42906, 33.43018, 33.43861, 33.45441, 
    33.46507, 33.47475, 33.48351, 33.49883, 33.51483, 33.53152, 33.96647,
  34.40163, 34.35985, 34.32531, 34.29802, 34.27793, 34.257, 34.23523, 
    34.21933, 34.2021, 34.18353, 34.1615, 34.13625, 34.10775, 34.08103, 
    34.04812, 34.00902, 33.97327, 33.93246, 33.88661, 33.84736, 33.80859, 
    33.77028, 33.7263, 33.68911, 33.65872, 33.62661, 33.60237, 33.586, 
    33.56979, 33.55745, 33.54897, 33.53837, 33.52825, 33.51862, 33.50566, 
    33.48993, 33.47142, 33.4602, 33.45151, 33.44537, 33.42632, 33.41147, 
    33.40083, 33.40548, 33.41516, 33.42984, 33.43058, 33.4388, 33.45451, 
    33.46508, 33.47475, 33.48351, 33.49883, 33.51483, 33.53152, 33.96647 ;

 salt_north =
  34.66766, 34.66767, 34.66498, 34.66027, 34.65579, 34.65334, 34.65135, 
    34.64808, 34.64547, 34.64398, 34.64197, 34.63961, 34.63744, 34.63489, 
    34.63248, 34.63154, 34.63239, 34.63386, 34.63428, 34.63214, 34.62042, 
    34.59029, 34.51262, 34.38235, 34.2407, 34.09169, 33.93779, 33.73247, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  34.65937, 34.65938, 34.65688, 34.65101, 34.64376, 34.6405, 34.63872, 
    34.63579, 34.63336, 34.63184, 34.62988, 34.62586, 34.6222, 34.61801, 
    34.61412, 34.61265, 34.61403, 34.61639, 34.61708, 34.61375, 34.60153, 
    34.56193, 34.47499, 34.34499, 34.20676, 34.06353, 33.89657, 33.688, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  34.65049, 34.65052, 34.64629, 34.63909, 34.63248, 34.62915, 34.626, 
    34.62081, 34.61655, 34.61403, 34.61076, 34.60711, 34.60382, 34.60006, 
    34.59658, 34.5953, 34.59657, 34.59877, 34.59949, 34.59649, 34.58361, 
    34.53589, 34.44282, 34.31306, 34.17775, 34.03211, 33.86129, 33.64988, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  34.63929, 34.63932, 34.63545, 34.62785, 34.61617, 34.61093, 34.60807, 
    34.60334, 34.59949, 34.59724, 34.59431, 34.59101, 34.58802, 34.58311, 
    34.57707, 34.57483, 34.57705, 34.58087, 34.58207, 34.57678, 34.55712, 
    34.51268, 34.41517, 34.28338, 34.14768, 34.00284, 33.8309, 33.58384, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  34.62931, 34.62934, 34.62248, 34.61075, 34.59996, 34.59514, 34.59252, 
    34.5882, 34.58374, 34.57997, 34.57494, 34.56922, 34.56398, 34.55806, 
    34.55252, 34.5505, 34.55251, 34.55606, 34.55722, 34.55223, 34.53415, 
    34.48149, 34.38313, 34.25136, 34.12064, 33.97743, 33.80135, 33.52318, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  34.61296, 34.61299, 34.60662, 34.59573, 34.58572, 34.57784, 34.57334, 
    34.56587, 34.55983, 34.55636, 34.5517, 34.54639, 34.54151, 34.53606, 
    34.53097, 34.52913, 34.53097, 34.53427, 34.5354, 34.53068, 34.51398, 
    34.45409, 34.35352, 34.22323, 34.09687, 33.95509, 33.75928, 33.46969, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  34.59832, 34.59836, 34.59243, 34.57983, 34.56274, 34.5551, 34.55093, 
    34.54402, 34.53843, 34.53524, 34.53091, 34.52596, 34.5214, 34.51637, 
    34.5111, 34.50835, 34.51105, 34.51477, 34.51587, 34.51049, 34.48583, 
    34.42958, 34.32703, 34.19804, 34.07559, 33.92952, 33.72155, 33.42165, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  34.58464, 34.58468, 34.57455, 34.55724, 34.54134, 34.53423, 34.53038, 
    34.52397, 34.5188, 34.51585, 34.51171, 34.50443, 34.49772, 34.49028, 
    34.48333, 34.4808, 34.48332, 34.48777, 34.48922, 34.48285, 34.45977, 
    34.40551, 34.3027, 34.17492, 34.05365, 33.89853, 33.68686, 33.33775, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  34.56137, 34.5614, 34.55197, 34.53586, 34.52106, 34.51447, 34.51073, 
    34.50129, 34.49367, 34.48934, 34.48341, 34.4766, 34.47032, 34.46345, 
    34.45703, 34.45472, 34.45706, 34.46119, 34.46253, 34.45667, 34.43509, 
    34.37562, 34.27567, 34.14901, 34.02743, 33.86917, 33.65397, 33.24246, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  34.53857, 34.53859, 34.52985, 34.5149, 34.49573, 34.48612, 34.48087, 
    34.47215, 34.46513, 34.46117, 34.45566, 34.44933, 34.44347, 34.43716, 
    34.43126, 34.42916, 34.43132, 34.43515, 34.43639, 34.43102, 34.4109, 
    34.34634, 34.24525, 34.1223, 34.00174, 33.8404, 33.60387, 33.14901, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  34.51549, 34.51552, 34.50559, 34.48406, 34.4643, 34.45547, 34.45064, 
    34.44267, 34.43626, 34.43266, 34.42759, 34.42174, 34.41631, 34.41056, 
    34.40323, 34.40049, 34.40327, 34.40814, 34.40964, 34.40278, 34.37654, 
    34.3167, 34.21448, 34.09527, 33.97574, 33.81128, 33.53454, 33.05449, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  34.48081, 34.48082, 34.46933, 34.44971, 34.43174, 34.42372, 34.41933, 
    34.41212, 34.40524, 34.40064, 34.39417, 34.38674, 34.37986, 34.37255, 
    34.3657, 34.36328, 34.36578, 34.37017, 34.3715, 34.36511, 34.34093, 
    34.28397, 34.1826, 34.06727, 33.94867, 33.75841, 33.46277, 32.91685, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  34.44171, 34.44172, 34.43139, 34.41376, 34.39347, 34.38335, 34.3778, 
    34.36872, 34.36147, 34.35749, 34.35173, 34.34508, 34.3389, 34.33247, 
    34.32644, 34.32435, 34.32655, 34.33045, 34.33159, 34.32568, 34.30366, 
    34.24081, 34.14454, 34.02956, 33.89999, 33.70089, 33.38317, 32.75711, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  34.39823, 34.39825, 34.38541, 34.36353, 34.34365, 34.33485, 34.33002, 
    34.32217, 34.31594, 34.3126, 34.30757, 34.30173, 34.29629, 34.28999, 
    34.28304, 34.28062, 34.28313, 34.28758, 34.28881, 34.28181, 34.25571, 
    34.19592, 34.10133, 33.98557, 33.84937, 33.64108, 33.18533, 32.59117, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  34.33959, 34.3397, 34.32869, 34.30987, 34.29289, 34.28379, 34.27827, 
    34.26935, 34.26235, 34.25869, 34.25312, 34.24662, 34.24053, 34.23444, 
    34.22867, 34.22673, 34.22876, 34.23246, 34.23337, 34.22684, 34.20332, 
    34.1451, 34.05731, 33.94057, 33.78552, 33.52402, 32.9838, 32.38899, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  34.2792, 34.27943, 34.26698, 34.24574, 34.22677, 34.21863, 34.21432, 
    34.20726, 34.20181, 34.19919, 34.19477, 34.18946, 34.1844, 34.17963, 
    34.17395, 34.17189, 34.17407, 34.17799, 34.17867, 34.17151, 34.14584, 
    34.08863, 33.99447, 33.86329, 33.69234, 33.40053, 32.69821, 32.1871, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  34.20464, 34.20523, 34.19534, 34.17819, 34.1608, 34.15195, 34.14743, 
    34.13984, 34.13413, 34.13162, 34.12713, 34.12166, 34.11646, 34.11179, 
    34.10735, 34.10635, 34.10833, 34.11178, 34.1127, 34.10653, 34.08429, 
    34.02407, 33.93114, 33.7829, 33.57646, 33.10933, 32.41041, 32.07688, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  34.12656, 34.12746, 34.11695, 34.09856, 34.08225, 34.07577, 34.07286, 
    34.06752, 34.06378, 34.06272, 34.0592, 34.05267, 34.04651, 34.04105, 
    34.03609, 34.03559, 34.03859, 34.04334, 34.04508, 34.03856, 34.01244, 
    33.95231, 33.83388, 33.66461, 33.4227, 32.76551, 32.15615, 32.03966, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  34.04645, 34.04764, 34.03715, 34.0162, 33.99675, 33.98871, 33.98518, 
    33.9781, 33.97314, 33.97176, 33.96843, 33.96413, 33.96011, 33.95748, 
    33.95547, 33.95724, 33.96071, 33.96581, 33.96877, 33.96461, 33.93475, 
    33.84853, 33.71637, 33.51746, 33.1027, 32.37551, 31.99468, 32.00937, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  33.95308, 33.95348, 33.94399, 33.92742, 33.90358, 33.89143, 33.88561, 
    33.87391, 33.8652, 33.86165, 33.85584, 33.84886, 33.8426, 33.83804, 
    33.83549, 33.83974, 33.84634, 33.85603, 33.86335, 33.86048, 33.82951, 
    33.72353, 33.57855, 33.30906, 32.68213, 32.09582, 31.96465, 32.00817, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  33.84758, 33.84616, 33.83211, 33.80852, 33.78439, 33.7729, 33.76585, 
    33.74723, 33.73278, 33.72549, 33.71579, 33.70467, 33.69471, 33.68666, 
    33.68298, 33.69065, 33.70155, 33.71791, 33.73196, 33.73103, 33.68971, 
    33.57403, 33.40798, 32.97905, 32.29026, 31.9689, 31.94553, 32.00717, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  33.72155, 33.71767, 33.69692, 33.66325, 33.62833, 33.61034, 33.60035, 
    33.58115, 33.56617, 33.55643, 33.54091, 33.5236, 33.50792, 33.49385, 
    33.48787, 33.50004, 33.51694, 33.54265, 33.56643, 33.56794, 33.5171, 
    33.39239, 33.1134, 32.51374, 32.01844, 31.95165, 31.94466, 32.00667, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  33.56034, 33.55441, 33.52392, 33.47512, 33.42605, 33.40062, 33.38583, 
    33.35739, 33.33394, 33.31836, 33.30423, 33.28111, 33.2555, 33.2288, 
    33.21579, 33.23171, 33.26046, 33.3021, 33.34104, 33.34499, 33.27457, 
    33.08128, 32.63927, 32.17152, 32.0137, 31.94572, 31.94396, 32.00658, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  33.31736, 33.31221, 33.26689, 33.19278, 33.12225, 33.08768, 33.06794, 
    33.02922, 32.99591, 32.97174, 32.95067, 32.92058, 32.88664, 32.84494, 
    32.81877, 32.82523, 32.87294, 32.93692, 32.99517, 33.00135, 32.88515, 
    32.56361, 32.26266, 32.08372, 32.01059, 31.94506, 31.94362, 32.00652, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  32.94391, 32.9424, 32.90029, 32.82822, 32.76496, 32.73141, 32.70568, 
    32.66984, 32.63469, 32.60318, 32.57518, 32.54998, 32.51975, 32.48688, 
    32.46146, 32.44347, 32.46487, 32.50056, 32.5414, 32.55213, 32.45293, 
    32.22535, 32.13184, 32.07829, 32.0098, 31.94454, 31.94338, 32.00646, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  32.68126, 32.67858, 32.67176, 32.66088, 32.65678, 32.64782, 32.63354, 
    32.62144, 32.60484, 32.58391, 32.5624, 32.53363, 32.49774, 32.46655, 
    32.43383, 32.39956, 32.34974, 32.31109, 32.28349, 32.26075, 32.21816, 
    32.15663, 32.12579, 32.07788, 32.00917, 31.94413, 31.94318, 32.00642, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  32.67618, 32.67316, 32.66665, 32.65665, 32.65358, 32.64487, 32.6305, 
    32.61883, 32.6027, 32.58213, 32.56107, 32.5328, 32.4973, 32.46612, 
    32.43322, 32.39861, 32.34748, 32.30772, 32.27923, 32.25281, 32.21008, 
    32.15317, 32.12558, 32.07753, 32.00866, 31.9438, 31.94305, 32.00642, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  32.67564, 32.67264, 32.66614, 32.65612, 32.65308, 32.64434, 32.62989, 
    32.61821, 32.60212, 32.58163, 32.5607, 32.5325, 32.49703, 32.46585, 
    32.43291, 32.39819, 32.34681, 32.30677, 32.27806, 32.25114, 32.20942, 
    32.1529, 32.12537, 32.07722, 32.00824, 31.94361, 31.94305, 32.00642, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  32.67534, 32.67232, 32.6658, 32.65578, 32.65274, 32.64396, 32.62941, 
    32.61771, 32.60164, 32.58119, 32.56036, 32.53221, 32.49672, 32.46555, 
    32.43258, 32.39781, 32.34643, 32.30638, 32.27765, 32.25072, 32.20904, 
    32.1526, 32.12515, 32.07697, 32.00809, 31.94361, 31.94305, 32.00642, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  32.6751, 32.67205, 32.66552, 32.65549, 32.65247, 32.64365, 32.62905, 
    32.61735, 32.60128, 32.58085, 32.56009, 32.53194, 32.49642, 32.46527, 
    32.43229, 32.3975, 32.34615, 32.3061, 32.27734, 32.25042, 32.20879, 
    32.15244, 32.12508, 32.07697, 32.00809, 31.94361, 31.94305, 32.00642, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 
    33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319, 33.97319,
  34.66774, 34.66775, 34.66506, 34.66038, 34.65593, 34.6535, 34.65153, 
    34.64827, 34.64568, 34.6442, 34.64215, 34.63977, 34.63757, 34.63499, 
    34.63257, 34.63162, 34.63252, 34.63402, 34.63445, 34.63238, 34.6208, 
    34.59076, 34.51299, 34.38117, 34.23828, 34.08714, 33.92694, 33.70988, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  34.65948, 34.65948, 34.65699, 34.65116, 34.64395, 34.64072, 34.63898, 
    34.63606, 34.63363, 34.63211, 34.63009, 34.62603, 34.62233, 34.61811, 
    34.6142, 34.61273, 34.61422, 34.61664, 34.61735, 34.61421, 34.60217, 
    34.5624, 34.47485, 34.34349, 34.20387, 34.05814, 33.88428, 33.66178, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  34.65063, 34.65064, 34.64644, 34.63929, 34.63272, 34.62943, 34.62634, 
    34.62115, 34.61689, 34.61436, 34.61103, 34.60732, 34.60397, 34.60018, 
    34.59668, 34.59539, 34.59684, 34.59914, 34.59989, 34.59718, 34.58445, 
    34.53635, 34.44225, 34.31127, 34.17444, 34.02535, 33.84776, 33.62055, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  34.63947, 34.63948, 34.63564, 34.6281, 34.61647, 34.61128, 34.60848, 
    34.60375, 34.59989, 34.59764, 34.59463, 34.59125, 34.5882, 34.58324, 
    34.57718, 34.57492, 34.57735, 34.58131, 34.58256, 34.57764, 34.55805, 
    34.51311, 34.41422, 34.2813, 34.14361, 33.99471, 33.8163, 33.53903, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  34.62951, 34.62954, 34.62271, 34.61105, 34.60032, 34.59555, 34.593, 
    34.58867, 34.58419, 34.58041, 34.5753, 34.5695, 34.56419, 34.5582, 
    34.55262, 34.55055, 34.55279, 34.55646, 34.55767, 34.55317, 34.53516, 
    34.48148, 34.38184, 34.24886, 34.11583, 33.96812, 33.78542, 33.46367, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  34.61321, 34.61323, 34.6069, 34.59608, 34.58613, 34.57832, 34.57388, 
    34.5664, 34.56034, 34.55685, 34.55209, 34.5467, 34.54175, 34.53621, 
    34.53105, 34.52915, 34.53122, 34.53465, 34.5358, 34.53168, 34.51506, 
    34.4537, 34.35193, 34.22036, 34.09141, 33.94473, 33.7401, 33.39721, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  34.59862, 34.59864, 34.59274, 34.58023, 34.56324, 34.55565, 34.55154, 
    34.54461, 34.53899, 34.53576, 34.53133, 34.52629, 34.52167, 34.51654, 
    34.51118, 34.50834, 34.51127, 34.51512, 34.51624, 34.51152, 34.48652, 
    34.42883, 34.32516, 34.19485, 34.06954, 33.91814, 33.69946, 33.33752, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  34.58497, 34.585, 34.57492, 34.55773, 34.5419, 34.53485, 34.53104, 
    34.52461, 34.5194, 34.51641, 34.51217, 34.50481, 34.49804, 34.49049, 
    34.48343, 34.48077, 34.48343, 34.48796, 34.48939, 34.48353, 34.46008, 
    34.40443, 34.30059, 34.17142, 34.04684, 33.88609, 33.66208, 33.23452, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  34.56178, 34.5618, 34.55242, 34.53642, 34.5217, 34.51516, 34.51146, 34.502, 
    34.49435, 34.48997, 34.48395, 34.47707, 34.47071, 34.46372, 34.45715, 
    34.45467, 34.45707, 34.46122, 34.46249, 34.45703, 34.43504, 34.37419, 
    34.27325, 34.14493, 34.01941, 33.85572, 33.62664, 33.11776, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  34.53906, 34.53907, 34.53038, 34.51554, 34.49646, 34.48691, 34.48169, 
    34.47296, 34.46592, 34.4619, 34.4563, 34.44988, 34.44394, 34.43748, 
    34.4314, 34.42908, 34.43123, 34.43501, 34.43613, 34.43106, 34.41051, 
    34.34455, 34.24247, 34.11755, 33.99251, 33.82595, 33.56669, 33.00325, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  34.51607, 34.51608, 34.50621, 34.48482, 34.46515, 34.45637, 34.45157, 
    34.44358, 34.43714, 34.43349, 34.42832, 34.42237, 34.41685, 34.41093, 
    34.40339, 34.40038, 34.40306, 34.40783, 34.40915, 34.40242, 34.37551, 
    34.31456, 34.21132, 34.08985, 33.9653, 33.79583, 33.47964, 32.88744, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  34.4815, 34.48151, 34.47008, 34.45059, 34.4327, 34.42473, 34.42037, 
    34.41314, 34.40624, 34.40159, 34.39504, 34.38752, 34.38052, 34.37302, 
    34.36591, 34.36314, 34.36537, 34.36953, 34.37057, 34.36404, 34.33923, 
    34.28144, 34.17906, 34.06115, 33.93698, 33.7393, 33.38954, 32.75301, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  34.44254, 34.44255, 34.43228, 34.41477, 34.39458, 34.38451, 34.37901, 
    34.36992, 34.36266, 34.35863, 34.3528, 34.34604, 34.33969, 34.33305, 
    34.32669, 34.32417, 34.32593, 34.32945, 34.3302, 34.32389, 34.30127, 
    34.2378, 34.14031, 34.02204, 33.88655, 33.67768, 33.29002, 32.60672, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  34.39921, 34.39923, 34.38646, 34.36472, 34.34493, 34.33617, 34.3314, 
    34.32356, 34.31733, 34.31394, 34.30886, 34.30289, 34.29722, 34.29068, 
    34.28334, 34.28038, 34.28229, 34.28621, 34.28693, 34.27925, 34.25257, 
    34.19241, 34.09617, 33.97622, 33.83411, 33.6136, 33.0508, 32.45477, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  34.34073, 34.34085, 34.32992, 34.31123, 34.29433, 34.28529, 34.27985, 
    34.27095, 34.26396, 34.26028, 34.25466, 34.24799, 34.24159, 34.23522, 
    34.22898, 34.2264, 34.22766, 34.23064, 34.23088, 34.22347, 34.1994, 
    34.14087, 34.0512, 33.92937, 33.76724, 33.46656, 32.80712, 32.30356, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  34.2805, 34.28076, 34.2684, 34.24732, 34.22841, 34.22032, 34.21611, 
    34.20909, 34.20366, 34.20103, 34.19656, 34.19104, 34.18559, 34.1805, 
    34.17429, 34.17146, 34.17269, 34.17574, 34.17557, 34.16729, 34.14095, 
    34.08344, 33.98614, 33.85054, 33.66814, 33.3098, 32.5528, 32.15454, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  34.20614, 34.20676, 34.19698, 34.17999, 34.16265, 34.1539, 34.14952, 
    34.14201, 34.13634, 34.13385, 34.12934, 34.12361, 34.11789, 34.11287, 
    34.10777, 34.10579, 34.10659, 34.10888, 34.10863, 34.1011, 34.07819, 
    34.01737, 33.92073, 33.76789, 33.53209, 32.95243, 32.31382, 32.05577, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  34.12845, 34.1294, 34.11905, 34.1009, 34.08461, 34.07818, 34.07541, 
    34.07013, 34.06643, 34.06541, 34.06189, 34.05514, 34.04839, 34.04257, 
    34.0368, 34.03497, 34.03637, 34.03954, 34.03962, 34.03124, 34.00395, 
    33.94355, 33.82257, 33.64263, 33.33435, 32.59477, 32.1355, 31.99894, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  34.04892, 34.05017, 34.03994, 34.01952, 34.00024, 33.99233, 33.98906, 
    33.98214, 33.97735, 33.97611, 33.97289, 33.96818, 33.9632, 33.96003, 
    33.95681, 33.95662, 33.9578, 33.96052, 33.96094, 33.95436, 33.92346, 
    33.83916, 33.70092, 33.46006, 32.92567, 32.26965, 32.00544, 31.95128, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  33.95723, 33.95774, 33.94854, 33.93241, 33.90908, 33.89737, 33.89208, 
    33.88089, 33.87268, 33.86957, 33.86427, 33.85704, 33.84966, 33.84465, 
    33.84047, 33.84164, 33.84453, 33.85025, 33.85335, 33.84693, 33.81559, 
    33.71159, 33.54789, 33.18167, 32.50335, 32.08941, 31.94112, 31.93421, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  33.85509, 33.85394, 33.84061, 33.8181, 33.79438, 33.78326, 33.77699, 
    33.75961, 33.74642, 33.74022, 33.73188, 33.72108, 33.71008, 33.7021, 
    33.69627, 33.69899, 33.70309, 33.71249, 33.71947, 33.71194, 33.66878, 
    33.5494, 33.32235, 32.76332, 32.19681, 31.98162, 31.89493, 31.92007, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  33.73506, 33.73186, 33.71275, 33.68148, 33.64796, 33.631, 33.62232, 
    33.60451, 33.59113, 33.58302, 33.56932, 33.55225, 33.53473, 33.52078, 
    33.51084, 33.51422, 33.51784, 33.53145, 33.54325, 33.53052, 33.46531, 
    33.31545, 32.91293, 32.32169, 32.04131, 31.9283, 31.87541, 31.91075, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  33.57859, 33.57421, 33.54448, 33.49615, 33.44585, 33.42102, 33.4086, 
    33.38186, 33.36123, 33.34958, 33.34034, 33.31832, 33.28952, 33.26406, 
    33.24398, 33.24354, 33.24406, 33.26191, 33.27838, 33.25362, 33.14559, 
    32.89086, 32.42783, 32.11504, 32.00648, 31.89709, 31.85984, 31.90548, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  33.32598, 33.32376, 33.27914, 33.20429, 33.12922, 33.0948, 33.0794, 
    33.04222, 33.01295, 32.99551, 32.98601, 32.96009, 32.92218, 32.88443, 
    32.84817, 32.83036, 32.82437, 32.84067, 32.85596, 32.81999, 32.6774, 
    32.37076, 32.17549, 32.04394, 31.97965, 31.87829, 31.84906, 31.90124, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  32.94015, 32.94197, 32.90414, 32.83712, 32.77621, 32.74636, 32.72551, 
    32.69344, 32.66335, 32.63793, 32.61737, 32.5927, 32.55795, 32.52768, 
    32.49437, 32.45917, 32.42844, 32.41117, 32.40362, 32.37941, 32.31016, 
    32.18259, 32.08445, 32.02081, 31.95996, 31.86322, 31.84065, 31.89784, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  32.68339, 32.68399, 32.67997, 32.6715, 32.66907, 32.66112, 32.64653, 
    32.63591, 32.62145, 32.60337, 32.58315, 32.55556, 32.52191, 32.49416, 
    32.46217, 32.42595, 32.37246, 32.32745, 32.2909, 32.23918, 32.18716, 
    32.12578, 32.06282, 32.01267, 31.94384, 31.85102, 31.83392, 31.89579, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  32.67185, 32.67384, 32.67139, 32.66447, 32.66415, 32.65604, 32.64011, 
    32.63041, 32.61671, 32.59904, 32.57957, 32.55368, 32.52139, 32.49374, 
    32.46177, 32.42548, 32.37177, 32.32508, 32.28543, 32.23032, 32.17117, 
    32.10898, 32.06149, 32.00575, 31.92942, 31.84126, 31.82954, 31.89579, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  32.67131, 32.67326, 32.67073, 32.66372, 32.66337, 32.6551, 32.63888, 
    32.62915, 32.61545, 32.59778, 32.57838, 32.55254, 32.52027, 32.49263, 
    32.46061, 32.42422, 32.37035, 32.32327, 32.28297, 32.22779, 32.16936, 
    32.10741, 32.05975, 31.99905, 31.91778, 31.83544, 31.82954, 31.89579, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  32.67076, 32.6727, 32.67012, 32.66304, 32.66269, 32.65436, 32.63804, 
    32.62827, 32.61453, 32.59683, 32.5774, 32.55141, 32.51888, 32.49119, 
    32.45906, 32.42252, 32.36833, 32.32104, 32.28062, 32.22551, 32.16689, 
    32.10461, 32.05764, 31.99378, 31.91347, 31.83544, 31.82954, 31.89579, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647,
  32.67041, 32.67231, 32.66971, 32.66259, 32.66224, 32.65387, 32.63749, 
    32.62767, 32.61392, 32.59623, 32.57677, 32.55062, 32.51777, 32.49004, 
    32.45783, 32.42115, 32.36662, 32.31908, 32.27853, 32.22337, 32.16491, 
    32.10314, 32.057, 31.99378, 31.91347, 31.83544, 31.82954, 31.89579, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 
    33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647, 33.96647 ;
}
