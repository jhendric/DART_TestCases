netcdf Test {
dimensions:
	latitude = 5 ;
	longitude = 6 ;
	height = 30 ;
	time = UNLIMITED ; // (1 currently)
variables:
	double latitude(latitude) ;
		latitude:units = "degrees_north" ;
		latitude:long_name = "latitude" ;
		latitude:standard_name = "latitude" ;
	double longitude(longitude) ;
		longitude:units = "degrees_east" ;
		longitude:long_name = "longitude" ;
		longitude:standard_name = "longitude" ;
	double height(height) ;
		height:units = "metres" ;
		height:long_name = "height" ;
		height:standard_name = "height" ;
	double time(time) ;
		time:units = "Days since 1601-01-01" ;
		time:long_name = "Time (UT)" ;
		time:standard_name = "Time" ;
	double Ne(height, latitude, longitude) ;
		Ne:grid_mapping = "standard" ;
		Ne:units = "1E11 e/m^3" ;
		Ne:long_name = "electron density" ;
		Ne:coordinates = "latitude longitude" ;
	double TEC(time, latitude, longitude) ;
		TEC:grid_mapping = "standard" ;
		TEC:units = "1E16 e/m^2" ;
		TEC:long_name = "total electron content" ;
		TEC:coordinates = "latitude longitude" ;
	double Variance(time, latitude, longitude) ;
		Variance:grid_mapping = "standard" ;
		Variance:units = "1E16 e/m^2" ;
		Variance:long_name = "Variance of total electron content" ;
		Variance:coordinates = "latitude longitude" ;
		Variance:standard_name = "TEC variance" ;

// global attributes:
		:Conventions = "CF-1.5" ;
data:

 latitude = -33, -23, -13, -3, 7 ;

 longitude = -85, -75, -65, -55, -45, -35 ;

 height = 0, 100000, 150000, 200000, 250000, 300000, 350000, 400000, 450000, 
    500000, 550000, 600000, 650000, 700000, 750000, 800000, 850000, 900000, 
    950000, 1000000, 1100000, 1200000, 1300000, 1400000, 1500000, 1600000, 
    1700000, 1800000, 1900000, 2000000 ;

 time = 148841.166666667 ;

 Ne =
  -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, -0,
  -0, -0, -0, -0, -0, 0,
  -0, -0, -0, -0, 0, 0,
  0.1834, 0.21859, 0.23895, 0.24, 0.2266, 0.21661,
  0.15765, 0.16073, 0.19797, 0.18955, 0.15125, 0.12585,
  0.09983, 0.12462, 0.1634, 0.11041, 0.08311, 0.04074,
  0.07594, 0.12256, 0.13626, 0.04707, 0.01051, -0.02368,
  0.07421, 0.10249, 0.09042, 0.0223, -0.04515, -0.1018,
  0.30159, 0.37261, 0.41266, 0.42, 0.40664, 0.39932,
  0.25323, 0.27248, 0.34216, 0.32708, 0.26904, 0.23385,
  0.15918, 0.20914, 0.27829, 0.18571, 0.14295, 0.07693,
  0.12208, 0.20246, 0.2283, 0.07497, 0.01295, -0.04345,
  0.11772, 0.16677, 0.14841, 0.03433, -0.08596, -0.1886,
  0.71149, 0.83635, 0.90953, 0.90864, 0.84894, 0.80212,
  0.61693, 0.61634, 0.7533, 0.72176, 0.5688, 0.46439,
  0.39169, 0.47975, 0.62543, 0.42464, 0.31687, 0.14923,
  0.29709, 0.47463, 0.52486, 0.18476, 0.04461, -0.08788,
  0.29172, 0.3992, 0.35105, 0.08856, -0.16479, -0.37614,
  0.77966, 0.72245, 0.7059, 0.62211, 0.42861, 0.24306,
  0.76477, 0.55505, 0.58049, 0.56429, 0.3238, 0.11215,
  0.50263, 0.46375, 0.54401, 0.40405, 0.2547, 0.01688,
  0.36686, 0.50648, 0.51271, 0.23835, 0.11281, -0.02991,
  0.38323, 0.46364, 0.38887, 0.13149, -0.0079, -0.09957,
  0.48038, 0.25657, 0.15235, 0.02026, -0.22344, -0.46822,
  0.55742, 0.22504, 0.11958, 0.12744, -0.09155, -0.31645,
  0.38102, 0.22551, 0.19783, 0.1894, 0.067, -0.1321,
  0.26618, 0.29881, 0.25523, 0.18174, 0.13162, 0.0461,
  0.2979, 0.31111, 0.24365, 0.11449, 0.16294, 0.24245,
  0.2553, 0.0113, -0.10644, -0.23001, -0.44208, -0.65868,
  0.35342, 0.04204, -0.09434, -0.07833, -0.24168, -0.42387,
  0.24981, 0.07991, 0.01405, 0.06116, -0.02404, -0.16472,
  0.16808, 0.15002, 0.0954, 0.11972, 0.11115, 0.06729,
  0.19928, 0.18222, 0.13218, 0.08304, 0.19789, 0.33033,
  0.12477, -0.07248, -0.16891, -0.26258, -0.41771, -0.57753,
  0.20838, -0.02783, -0.14459, -0.12938, -0.23851, -0.36663,
  0.15159, 0.01414, -0.04995, 0.00526, -0.04895, -0.13945,
  0.09875, 0.06784, 0.02153, 0.07294, 0.08002, 0.05958,
  0.12294, 0.09958, 0.06628, 0.05443, 0.16612, 0.2871,
  0.06716, -0.07028, -0.13778, -0.20154, -0.30568, -0.41334,
  0.12646, -0.03438, -0.11731, -0.10616, -0.17664, -0.26128,
  0.09342, -0.00238, -0.04967, -0.00705, -0.04126, -0.09869,
  0.05981, 0.03431, 0.00152, 0.04504, 0.05337, 0.04277,
  0.07642, 0.05782, 0.03635, 0.03485, 0.11724, 0.20491,
  0.04386, -0.04748, -0.09234, -0.13466, -0.20371, -0.27511,
  0.08331, -0.02343, -0.0786, -0.07117, -0.1178, -0.17386,
  0.06161, -0.00206, -0.03358, -0.0051, -0.0277, -0.06564,
  0.03939, 0.0223, 0.00049, 0.02971, 0.03537, 0.02847,
  0.05042, 0.03797, 0.02377, 0.02304, 0.07797, 0.13636,
  0.03322, -0.02882, -0.05925, -0.08825, -0.13585, -0.18499,
  0.05984, -0.01332, -0.05052, -0.04557, -0.07821, -0.11709,
  0.04396, 0.00072, -0.02024, -0.00161, -0.01758, -0.04433,
  0.02832, 0.01739, 0.00267, 0.02118, 0.02444, 0.01912,
  0.03585, 0.0278, 0.01785, 0.01618, 0.05271, 0.09179,
  0.0273, -0.01737, -0.03922, -0.06035, -0.09529, -0.1313,
  0.04628, -0.00703, -0.03354, -0.03007, -0.05451, -0.0833,
  0.03373, 0.00261, -0.01203, 0.00067, -0.01143, -0.03165,
  0.02192, 0.01473, 0.00422, 0.01624, 0.018, 0.01355,
  0.02739, 0.02199, 0.01453, 0.01218, 0.03769, 0.06524,
  0.02351, -0.01092, -0.02773, -0.04421, -0.07164, -0.09986,
  0.03802, -0.00355, -0.02379, -0.02118, -0.04072, -0.06349,
  0.02753, 0.00354, -0.00742, 0.00185, -0.00792, -0.02421,
  0.01802, 0.01297, 0.00494, 0.01324, 0.01418, 0.01029,
  0.02227, 0.0184, 0.01243, 0.00977, 0.02887, 0.04969,
  0.02093, -0.00737, -0.02117, -0.03484, -0.0577, -0.08121,
  0.03277, -0.0017, -0.01821, -0.01612, -0.03263, -0.05172,
  0.02362, 0.0039, -0.00489, 0.00239, -0.00593, -0.01978,
  0.01555, 0.01172, 0.00515, 0.01135, 0.01185, 0.00836,
  0.01906, 0.01606, 0.01102, 0.00828, 0.02361, 0.04046,
  0.01913, -0.00542, -0.01736, -0.0293, -0.04932, -0.06988,
  0.02934, -0.00074, -0.01498, -0.01319, -0.02778, -0.04457,
  0.02109, 0.00399, -0.00351, 0.0026, -0.00479, -0.01708,
  0.01393, 0.0108, 0.00513, 0.01013, 0.01039, 0.00719,
  0.01698, 0.0145, 0.01004, 0.00733, 0.0204, 0.03484,
  0.01785, -0.00434, -0.01513, -0.02596, -0.04417, -0.06285,
  0.02705, -0.00024, -0.01307, -0.01147, -0.02481, -0.04012,
  0.0194, 0.00395, -0.00276, 0.00265, -0.00413, -0.01539,
  0.01284, 0.01013, 0.00502, 0.00932, 0.00946, 0.00646,
  0.01561, 0.01343, 0.00935, 0.00672, 0.0184, 0.03136,
  0.01693, -0.00375, -0.0138, -0.02391, -0.04094, -0.05841,
  0.02549, -0, -0.01193, -0.01045, -0.02297, -0.0373,
  0.01826, 0.00386, -0.00234, 0.00263, -0.00374, -0.01432,
  0.0121, 0.00963, 0.00488, 0.00877, 0.00885, 0.006,
  0.01469, 0.01269, 0.00886, 0.0063, 0.01712, 0.02915,
  0.01627, -0.00343, -0.013, -0.02264, -0.03889, -0.05556,
  0.02441, 0.00011, -0.01125, -0.00983, -0.0218, -0.03549,
  0.01749, 0.00377, -0.00213, 0.00259, -0.00351, -0.01363,
  0.01159, 0.00927, 0.00474, 0.00839, 0.00845, 0.00571,
  0.01406, 0.01217, 0.00851, 0.00603, 0.0163, 0.02773,
  0.01579, -0.00326, -0.01252, -0.02185, -0.03758, -0.05371,
  0.02367, 0.00014, -0.01083, -0.00947, -0.02106, -0.03431,
  0.01695, 0.00368, -0.00202, 0.00253, -0.00338, -0.01318,
  0.01124, 0.009, 0.00463, 0.00814, 0.00818, 0.00552,
  0.01362, 0.0118, 0.00826, 0.00584, 0.01576, 0.02681,
  0.01544, -0.00318, -0.01223, -0.02136, -0.03674, -0.05251,
  0.02315, 0.00015, -0.01059, -0.00925, -0.02059, -0.03354,
  0.01657, 0.0036, -0.00197, 0.00248, -0.0033, -0.01289,
  0.01099, 0.0088, 0.00453, 0.00796, 0.008, 0.00539,
  0.01332, 0.01155, 0.00808, 0.00571, 0.01541, 0.02621,
  0.01501, -0.00314, -0.01196, -0.02086, -0.03584, -0.05121,
  0.02253, 0.00011, -0.01035, -0.00905, -0.02009, -0.03271,
  0.01613, 0.00348, -0.00195, 0.00239, -0.00323, -0.01256,
  0.0107, 0.00856, 0.00439, 0.00774, 0.00779, 0.00526,
  0.01297, 0.01123, 0.00786, 0.00556, 0.01503, 0.02556,
  0.01479, -0.00316, -0.01188, -0.02067, -0.03547, -0.05066,
  0.02222, 7e-05, -0.01028, -0.00899, -0.01989, -0.03235,
  0.01591, 0.00341, -0.00196, 0.00234, -0.00321, -0.01242,
  0.01055, 0.00842, 0.0043, 0.00764, 0.0077, 0.0052,
  0.01279, 0.01107, 0.00774, 0.00549, 0.01486, 0.02528,
  0.01468, -0.00318, -0.01186, -0.0206, -0.03532, -0.05042,
  0.02207, 4e-05, -0.01026, -0.00898, -0.01981, -0.0322,
  0.01581, 0.00337, -0.00198, 0.00231, -0.00321, -0.01236,
  0.01048, 0.00835, 0.00425, 0.00759, 0.00765, 0.00518,
  0.01271, 0.01099, 0.00768, 0.00545, 0.01478, 0.02516,
  0.01462, -0.0032, -0.01186, -0.02057, -0.03525, -0.05031,
  0.02199, 2e-05, -0.01026, -0.00898, -0.01977, -0.03213,
  0.01576, 0.00335, -0.002, 0.00229, -0.00321, -0.01234,
  0.01044, 0.00832, 0.00422, 0.00757, 0.00763, 0.00517,
  0.01267, 0.01095, 0.00765, 0.00544, 0.01475, 0.02511,
  0.01459, -0.00321, -0.01186, -0.02057, -0.03523, -0.05027,
  0.02195, 1e-05, -0.01026, -0.00898, -0.01976, -0.0321,
  0.01573, 0.00333, -0.00201, 0.00228, -0.00321, -0.01233,
  0.01042, 0.0083, 0.00421, 0.00755, 0.00762, 0.00516,
  0.01265, 0.01093, 0.00763, 0.00543, 0.01474, 0.02509,
  0.01457, -0.00322, -0.01186, -0.02056, -0.03522, -0.05025,
  0.02194, 0, -0.01026, -0.00898, -0.01976, -0.03209,
  0.01572, 0.00333, -0.00201, 0.00227, -0.00321, -0.01232,
  0.01042, 0.00829, 0.0042, 0.00755, 0.00762, 0.00516,
  0.01264, 0.01092, 0.00763, 0.00543, 0.01473, 0.02508,
  0.01456, -0.00322, -0.01187, -0.02056, -0.03521, -0.05024,
  0.02193, 0, -0.01026, -0.00898, -0.01975, -0.03208,
  0.01571, 0.00332, -0.00201, 0.00227, -0.00321, -0.01232,
  0.01041, 0.00829, 0.0042, 0.00754, 0.00761, 0.00516,
  0.01263, 0.01092, 0.00762, 0.00542, 0.01473, 0.02507,
  0.01456, -0.00322, -0.01187, -0.02056, -0.03521, -0.05024,
  0.02192, -0, -0.01026, -0.00899, -0.01975, -0.03208,
  0.01571, 0.00332, -0.00202, 0.00227, -0.00322, -0.01232,
  0.01041, 0.00828, 0.0042, 0.00754, 0.00761, 0.00516,
  0.01263, 0.01091, 0.00762, 0.00542, 0.01473, 0.02507,
  0.01456, -0.00323, -0.01187, -0.02056, -0.03521, -0.05024,
  0.02192, -0, -0.01026, -0.00899, -0.01975, -0.03208,
  0.01571, 0.00332, -0.00202, 0.00227, -0.00322, -0.01232,
  0.01041, 0.00828, 0.0042, 0.00754, 0.00761, 0.00516,
  0.01263, 0.01091, 0.00762, 0.00542, 0.01473, 0.02507,
  0.01456, -0.00323, -0.01187, -0.02056, -0.03521, -0.05024,
  0.02192, -0, -0.01027, -0.00899, -0.01975, -0.03208,
  0.01571, 0.00332, -0.00202, 0.00227, -0.00322, -0.01232,
  0.01041, 0.00828, 0.00419, 0.00754, 0.00761, 0.00516,
  0.01263, 0.01091, 0.00762, 0.00542, 0.01473, 0.02507 ;

 TEC =
  1.76592, 1.0933425, 0.78511, 0.363645, -0.433075, -1.22896,
  1.980425, 0.9204, 0.629235, 0.6439, -0.104725, -0.8561725,
  1.343835, 0.876945, 0.8366375, 0.7436775, 0.3178975, -0.3721275,
  0.9465175, 1.108995, 0.9865675, 0.6402975, 0.4343775, 0.1180575,
  1.0458625, 1.12339, 0.89244, 0.3942075, 0.465325, 0.6492875 ;

 Variance =
  22.4247280968008, 18.1858931308528, 14.9015471754668, 19.7896683978711, 
    16.7584127684643, 22.2977131707742,
  10.2268936775311, 4.36274813036854, 2.57970461420597, 5.97278948745223, 
    3.55583542580556, 15.390178636927,
  13.1743417574975, 7.5747651689139, 3.89180540387229, 1.82610318408633, 
    1.10799298654775, 8.9919813713478,
  18.2628993334102, 12.9084936434282, 2.46832689076766, 1, 1.5803853965816, 
    10.5128331898955,
  22.5883201513858, 22.3057730440516, 17.7044063463173, 7.6139520192543, 
    3.31843539395211, 14.9400267236203 ;
}
